* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt pixel gring VDD GND VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT CSA_VREF
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=7.5 as=24.809025 ps=56.34 w=2 l=1.44
X1 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.995 ps=8.8 w=1 l=0.8
X2 a_5720_n730# a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.25 pd=1.5 as=0.35 ps=2.7 w=1 l=1
X3 a_4330_n30# a_3852_n32# a_3852_n32# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.23 pd=1.65 as=0.3927 ps=2.8 w=1 l=2
X4 VDD SF_IB a_5720_n730# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.25 ps=1.5 w=1 l=1
X5 a_5460_10# a_4330_n30# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X6 a_3852_n32# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.76 ps=8.8 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=1
X8 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=1.995 pd=8.8 as=1.4 ps=7.4 w=7 l=0.15
X9 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.119375 pd=7.15 as=0 ps=0 w=2 l=3.35
X10 a_4120_n520# a_3852_n32# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X11 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=3.1 as=0.42 ps=3.1 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=2.95 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# VREF a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=1.4 pd=7.4 as=1.76 ps=8.8 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1.15
X16 VDD a_4330_n30# a_4330_n30# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.23 ps=1.65 w=1 l=2
X17 VDD a_5720_n730# a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.6 ps=2.95 w=1 l=0.15
X18 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X19 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=10.715 pd=15.9 as=0 ps=0 w=2.6 l=0.35
.ends

.subckt pixel_array VBIAS VREF NB2 VDD SF_IB CSA_VREF ROW_SEL0 ROW_SEL1 ROW_SEL2 PIX0_IN
+ GRING PIX1_IN PIX2_IN PIX3_IN PIX4_IN PIX5_IN PIX6_IN PIX_OUT0 PIX7_IN PIX_OUT1
+ PIX8_IN PIX_OUT2 ARRAY_OUT COL_SEL0 COL_SEl1 COL_SEL2 GND NB1
Xpixel_0 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX0_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel
Xpixel_1 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX1_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel
Xpixel_2 GRING VDD GND VREF ROW_SEL0 NB1 VBIAS NB2 PIX2_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel
Xpixel_3 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX3_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel
Xpixel_4 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX4_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel
Xpixel_5 GRING VDD GND VREF ROW_SEL1 NB1 VBIAS NB2 PIX5_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel
Xpixel_6 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX6_IN SF_IB PIX_OUT0 CSA_VREF
+ pixel
Xpixel_7 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX7_IN SF_IB PIX_OUT1 CSA_VREF
+ pixel
Xpixel_8 GRING VDD GND VREF ROW_SEL2 NB1 VBIAS NB2 PIX8_IN SF_IB PIX_OUT2 CSA_VREF
+ pixel
X0 PIX_OUT2 COL_SEL2 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X1 PIX_OUT1 COL_SEl1 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X2 PIX_OUT0 COL_SEL0 ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt shift_registerC COL_SEL[0] COL_SEL[10] COL_SEL[11] COL_SEL[12] COL_SEL[13]
+ COL_SEL[14] COL_SEL[15] COL_SEL[16] COL_SEL[17] COL_SEL[18] COL_SEL[19] COL_SEL[1]
+ COL_SEL[20] COL_SEL[21] COL_SEL[22] COL_SEL[23] COL_SEL[24] COL_SEL[25] COL_SEL[26]
+ COL_SEL[27] COL_SEL[28] COL_SEL[29] COL_SEL[2] COL_SEL[30] COL_SEL[31] COL_SEL[32]
+ COL_SEL[33] COL_SEL[34] COL_SEL[35] COL_SEL[36] COL_SEL[37] COL_SEL[38] COL_SEL[39]
+ COL_SEL[3] COL_SEL[40] COL_SEL[41] COL_SEL[42] COL_SEL[43] COL_SEL[44] COL_SEL[45]
+ COL_SEL[46] COL_SEL[47] COL_SEL[48] COL_SEL[49] COL_SEL[4] COL_SEL[50] COL_SEL[51]
+ COL_SEL[52] COL_SEL[53] COL_SEL[54] COL_SEL[55] COL_SEL[56] COL_SEL[57] COL_SEL[58]
+ COL_SEL[59] COL_SEL[5] COL_SEL[60] COL_SEL[61] COL_SEL[62] COL_SEL[63] COL_SEL[64]
+ COL_SEL[65] COL_SEL[66] COL_SEL[67] COL_SEL[68] COL_SEL[69] COL_SEL[6] COL_SEL[70]
+ COL_SEL[71] COL_SEL[72] COL_SEL[73] COL_SEL[74] COL_SEL[75] COL_SEL[76] COL_SEL[77]
+ COL_SEL[78] COL_SEL[79] COL_SEL[7] COL_SEL[80] COL_SEL[81] COL_SEL[82] COL_SEL[83]
+ COL_SEL[84] COL_SEL[85] COL_SEL[86] COL_SEL[87] COL_SEL[88] COL_SEL[89] COL_SEL[8]
+ COL_SEL[90] COL_SEL[91] COL_SEL[92] COL_SEL[93] COL_SEL[94] COL_SEL[95] COL_SEL[96]
+ COL_SEL[97] COL_SEL[98] COL_SEL[99] COL_SEL[9] clk data_in data_out ena rst VDD
+ GND
XFILLER_3_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_501_ _727_/Q _726_/Q _503_/S GND GND VDD VDD _502_/A sky130_fd_sc_hd__mux2_1
X_432_ _758_/Q _757_/Q _436_/S GND GND VDD VDD _433_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_363_ _789_/Q _788_/Q _369_/S GND GND VDD VDD _364_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2524 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2629 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1730 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_648 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_415_ _415_/A GND GND VDD VDD _766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3011 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3044 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_2310 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3105 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2343 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_3077 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1620 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1653 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2993 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1357 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1368 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_556 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2151 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_220 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_669 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_680_ _683_/A GND GND VDD VDD _680_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1110 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1154 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_397 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2220 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2097 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1341 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_732_ _773_/CLK _732_/D _618_/Y GND GND VDD VDD _732_/Q sky130_fd_sc_hd__dfrtp_1
X_663_ _664_/A GND GND VDD VDD _663_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_594_ _596_/A GND GND VDD VDD _594_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_868 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_5 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_3_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1625 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2094 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_359 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2871 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput7 _787_/Q GND GND VDD VDD COL_SEL[12] sky130_fd_sc_hd__clkbuf_1
Xoutput20 _699_/Q GND GND VDD VDD COL_SEL[24] sky130_fd_sc_hd__clkbuf_1
Xoutput31 _709_/Q GND GND VDD VDD COL_SEL[34] sky130_fd_sc_hd__clkbuf_1
Xoutput42 _719_/Q GND GND VDD VDD COL_SEL[44] sky130_fd_sc_hd__clkbuf_1
Xoutput53 _729_/Q GND GND VDD VDD COL_SEL[54] sky130_fd_sc_hd__clkbuf_1
Xoutput64 _739_/Q GND GND VDD VDD COL_SEL[64] sky130_fd_sc_hd__clkbuf_1
Xoutput75 _749_/Q GND GND VDD VDD COL_SEL[74] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput86 _759_/Q GND GND VDD VDD COL_SEL[84] sky130_fd_sc_hd__clkbuf_1
Xoutput97 _769_/Q GND GND VDD VDD COL_SEL[94] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_715_ _795_/CLK _715_/D _596_/Y GND GND VDD VDD _715_/Q sky130_fd_sc_hd__dfrtp_1
X_646_ _646_/A GND GND VDD VDD _646_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_577_ _578_/A GND GND VDD VDD _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2657 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_808 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1709 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2189 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_500_ _500_/A GND GND VDD VDD _728_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_6__f_clk clkbuf_0_clk/X GND GND VDD VDD _775_/CLK sky130_fd_sc_hd__clkbuf_16
X_431_ _431_/A GND GND VDD VDD _759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_362_ _362_/A GND GND VDD VDD _790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1802 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1929 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_963 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_629_ _633_/A GND GND VDD VDD _629_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1786 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2885 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_414_ _766_/Q _765_/Q _414_/S GND GND VDD VDD _415_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2405 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2377 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1676 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_281 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_579 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2163 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_276 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1166 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_332 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2508 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2232 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1397 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_445 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_731_ _773_/CLK _731_/D _617_/Y GND GND VDD VDD _731_/Q sky130_fd_sc_hd__dfrtp_1
X_662_ _664_/A GND GND VDD VDD _662_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_593_ _596_/A GND GND VDD VDD _593_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2585 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_8_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_6 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_3_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput8 _788_/Q GND GND VDD VDD COL_SEL[13] sky130_fd_sc_hd__clkbuf_1
Xoutput10 _790_/Q GND GND VDD VDD COL_SEL[15] sky130_fd_sc_hd__clkbuf_1
Xoutput21 _700_/Q GND GND VDD VDD COL_SEL[25] sky130_fd_sc_hd__clkbuf_1
Xoutput32 _710_/Q GND GND VDD VDD COL_SEL[35] sky130_fd_sc_hd__clkbuf_1
Xoutput43 _720_/Q GND GND VDD VDD COL_SEL[45] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput54 _730_/Q GND GND VDD VDD COL_SEL[55] sky130_fd_sc_hd__clkbuf_1
Xoutput65 _740_/Q GND GND VDD VDD COL_SEL[65] sky130_fd_sc_hd__clkbuf_1
Xoutput76 _750_/Q GND GND VDD VDD COL_SEL[75] sky130_fd_sc_hd__clkbuf_1
Xoutput87 _760_/Q GND GND VDD VDD COL_SEL[85] sky130_fd_sc_hd__clkbuf_1
Xoutput98 _770_/Q GND GND VDD VDD COL_SEL[95] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_714_ _786_/CLK _714_/D _595_/Y GND GND VDD VDD _714_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_611 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_645_ _646_/A GND GND VDD VDD _645_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_576_ _578_/A GND GND VDD VDD _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1401 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2124 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1423 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_430_ _759_/Q _758_/Q _436_/S GND GND VDD VDD _431_/A sky130_fd_sc_hd__mux2_1
X_361_ _790_/Q _789_/Q _369_/S GND GND VDD VDD _362_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_920 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_628_ _628_/A GND GND VDD VDD _633_/A sky130_fd_sc_hd__buf_2
XFILLER_18_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_559_ _701_/Q _700_/Q _559_/S GND GND VDD VDD _560_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2488 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_413_ _413_/A GND GND VDD VDD _767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2797 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1705 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_293 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2049 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_981 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3273 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2572 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1893 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2082 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2756 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_377 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_388 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_730_ _774_/CLK _730_/D _615_/Y GND GND VDD VDD _730_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_661_ _664_/A GND GND VDD VDD _661_/Y sky130_fd_sc_hd__inv_2
X_592_ _596_/A GND GND VDD VDD _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2807 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_7 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_3_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_317 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1173 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2895 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput9 _789_/Q GND GND VDD VDD COL_SEL[14] sky130_fd_sc_hd__clkbuf_1
Xoutput11 _791_/Q GND GND VDD VDD COL_SEL[16] sky130_fd_sc_hd__clkbuf_1
Xoutput22 _701_/Q GND GND VDD VDD COL_SEL[26] sky130_fd_sc_hd__clkbuf_1
Xoutput33 _711_/Q GND GND VDD VDD COL_SEL[36] sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_221 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xoutput44 _721_/Q GND GND VDD VDD COL_SEL[46] sky130_fd_sc_hd__clkbuf_1
Xoutput55 _731_/Q GND GND VDD VDD COL_SEL[56] sky130_fd_sc_hd__clkbuf_1
Xoutput66 _741_/Q GND GND VDD VDD COL_SEL[66] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput77 _751_/Q GND GND VDD VDD COL_SEL[76] sky130_fd_sc_hd__clkbuf_1
Xoutput88 _761_/Q GND GND VDD VDD COL_SEL[86] sky130_fd_sc_hd__clkbuf_1
Xoutput99 _771_/Q GND GND VDD VDD COL_SEL[96] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_713_ _786_/CLK _713_/D _594_/Y GND GND VDD VDD _713_/Q sky130_fd_sc_hd__dfrtp_1
X_644_ _646_/A GND GND VDD VDD _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_575_ _578_/A GND GND VDD VDD _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2615 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1903 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3285 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_409 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_360_ _393_/A GND GND VDD VDD _369_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2946 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_910 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_627_ _627_/A GND GND VDD VDD _627_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_558_ _558_/A GND GND VDD VDD _702_/D sky130_fd_sc_hd__clkbuf_1
X_489_ _489_/A GND GND VDD VDD _733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1243 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1254 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2710 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_412_ _767_/Q _766_/Q _414_/S GND GND VDD VDD _413_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_809 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2880 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2176 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2237 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2735 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2768 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1261 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_660_ _664_/A GND GND VDD VDD _660_/Y sky130_fd_sc_hd__inv_2
X_591_ _597_/A GND GND VDD VDD _596_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_827 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_304 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2819 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2598 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_8 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_10_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_789_ _791_/CLK _789_/D _688_/Y GND GND VDD VDD _789_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2031 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2086 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1116 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput12 _792_/Q GND GND VDD VDD COL_SEL[17] sky130_fd_sc_hd__clkbuf_1
Xoutput23 _702_/Q GND GND VDD VDD COL_SEL[27] sky130_fd_sc_hd__clkbuf_1
Xoutput34 _712_/Q GND GND VDD VDD COL_SEL[37] sky130_fd_sc_hd__clkbuf_1
Xoutput45 _722_/Q GND GND VDD VDD COL_SEL[47] sky130_fd_sc_hd__clkbuf_1
Xoutput56 _732_/Q GND GND VDD VDD COL_SEL[57] sky130_fd_sc_hd__clkbuf_1
Xoutput67 _742_/Q GND GND VDD VDD COL_SEL[67] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput78 _752_/Q GND GND VDD VDD COL_SEL[77] sky130_fd_sc_hd__clkbuf_1
Xoutput89 _762_/Q GND GND VDD VDD COL_SEL[87] sky130_fd_sc_hd__clkbuf_1
XFILLER_20_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_277 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_712_ _791_/CLK _712_/D _593_/Y GND GND VDD VDD _712_/Q sky130_fd_sc_hd__dfrtp_1
X_643_ _646_/A GND GND VDD VDD _643_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_574_ _578_/A GND GND VDD VDD _574_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2638 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_626_ _627_/A GND GND VDD VDD _626_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_557_ _702_/Q _701_/Q _559_/S GND GND VDD VDD _558_/A sky130_fd_sc_hd__mux2_1
X_488_ _733_/Q _732_/Q _492_/S GND GND VDD VDD _489_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1745 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2181 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_411_ _411_/A GND GND VDD VDD _768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3037 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_609_ _609_/A GND GND VDD VDD _609_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2265 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_416 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1597 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_1586 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2007 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1537 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_1476 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2040 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2051 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2095 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_780 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_357 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2013 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1284 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_590_ _590_/A GND GND VDD VDD _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_9 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_10_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_8 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_788_ _792_/CLK _788_/D _687_/Y GND GND VDD VDD _788_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2043 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2076 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2864 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1128 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput13 _793_/Q GND GND VDD VDD COL_SEL[18] sky130_fd_sc_hd__clkbuf_1
Xoutput24 _703_/Q GND GND VDD VDD COL_SEL[28] sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput35 _713_/Q GND GND VDD VDD COL_SEL[38] sky130_fd_sc_hd__clkbuf_1
Xoutput46 _723_/Q GND GND VDD VDD COL_SEL[48] sky130_fd_sc_hd__clkbuf_1
Xoutput57 _733_/Q GND GND VDD VDD COL_SEL[58] sky130_fd_sc_hd__clkbuf_1
Xoutput68 _743_/Q GND GND VDD VDD COL_SEL[68] sky130_fd_sc_hd__clkbuf_1
Xoutput79 _753_/Q GND GND VDD VDD COL_SEL[78] sky130_fd_sc_hd__clkbuf_1
X_711_ _786_/CLK _711_/D _592_/Y GND GND VDD VDD _711_/Q sky130_fd_sc_hd__dfrtp_1
X_642_ _646_/A GND GND VDD VDD _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_573_ _597_/A GND GND VDD VDD _578_/A sky130_fd_sc_hd__buf_2
XFILLER_16_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1916 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_clk clkbuf_0_clk/X GND GND VDD VDD _795_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1415 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2904 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2959 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_625_ _627_/A GND GND VDD VDD _625_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_956 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_556_ _556_/A GND GND VDD VDD _703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1702 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_487_ _487_/A GND GND VDD VDD _734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_410_ _768_/Q _767_/Q _414_/S GND GND VDD VDD _411_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_2723 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2778 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3005 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2337 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1625 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_608_ _609_/A GND GND VDD VDD _608_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_539_ _561_/A GND GND VDD VDD _548_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1565 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2965 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1885 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1373 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2940 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1513 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2069 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1313 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_818 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_787_ _795_/CLK _787_/D _686_/Y GND GND VDD VDD _787_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2055 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1093 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput14 _794_/Q GND GND VDD VDD COL_SEL[19] sky130_fd_sc_hd__clkbuf_1
Xoutput25 _704_/Q GND GND VDD VDD COL_SEL[29] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput36 _714_/Q GND GND VDD VDD COL_SEL[39] sky130_fd_sc_hd__clkbuf_1
Xoutput47 _724_/Q GND GND VDD VDD COL_SEL[49] sky130_fd_sc_hd__clkbuf_1
Xoutput58 _734_/Q GND GND VDD VDD COL_SEL[59] sky130_fd_sc_hd__clkbuf_1
Xoutput69 _744_/Q GND GND VDD VDD COL_SEL[69] sky130_fd_sc_hd__clkbuf_1
X_710_ _792_/CLK _710_/D _590_/Y GND GND VDD VDD _710_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_641_ _659_/A GND GND VDD VDD _646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_604 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_572_ _665_/A GND GND VDD VDD _597_/A sky130_fd_sc_hd__buf_2
XFILLER_16_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1630 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_0 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2117 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_624_ _627_/A GND GND VDD VDD _624_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_555_ _703_/Q _702_/Q _559_/S GND GND VDD VDD _556_/A sky130_fd_sc_hd__mux2_1
X_486_ _734_/Q _733_/Q _492_/S GND GND VDD VDD _487_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1758 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1268 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1648 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_607_ _609_/A GND GND VDD VDD _607_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_538_ _538_/A GND GND VDD VDD _711_/D sky130_fd_sc_hd__clkbuf_1
X_469_ _469_/A GND GND VDD VDD _742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2919 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1087 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2565 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2124 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_2157 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_1401 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_584 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2952 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2741 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2749 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1369 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2760 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_417 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_786_ _786_/CLK _786_/D _685_/Y GND GND VDD VDD _786_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_340 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2170 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput15 _776_/Q GND GND VDD VDD COL_SEL[1] sky130_fd_sc_hd__clkbuf_1
Xoutput26 _777_/Q GND GND VDD VDD COL_SEL[2] sky130_fd_sc_hd__clkbuf_1
Xoutput37 _778_/Q GND GND VDD VDD COL_SEL[3] sky130_fd_sc_hd__clkbuf_1
Xoutput48 _779_/Q GND GND VDD VDD COL_SEL[4] sky130_fd_sc_hd__clkbuf_1
Xoutput59 _780_/Q GND GND VDD VDD COL_SEL[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_640_ _640_/A GND GND VDD VDD _640_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_571_ _571_/A GND GND VDD VDD _696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1642 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_781 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_769_ _771_/CLK _769_/D _663_/Y GND GND VDD VDD _769_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_1 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1940 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_623_ _627_/A GND GND VDD VDD _623_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_936 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_554_ _554_/A GND GND VDD VDD _704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_485_ _485_/A GND GND VDD VDD _735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2195 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_980 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2950 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2736 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_606_ _609_/A GND GND VDD VDD _606_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_537_ _711_/Q _710_/Q _537_/S GND GND VDD VDD _538_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2202 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2257 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_468_ _742_/Q _741_/Q _470_/S GND GND VDD VDD _469_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1578 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_399_ _399_/A GND GND VDD VDD _773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_920 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2577 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_clk clkbuf_0_clk/X GND GND VDD VDD _773_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1424 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_249 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2964 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2797 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_360 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_1298 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2772 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3273 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_785_ _792_/CLK _785_/D _683_/Y GND GND VDD VDD _785_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1145 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1109 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput16 _795_/Q GND GND VDD VDD COL_SEL[20] sky130_fd_sc_hd__clkbuf_1
Xoutput27 _705_/Q GND GND VDD VDD COL_SEL[30] sky130_fd_sc_hd__clkbuf_1
Xoutput38 _715_/Q GND GND VDD VDD COL_SEL[40] sky130_fd_sc_hd__clkbuf_1
Xoutput49 _725_/Q GND GND VDD VDD COL_SEL[50] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_570_ _696_/Q _795_/Q _570_/S GND GND VDD VDD _571_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2090 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_768_ _775_/CLK _768_/D _662_/Y GND GND VDD VDD _768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_699_ _786_/CLK _699_/D _577_/Y GND GND VDD VDD _699_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk GND GND VDD VDD clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_15_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_622_ _628_/A GND GND VDD VDD _627_/A sky130_fd_sc_hd__clkbuf_2
X_553_ _704_/Q _703_/Q _559_/S GND GND VDD VDD _554_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_484_ _735_/Q _734_/Q _492_/S GND GND VDD VDD _485_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_992 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2962 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2494 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1782 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_605_ _609_/A GND GND VDD VDD _605_/Y sky130_fd_sc_hd__inv_2
X_536_ _536_/A GND GND VDD VDD _712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_467_ _467_/A GND GND VDD VDD _743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_398_ _773_/Q _772_/Q _402_/S GND GND VDD VDD _399_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2852 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2100 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2209 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1469 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_519_ _519_/A GND GND VDD VDD _720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1387 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1970 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2729 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_851 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_1200 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1233 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_394 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2784 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_29 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_1_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2573 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_784_ _795_/CLK _784_/D _682_/Y GND GND VDD VDD _784_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_865 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2857 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput17 _696_/Q GND GND VDD VDD COL_SEL[21] sky130_fd_sc_hd__clkbuf_1
Xoutput28 _706_/Q GND GND VDD VDD COL_SEL[31] sky130_fd_sc_hd__clkbuf_1
Xoutput39 _716_/Q GND GND VDD VDD COL_SEL[41] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_249 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1677 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_767_ _771_/CLK _767_/D _661_/Y GND GND VDD VDD _767_/Q sky130_fd_sc_hd__dfrtp_1
X_698_ _795_/CLK _698_/D _576_/Y GND GND VDD VDD _698_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_621_ _621_/A GND GND VDD VDD _621_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_415 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_437 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_949 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_552_ _552_/A GND GND VDD VDD _705_/D sky130_fd_sc_hd__clkbuf_1
X_483_ _505_/A GND GND VDD VDD _492_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2153 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2974 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1761 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_604_ _628_/A GND GND VDD VDD _609_/A sky130_fd_sc_hd__buf_2
XFILLER_18_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_535_ _712_/Q _711_/Q _537_/S GND GND VDD VDD _536_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1503 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_466_ _743_/Q _742_/Q _470_/S GND GND VDD VDD _467_/A sky130_fd_sc_hd__mux2_1
X_397_ _397_/A GND GND VDD VDD _774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2893 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2524 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1801 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2112 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_518_ _720_/Q _719_/Q _526_/S GND GND VDD VDD _519_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2045 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_449_ _449_/A GND GND VDD VDD _458_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_785 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1620 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1256 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2796 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1873 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1804 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_921 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_783_ _795_/CLK _783_/D _681_/Y GND GND VDD VDD _783_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_822 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_354 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1042 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput18 _697_/Q GND GND VDD VDD COL_SEL[22] sky130_fd_sc_hd__clkbuf_1
Xoutput29 _707_/Q GND GND VDD VDD COL_SEL[32] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_766_ _773_/CLK _766_/D _660_/Y GND GND VDD VDD _766_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_697_ _792_/CLK _697_/D _575_/Y GND GND VDD VDD _697_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2611 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_620_ _621_/A GND GND VDD VDD _620_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_551_ _705_/Q _704_/Q _559_/S GND GND VDD VDD _552_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_449 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_482_ _482_/A GND GND VDD VDD _736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_2110 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_749_ _774_/CLK _749_/D _639_/Y GND GND VDD VDD _749_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2986 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1228 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2474 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1740 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_603_ _665_/A GND GND VDD VDD _628_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_534_ _534_/A GND GND VDD VDD _713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1515 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_465_ _465_/A GND GND VDD VDD _744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_396_ _796_/A _773_/Q _402_/S GND GND VDD VDD _397_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2937 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2783 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2536 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2124 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1581 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_577 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_517_ _561_/A GND GND VDD VDD _526_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2901 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_208 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_448_ _448_/A GND GND VDD VDD _751_/D sky130_fd_sc_hd__clkbuf_1
X_379_ _379_/A GND GND VDD VDD _782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_720 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_742 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_308 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2208 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1676 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_875 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_897 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3193 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1816 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_561 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_782_ _791_/CLK _782_/D _680_/Y GND GND VDD VDD _782_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_977 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_834 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_366 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1451 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2185 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1065 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput19 _698_/Q GND GND VDD VDD COL_SEL[23] sky130_fd_sc_hd__clkbuf_1
XFILLER_6_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_765_ _775_/CLK _765_/D _658_/Y GND GND VDD VDD _765_/Q sky130_fd_sc_hd__dfrtp_1
X_696_ _786_/CLK _696_/D _574_/Y GND GND VDD VDD _696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_5 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2870 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_550_ _561_/A GND GND VDD VDD _559_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_428 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_481_ _736_/Q _735_/Q _481_/S GND GND VDD VDD _482_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2188 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_748_ _771_/CLK _748_/D _638_/Y GND GND VDD VDD _748_/Q sky130_fd_sc_hd__dfrtp_1
X_679_ _683_/A GND GND VDD VDD _679_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_450 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_602_ _602_/A GND GND VDD VDD _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_533_ _713_/Q _712_/Q _537_/S GND GND VDD VDD _534_/A sky130_fd_sc_hd__mux2_1
X_464_ _744_/Q _743_/Q _470_/S GND GND VDD VDD _465_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1527 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_395_ _395_/A GND GND VDD VDD _775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2811 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1004 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2795 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_2__f_clk clkbuf_0_clk/X GND GND VDD VDD _786_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2548 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2129 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_516_ _516_/A GND GND VDD VDD _561_/A sky130_fd_sc_hd__buf_2
XFILLER_18_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1313 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2058 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_447_ _751_/Q _750_/Q _447_/S GND GND VDD VDD _448_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_378_ _782_/Q _781_/Q _380_/S GND GND VDD VDD _379_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1379 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2713 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2685 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2592 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1611 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_353 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_375 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_887 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_386 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2460 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_551 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_584 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_781_ _795_/CLK _781_/D _679_/Y GND GND VDD VDD _781_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1430 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_378 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1463 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2017 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1088 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2083 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_753 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_764_ _771_/CLK _764_/D _657_/Y GND GND VDD VDD _764_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_695_ _695_/A GND GND VDD VDD _695_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_6 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2181 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_480_ _480_/A GND GND VDD VDD _737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_747_ _773_/CLK _747_/D _637_/Y GND GND VDD VDD _747_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_678_ _690_/A GND GND VDD VDD _683_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_462 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2487 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1775 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_601_ _602_/A GND GND VDD VDD _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_532_ _532_/A GND GND VDD VDD _714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_463_ _463_/A GND GND VDD VDD _745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_394_ _775_/Q input1/X _402_/S GND GND VDD VDD _395_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1252 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2801 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2823 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_925 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2516 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1815 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_515_ _515_/A GND GND VDD VDD _721_/D sky130_fd_sc_hd__clkbuf_1
X_446_ _446_/A GND GND VDD VDD _752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_377_ _377_/A GND GND VDD VDD _783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1093 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2697 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_1985 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2769 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_844 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_429_ _429_/A GND GND VDD VDD _760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_2891 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xinput1 data_in GND GND VDD VDD input1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3245 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_780_ _795_/CLK _780_/D _677_/Y GND GND VDD VDD _780_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_313 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1475 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1012 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1117 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_360 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_393 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_763_ _771_/CLK _763_/D _656_/Y GND GND VDD VDD _763_/Q sky130_fd_sc_hd__dfrtp_1
X_694_ _695_/A GND GND VDD VDD _694_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_7 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1250 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1681 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_408 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1481 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1423 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_746_ _773_/CLK _746_/D _636_/Y GND GND VDD VDD _746_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_677_ _677_/A GND GND VDD VDD _677_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1754 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_600_ _602_/A GND GND VDD VDD _600_/Y sky130_fd_sc_hd__inv_2
X_531_ _714_/Q _713_/Q _537_/S GND GND VDD VDD _532_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_462_ _745_/Q _744_/Q _470_/S GND GND VDD VDD _463_/A sky130_fd_sc_hd__mux2_1
X_393_ _393_/A GND GND VDD VDD _402_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_12_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1264 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2857 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_729_ _773_/CLK _729_/D _614_/Y GND GND VDD VDD _729_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2720 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2753 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_948 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1827 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1595 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_514_ _721_/Q _720_/Q _514_/S GND GND VDD VDD _515_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_445_ _752_/Q _751_/Q _447_/S GND GND VDD VDD _446_/A sky130_fd_sc_hd__mux2_1
X_376_ _783_/Q _782_/Q _380_/S GND GND VDD VDD _377_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_701 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1205 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1112 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_428_ _760_/Q _759_/Q _436_/S GND GND VDD VDD _429_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1145 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_359_ _359_/A GND GND VDD VDD _791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xinput2 ena GND GND VDD VDD _516_/A sky130_fd_sc_hd__buf_6
XFILLER_0_2545 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_520 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1690 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2122 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_347 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1487 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1024 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3021 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_762_ _773_/CLK _762_/D _655_/Y GND GND VDD VDD _762_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_693_ _695_/A GND GND VDD VDD _693_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_8 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2604 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1947 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_585 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_745_ _771_/CLK _745_/D _633_/Y GND GND VDD VDD _745_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_676_ _677_/A GND GND VDD VDD _676_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_530_ _530_/A GND GND VDD VDD _715_/D sky130_fd_sc_hd__clkbuf_1
X_461_ _505_/A GND GND VDD VDD _470_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_392_ _392_/A GND GND VDD VDD _776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1276 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_728_ _773_/CLK _728_/D _613_/Y GND GND VDD VDD _728_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_659_ _659_/A GND GND VDD VDD _664_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_2710 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2776 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1839 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_513_ _513_/A GND GND VDD VDD _722_/D sky130_fd_sc_hd__clkbuf_1
X_444_ _444_/A GND GND VDD VDD _753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2916 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_375_ _375_/A GND GND VDD VDD _784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2677 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_581 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1625 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2050 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1228 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2860 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_427_ _449_/A GND GND VDD VDD _436_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_358_ _791_/Q _790_/Q _358_/S GND GND VDD VDD _359_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xinput3 rst GND GND VDD VDD _665_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1845 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_326 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_2145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1499 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3077 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2321 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1592 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1606 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_30 _771_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_761_ _775_/CLK _761_/D _654_/Y GND GND VDD VDD _761_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_692_ _695_/A GND GND VDD VDD _692_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_602 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_9 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2885 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1274 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_744_ _773_/CLK _744_/D _632_/Y GND GND VDD VDD _744_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_675_ _677_/A GND GND VDD VDD _675_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_421 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_443 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2936 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1060 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_281 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_460_ _516_/A GND GND VDD VDD _505_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_391_ _776_/Q _775_/Q _391_/S GND GND VDD VDD _392_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1244 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_1288 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_361 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2837 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2909 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_727_ _775_/CLK _727_/D _612_/Y GND GND VDD VDD _727_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_658_ _658_/A GND GND VDD VDD _658_/Y sky130_fd_sc_hd__inv_2
X_589_ _590_/A GND GND VDD VDD _589_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2766 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2210 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_512_ _722_/Q _721_/Q _514_/S GND GND VDD VDD _513_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_443_ _753_/Q _752_/Q _447_/S GND GND VDD VDD _444_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_374_ _784_/Q _783_/Q _380_/S GND GND VDD VDD _375_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2928 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1900 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2689 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_1977 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1704 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_368 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_426_ _426_/A GND GND VDD VDD _761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_357_ _357_/A GND GND VDD VDD _792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3165 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1534 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_949 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2157 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_611 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2680 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_409_ _409_/A GND GND VDD VDD _769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2250 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1621 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2377 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_20 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2076 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_760_ _773_/CLK _760_/D _652_/Y GND GND VDD VDD _760_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_691_ _695_/A GND GND VDD VDD _691_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_614 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1220 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2897 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_452 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1927 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1640 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_743_ _774_/CLK _743_/D _631_/Y GND GND VDD VDD _743_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_674_ _677_/A GND GND VDD VDD _674_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_956 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1960 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1768 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_390_ _390_/A GND GND VDD VDD _777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_726_ _773_/CLK _726_/D _611_/Y GND GND VDD VDD _726_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_657_ _658_/A GND GND VDD VDD _657_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_588_ _590_/A GND GND VDD VDD _588_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1808 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_511_ _511_/A GND GND VDD VDD _723_/D sky130_fd_sc_hd__clkbuf_1
X_442_ _442_/A GND GND VDD VDD _754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_373_ _373_/A GND GND VDD VDD _785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_709_ _792_/CLK _709_/D _589_/Y GND GND VDD VDD _709_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_594 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2041 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_425_ _761_/Q _760_/Q _425_/S GND GND VDD VDD _426_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1126 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_356_ _792_/Q _791_/Q _358_/S GND GND VDD VDD _357_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_2748 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3144 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_589 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_10_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_408_ _769_/Q _768_/Q _414_/S GND GND VDD VDD _409_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2262 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1677 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1619 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XANTENNA_21 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_10 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_725 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_690_ _690_/A GND GND VDD VDD _695_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_626 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_475 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2618 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1652 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2153 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1416 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_742_ _774_/CLK _742_/D _630_/Y GND GND VDD VDD _742_/Q sky130_fd_sc_hd__dfrtp_1
X_673_ _677_/A GND GND VDD VDD _673_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_968 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1972 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_261 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1747 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_725_ _773_/CLK _725_/D _609_/Y GND GND VDD VDD _725_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_656_ _658_/A GND GND VDD VDD _656_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_587_ _590_/A GND GND VDD VDD _587_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1780 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2223 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_510_ _723_/Q _722_/Q _514_/S GND GND VDD VDD _511_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_441_ _754_/Q _753_/Q _447_/S GND GND VDD VDD _442_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_372_ _785_/Q _784_/Q _380_/S GND GND VDD VDD _373_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_193 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_708_ _792_/CLK _708_/D _588_/Y GND GND VDD VDD _708_/Q sky130_fd_sc_hd__dfrtp_1
X_639_ _640_/A GND GND VDD VDD _639_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1639 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2064 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1396 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_805 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_304 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_424_ _424_/A GND GND VDD VDD _762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_2852 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_355_ _355_/A GND GND VDD VDD _793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3112 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3217 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2444 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3156 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_3178 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1732 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_893 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_clk clkbuf_0_clk/X GND GND VDD VDD _792_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_407_ _407_/A GND GND VDD VDD _770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_22 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_11 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_20_332 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1491 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1480 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_638 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1108 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_410 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_465 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_487 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1664 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1453 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_501 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_741_ _774_/CLK _741_/D _629_/Y GND GND VDD VDD _741_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_672_ _690_/A GND GND VDD VDD _677_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1984 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_295 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_724_ _775_/CLK _724_/D _608_/Y GND GND VDD VDD _724_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_2829 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_655_ _658_/A GND GND VDD VDD _655_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_586_ _590_/A GND GND VDD VDD _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2482 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1792 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2235 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_440_ _440_/A GND GND VDD VDD _755_/D sky130_fd_sc_hd__clkbuf_1
X_371_ _393_/A GND GND VDD VDD _380_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2780 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_707_ _792_/CLK _707_/D _587_/Y GND GND VDD VDD _707_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_638_ _640_/A GND GND VDD VDD _638_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_574 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_569_ _569_/A GND GND VDD VDD _697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2599 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_423_ _762_/Q _761_/Q _425_/S GND GND VDD VDD _424_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_354_ _793_/Q _792_/Q _358_/S GND GND VDD VDD _355_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3124 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2412 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2517 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_371 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_603 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_406_ _770_/Q _769_/Q _414_/S GND GND VDD VDD _407_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_341 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1971 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2297 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XANTENNA_23 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_12 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1201 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2881 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_499 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1621 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1676 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_174 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_740_ _771_/CLK _740_/D _627_/Y GND GND VDD VDD _740_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_557 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_671_ _671_/A GND GND VDD VDD _671_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_915 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_937 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_436 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2929 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1086 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_274 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2185 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_2196 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2940 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_723_ _792_/CLK _723_/D _607_/Y GND GND VDD VDD _723_/Q sky130_fd_sc_hd__dfrtp_1
X_654_ _658_/A GND GND VDD VDD _654_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_585_ _597_/A GND GND VDD VDD _590_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_370_ _370_/A GND GND VDD VDD _786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2792 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_706_ _792_/CLK _706_/D _586_/Y GND GND VDD VDD _706_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_637_ _640_/A GND GND VDD VDD _637_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_568_ _697_/Q _696_/Q _570_/S GND GND VDD VDD _569_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_499_ _728_/Q _727_/Q _503_/S GND GND VDD VDD _500_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_729 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_829 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_422_ _422_/A GND GND VDD VDD _763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_353_ _353_/A GND GND VDD VDD _794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_862 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1817 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_383 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2991 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_320 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_405_ _449_/A GND GND VDD VDD _414_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1983 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3049 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1564 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2150 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_13 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_18_2183 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_24 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2069 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1213 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1909 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2492 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1780 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2040 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1394 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_197 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_186 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_5_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_670_ _671_/A GND GND VDD VDD _670_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1920 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1180 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1285 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2952 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_333 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_722_ _786_/CLK _722_/D _606_/Y GND GND VDD VDD _722_/Q sky130_fd_sc_hd__dfrtp_1
X_653_ _659_/A GND GND VDD VDD _658_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_584_ _584_/A GND GND VDD VDD _584_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2473 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_705_ _792_/CLK _705_/D _584_/Y GND GND VDD VDD _705_/Q sky130_fd_sc_hd__dfrtp_1
X_636_ _640_/A GND GND VDD VDD _636_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_565 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_567_ _567_/A GND GND VDD VDD _698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_708 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_498_ _498_/A GND GND VDD VDD _729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2579 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1889 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_329 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_421_ _763_/Q _762_/Q _425_/S GND GND VDD VDD _422_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_2844 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_352_ _794_/Q _793_/Q _358_/S GND GND VDD VDD _353_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1119 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_6_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3137 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_852 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_619_ _621_/A GND GND VDD VDD _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_538 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1406 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2641 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_404_ _516_/A GND GND VDD VDD _449_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1995 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2349 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_14 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_25 _796_/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_11_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2460 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2081 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1340 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2096 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1409 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2880 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_928 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2622 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_950 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1420 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1192 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2964 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_389 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_721_ _786_/CLK _721_/D _605_/Y GND GND VDD VDD _721_/Q sky130_fd_sc_hd__dfrtp_1
X_652_ _652_/A GND GND VDD VDD _652_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_583_ _584_/A GND GND VDD VDD _583_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1061 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2761 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_704_ _792_/CLK _704_/D _583_/Y GND GND VDD VDD _704_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_635_ _659_/A GND GND VDD VDD _640_/A sky130_fd_sc_hd__buf_2
X_566_ _698_/Q _697_/Q _570_/S GND GND VDD VDD _567_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2514 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_497_ _729_/Q _728_/Q _503_/S GND GND VDD VDD _498_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2901 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2057 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_420_ _420_/A GND GND VDD VDD _764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_351_ _351_/A GND GND VDD VDD _795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_2867 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2437 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_330 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_618_ _621_/A GND GND VDD VDD _618_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_549_ _549_/A GND GND VDD VDD _706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1632 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_617 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_403_ _403_/A GND GND VDD VDD _771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_355 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1544 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1649 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_26 _770_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_15 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_11_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput100 _772_/Q GND GND VDD VDD COL_SEL[97] sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1237 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_892 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1793 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2125 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_144 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1270 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2634 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_962 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2280 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1432 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_720_ _786_/CLK _720_/D _602_/Y GND GND VDD VDD _720_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_651_ _652_/A GND GND VDD VDD _651_/Y sky130_fd_sc_hd__inv_2
X_582_ _584_/A GND GND VDD VDD _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2729 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1752 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3300 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_165 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_703_ _795_/CLK _703_/D _582_/Y GND GND VDD VDD _703_/Q sky130_fd_sc_hd__dfrtp_1
X_634_ _665_/A GND GND VDD VDD _659_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2526 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_565_ _565_/A GND GND VDD VDD _699_/D sky130_fd_sc_hd__clkbuf_1
X_496_ _496_/A GND GND VDD VDD _730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_350_ _795_/Q _794_/Q _358_/S GND GND VDD VDD _351_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1704 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_617_ _621_/A GND GND VDD VDD _617_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_364 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_548_ _706_/Q _705_/Q _548_/S GND GND VDD VDD _549_/A sky130_fd_sc_hd__mux2_1
X_479_ _737_/Q _736_/Q _481_/S GND GND VDD VDD _480_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1666 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2972 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2109 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1110 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_17_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_402_ _771_/Q _770_/Q _402_/S GND GND VDD VDD _403_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_40 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_334 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1964 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1556 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_304 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XANTENNA_27 _665_/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_16 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_20_337 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput101 _773_/Q GND GND VDD VDD COL_SEL[98] sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_437 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2010 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1425 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_156 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_429 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2646 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_796_ _796_/A GND GND VDD VDD _796_/X sky130_fd_sc_hd__buf_6
XFILLER_1_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_974 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2292 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1444 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_650_ _652_/A GND GND VDD VDD _650_/Y sky130_fd_sc_hd__inv_2
X_581_ _584_/A GND GND VDD VDD _581_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_779_ _791_/CLK _779_/D _676_/Y GND GND VDD VDD _779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_702_ _792_/CLK _702_/D _581_/Y GND GND VDD VDD _702_/Q sky130_fd_sc_hd__dfrtp_1
X_633_ _633_/A GND GND VDD VDD _633_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_564_ _699_/Q _698_/Q _570_/S GND GND VDD VDD _565_/A sky130_fd_sc_hd__mux2_1
X_495_ _730_/Q _729_/Q _503_/S GND GND VDD VDD _496_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2538 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2240 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2825 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2428 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_616_ _628_/A GND GND VDD VDD _621_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_547_ _547_/A GND GND VDD VDD _707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_508 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_478_ _478_/A GND GND VDD VDD _738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1678 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1100 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2880 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2600 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_30 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_401_ _401_/A GND GND VDD VDD _772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_2633 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_41 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_641 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_2269 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2176 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XANTENNA_28 _771_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_17 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_9_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput102 _796_/A GND GND VDD VDD COL_SEL[99] sky130_fd_sc_hd__clkbuf_1
XFILLER_9_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2853 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1228 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2073 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2894 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_529 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1913 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_795_ _795_/CLK _795_/D _695_/Y GND GND VDD VDD _795_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xclkbuf_3_4__f_clk clkbuf_0_clk/X GND GND VDD VDD _771_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1401 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1201 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_1173 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_580_ _584_/A GND GND VDD VDD _580_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_893 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_778_ _791_/CLK _778_/D _675_/Y GND GND VDD VDD _778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_701_ _795_/CLK _701_/D _580_/Y GND GND VDD VDD _701_/Q sky130_fd_sc_hd__dfrtp_1
X_632_ _633_/A GND GND VDD VDD _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_563_ _563_/A GND GND VDD VDD _700_/D sky130_fd_sc_hd__clkbuf_1
X_494_ _505_/A GND GND VDD VDD _503_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_13_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2252 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2915 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_615_ _615_/A GND GND VDD VDD _615_/Y sky130_fd_sc_hd__inv_2
X_546_ _707_/Q _706_/Q _548_/S GND GND VDD VDD _547_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_477_ _738_/Q _737_/Q _481_/S GND GND VDD VDD _478_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_400_ _772_/Q _771_/Q _402_/S GND GND VDD VDD _401_/A sky130_fd_sc_hd__mux2_1
XPHY_20 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_31 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_2656 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1900 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1569 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_529_ _715_/Q _714_/Q _537_/S GND GND VDD VDD _530_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1432 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_29 _771_/Q GND GND VDD VDD sky130_fd_sc_hd__diode_2
XANTENNA_18 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_14_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput103 _784_/Q GND GND VDD VDD COL_SEL[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_9_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_22 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2453 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2045 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1355 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1251 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2615 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1936 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_794_ _795_/CLK _794_/D _694_/Y GND GND VDD VDD _794_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_943 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2125 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_15_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1560 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_7_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1257 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_291 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_305 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_777_ _792_/CLK _777_/D _674_/Y GND GND VDD VDD _777_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2754 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_700_ _792_/CLK _700_/D _578_/Y GND GND VDD VDD _700_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_631_ _633_/A GND GND VDD VDD _631_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_562_ _700_/Q _699_/Q _570_/S GND GND VDD VDD _563_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2507 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1806 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_493_ _493_/A GND GND VDD VDD _731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2264 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_592 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2927 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_813 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_614_ _615_/A GND GND VDD VDD _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_545_ _545_/A GND GND VDD VDD _708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1603 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_476_ _476_/A GND GND VDD VDD _739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2997 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_3_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2860 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2624 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_10 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_21 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_2668 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_32 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_348 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1956 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_528_ _561_/A GND GND VDD VDD _537_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1411 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XANTENNA_19 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_18_1444 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_459_ _459_/A GND GND VDD VDD _746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput104 _796_/X GND GND VDD VDD data_out sky130_fd_sc_hd__clkbuf_1
XFILLER_9_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_885 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_34 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1731 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1628 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_974 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_137 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2685 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_1005 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_660 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1948 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_793_ _795_/CLK _793_/D _693_/Y GND GND VDD VDD _793_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3161 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1745 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_776_ _791_/CLK _776_/D _673_/Y GND GND VDD VDD _776_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1033 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_630_ _633_/A GND GND VDD VDD _630_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_561_ _561_/A GND GND VDD VDD _570_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_492_ _731_/Q _730_/Q _492_/S GND GND VDD VDD _493_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_759_ _773_/CLK _759_/D _651_/Y GND GND VDD VDD _759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1096 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2585 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_613_ _615_/A GND GND VDD VDD _613_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_346 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_544_ _708_/Q _707_/Q _548_/S GND GND VDD VDD _545_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_357 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_475_ _739_/Q _738_/Q _481_/S GND GND VDD VDD _476_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1648 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2095 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_880 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_11 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_22 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_33 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_327 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_633 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_1516 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_527_ _527_/A GND GND VDD VDD _716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_458_ _746_/Q _745_/Q _458_/S GND GND VDD VDD _459_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1456 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_389_ _777_/Q _776_/Q _391_/S GND GND VDD VDD _390_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_371 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_897 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_46 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_11_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1743 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_953 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1368 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1220 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2570 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1985 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_1927 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_805 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_792_ _792_/CLK _792_/D _692_/Y GND GND VDD VDD _792_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1061 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2461 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_1768 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_775_ _775_/CLK _775_/D _671_/Y GND GND VDD VDD _775_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2082 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_81 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1089 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_11_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_137 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_560_ _560_/A GND GND VDD VDD _701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_491_ _491_/A GND GND VDD VDD _732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_758_ _771_/CLK _758_/D _650_/Y GND GND VDD VDD _758_/Q sky130_fd_sc_hd__dfrtp_1
X_689_ _689_/A GND GND VDD VDD _689_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_612_ _615_/A GND GND VDD VDD _612_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1709 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_826 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_543_ _543_/A GND GND VDD VDD _709_/D sky130_fd_sc_hd__clkbuf_1
X_474_ _474_/A GND GND VDD VDD _740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_892 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2905 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_12 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_23 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_34 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1513 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1528 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_526_ _716_/Q _715_/Q _526_/S GND GND VDD VDD _527_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_309 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_457_ _457_/A GND GND VDD VDD _747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1424 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_2169 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_383 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_1468 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_388_ _388_/A GND GND VDD VDD _778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1393 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2445 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1788 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2088 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1533 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_921 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_509_ _509_/A GND GND VDD VDD _724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2887 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3261 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_791_ _791_/CLK _791_/D _691_/Y GND GND VDD VDD _791_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_935 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1761 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_470 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_774_ _774_/CLK _774_/D _670_/Y GND GND VDD VDD _796_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2768 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1981 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_490_ _732_/Q _731_/Q _492_/S GND GND VDD VDD _491_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2457 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_757_ _773_/CLK _757_/D _649_/Y GND GND VDD VDD _757_/Q sky130_fd_sc_hd__dfrtp_1
X_688_ _689_/A GND GND VDD VDD _688_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_2009 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1897 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_611_ _615_/A GND GND VDD VDD _611_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_542_ _709_/Q _708_/Q _548_/S GND GND VDD VDD _543_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_473_ _740_/Q _739_/Q _481_/S GND GND VDD VDD _474_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1341 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1385 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1085 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_13 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_24 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_35 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_2649 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_1650 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_525_ _525_/A GND GND VDD VDD _717_/D sky130_fd_sc_hd__clkbuf_1
X_456_ _747_/Q _746_/Q _458_/S GND GND VDD VDD _457_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_340 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_387_ _778_/Q _777_/Q _391_/S GND GND VDD VDD _388_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2825 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1723 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1767 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2027 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_421 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_966 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_508_ _724_/Q _723_/Q _514_/S GND GND VDD VDD _509_/A sky130_fd_sc_hd__mux2_1
X_439_ _755_/Q _754_/Q _447_/S GND GND VDD VDD _440_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_1277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2608 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_790_ _792_/CLK _790_/D _689_/Y GND GND VDD VDD _790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2577 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2210 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1397 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_69 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1704 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1759 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_637 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_865 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_773_ _773_/CLK _773_/D _669_/Y GND GND VDD VDD _773_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1673 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_1383 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2149 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2293 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2202 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1534 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1589 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_445 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_756_ _775_/CLK _756_/D _648_/Y GND GND VDD VDD _756_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_687_ _689_/A GND GND VDD VDD _687_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_15_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2577 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_610_ _628_/A GND GND VDD VDD _615_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_839 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_3009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_541_ _541_/A GND GND VDD VDD _710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_472_ _505_/A GND GND VDD VDD _481_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_1353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1397 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_12_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2233 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_2277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2979 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_739_ _771_/CLK _739_/D _626_/Y GND GND VDD VDD _739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_14 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_25 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_36 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1949 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1662 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_614 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_524_ _717_/Q _716_/Q _526_/S GND GND VDD VDD _525_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_2138 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_455_ _455_/A GND GND VDD VDD _748_/D sky130_fd_sc_hd__clkbuf_1
X_386_ _386_/A GND GND VDD VDD _779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2041 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput90 _763_/Q GND GND VDD VDD COL_SEL[88] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2661 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_878 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1481 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_945 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_466 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_507_ _507_/A GND GND VDD VDD _725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_438_ _449_/A GND GND VDD VDD _447_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_19_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_108 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_369_ _786_/Q _785_/Q _369_/S GND GND VDD VDD _370_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2601 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1861 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1872 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2244 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1587 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_10_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_775 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_19_753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1229 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_19_797 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1075 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2821 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1691 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1917 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_772_ _773_/CLK _772_/D _668_/Y GND GND VDD VDD _772_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2041 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1593 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_16_2269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_413 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_641 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_755_ _774_/CLK _755_/D _646_/Y GND GND VDD VDD _755_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_686_ _689_/A GND GND VDD VDD _686_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1089 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_5__f_clk clkbuf_0_clk/X GND GND VDD VDD _774_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_2501 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_540_ _710_/Q _709_/Q _548_/S GND GND VDD VDD _541_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_306 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_471_ _471_/A GND GND VDD VDD _741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1677 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1365 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_777 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2289 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_738_ _771_/CLK _738_/D _625_/Y GND GND VDD VDD _738_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_669_ _671_/A GND GND VDD VDD _669_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_309 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_15 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_26 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_37 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1674 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_1509 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_523_ _523_/A GND GND VDD VDD _718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_454_ _748_/Q _747_/Q _458_/S GND GND VDD VDD _455_/A sky130_fd_sc_hd__mux2_1
X_385_ _779_/Q _778_/Q _391_/S GND GND VDD VDD _386_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_81 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1140 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_1173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput80 _754_/Q GND GND VDD VDD COL_SEL[79] sky130_fd_sc_hd__clkbuf_1
Xoutput91 _764_/Q GND GND VDD VDD COL_SEL[89] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2097 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_813 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_12_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_434 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_506_ _725_/Q _724_/Q _514_/S GND GND VDD VDD _507_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_489 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_437_ _437_/A GND GND VDD VDD _756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_368_ _368_/A GND GND VDD VDD _787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2657 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1901 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2481 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_676 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1677 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2513 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2234 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_2256 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1408 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_853 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_897 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1609 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_721 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_765 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1953 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1817 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2877 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3133 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_27 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2429 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1441 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1929 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_771_ _771_/CLK _771_/D _667_/Y GND GND VDD VDD _771_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1396 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2573 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1005 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2738 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3185 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_3005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1625 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1761 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_2641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_281 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_469 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_697 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_754_ _775_/CLK _754_/D _645_/Y GND GND VDD VDD _754_/Q sky130_fd_sc_hd__dfrtp_1
X_685_ _689_/A GND GND VDD VDD _685_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1057 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1901 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1945 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1989 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2961 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_370 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_17_2557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_808 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_2493 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_470_ _741_/Q _740_/Q _470_/S GND GND VDD VDD _471_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2001 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2045 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_9_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1300 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_737_ _771_/CLK _737_/D _624_/Y GND GND VDD VDD _737_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_668_ _671_/A GND GND VDD VDD _668_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_599_ _602_/A GND GND VDD VDD _599_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2844 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_0 _690_/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_8_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_16 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_27 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_38 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1620 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_522_ _718_/Q _717_/Q _526_/S GND GND VDD VDD _523_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_453_ _453_/A GND GND VDD VDD _749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_384_ _384_/A GND GND VDD VDD _780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_93 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1005 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1049 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_553 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput70 _781_/Q GND GND VDD VDD COL_SEL[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2065 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput81 _782_/Q GND GND VDD VDD COL_SEL[7] sky130_fd_sc_hd__clkbuf_1
Xoutput92 _783_/Q GND GND VDD VDD COL_SEL[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_4_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2685 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_2505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1962 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_836 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1369 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_589 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2205 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_2249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1329 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_505_ _505_/A GND GND VDD VDD _514_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_436_ _756_/Q _755_/Q _436_/S GND GND VDD VDD _437_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_367_ _787_/Q _786_/Q _369_/S GND GND VDD VDD _368_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2869 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_13_3261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2531 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1957 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_18_2493 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_1645 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_688 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1509 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_917 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_928 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_405 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_449 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2268 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1578 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1280 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_10_165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1133 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_865 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2057 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_265 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_419_ _764_/Q _763_/Q _425_/S GND GND VDD VDD _420_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2633 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1088 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_1099 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_11_1829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3084 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2433 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_39 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3189 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_3109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1453 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1497 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_770_ _775_/CLK _770_/D _664_/Y GND GND VDD VDD _770_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_725 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_769 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_441 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_2953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2997 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2541 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_485 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2585 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_3017 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_1773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1637 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_109 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_6_2653 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2216 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1705 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1749 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_753_ _774_/CLK _753_/D _644_/Y GND GND VDD VDD _753_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2185 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_684_ _690_/A GND GND VDD VDD _689_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_533 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1957 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2393 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2569 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1401 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1581 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2013 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1312 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_473 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_736_ _773_/CLK _736_/D _623_/Y GND GND VDD VDD _736_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1281 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_667_ _671_/A GND GND VDD VDD _667_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_330 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_1_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_598_ _602_/A GND GND VDD VDD _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_897 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_1_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3101 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_2709 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_2867 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_3145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1721 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_3189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_1 _690_/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_6_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1765 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_17 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_28 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_39 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1643 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_3213 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1833 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_521_ _521_/A GND GND VDD VDD _719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_452_ _749_/Q _748_/Q _458_/S GND GND VDD VDD _453_/A sky130_fd_sc_hd__mux2_1
X_383_ _780_/Q _779_/Q _391_/S GND GND VDD VDD _384_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput60 _735_/Q GND GND VDD VDD COL_SEL[60] sky130_fd_sc_hd__clkbuf_1
Xoutput71 _745_/Q GND GND VDD VDD COL_SEL[70] sky130_fd_sc_hd__clkbuf_1
Xoutput82 _755_/Q GND GND VDD VDD COL_SEL[80] sky130_fd_sc_hd__clkbuf_1
Xoutput93 _765_/Q GND GND VDD VDD COL_SEL[90] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_719_ _786_/CLK _719_/D _601_/Y GND GND VDD VDD _719_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2631 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1974 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_609 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_3129 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2196 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_1337 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_458 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_504_ _504_/A GND GND VDD VDD _726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_435_ _435_/A GND GND VDD VDD _757_/D sky130_fd_sc_hd__clkbuf_1
X_366_ _366_/A GND GND VDD VDD _788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1449 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3211 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_3233 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_3244 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_3277 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_970 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_18_981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1886 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_612 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2325 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2093 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_417 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_1101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_177 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1145 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1189 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_321 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_877 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2069 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1116 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_277 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_418_ _418_/A GND GND VDD VDD _765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_349_ _393_/A GND GND VDD VDD _358_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_13_3081 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2689 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_693 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1213 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1257 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3096 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2384 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2489 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1733 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1421 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_486 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1329 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_3193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_225 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_737 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2033 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_16_2932 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1376 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3221 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2829 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_497 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2597 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1785 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1649 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1021 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2253 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2228 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1273 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_752_ _775_/CLK _752_/D _643_/Y GND GND VDD VDD _752_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_683_ _683_/A GND GND VDD VDD _683_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_2197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_501 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_545 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2773 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_261 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1925 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2361 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_961 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1413 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1593 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1457 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2902 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2058 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_2913 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_2681 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_735_ _771_/CLK _735_/D _621_/Y GND GND VDD VDD _735_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_666_ _690_/A GND GND VDD VDD _671_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_597_ _597_/A GND GND VDD VDD _602_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_581 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_3157 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_2 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_12_1733 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1777 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_2793 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_18 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_29 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_2345 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_1633 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_2389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2209 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3269 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1845 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_607 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1889 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_520_ _719_/Q _718_/Q _526_/S GND GND VDD VDD _521_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_451_ _451_/A GND GND VDD VDD _750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_382_ _393_/A GND GND VDD VDD _391_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1029 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput4 _775_/Q GND GND VDD VDD COL_SEL[0] sky130_fd_sc_hd__clkbuf_1
Xoutput50 _726_/Q GND GND VDD VDD COL_SEL[51] sky130_fd_sc_hd__clkbuf_1
Xoutput61 _736_/Q GND GND VDD VDD COL_SEL[61] sky130_fd_sc_hd__clkbuf_1
Xoutput72 _746_/Q GND GND VDD VDD COL_SEL[71] sky130_fd_sc_hd__clkbuf_1
Xoutput83 _756_/Q GND GND VDD VDD COL_SEL[81] sky130_fd_sc_hd__clkbuf_1
Xoutput94 _766_/Q GND GND VDD VDD COL_SEL[91] sky130_fd_sc_hd__clkbuf_1
XFILLER_4_2933 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_718_ _786_/CLK _718_/D _600_/Y GND GND VDD VDD _718_/Q sky130_fd_sc_hd__dfrtp_1
X_649_ _652_/A GND GND VDD VDD _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_673 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2698 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2529 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1541 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_109 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1430 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2017 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_503_ _726_/Q _725_/Q _503_/S GND GND VDD VDD _504_/A sky130_fd_sc_hd__mux2_1
X_434_ _757_/Q _756_/Q _436_/S GND GND VDD VDD _435_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1227 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_365_ _788_/Q _787_/Q _369_/S GND GND VDD VDD _366_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_3241 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_2849 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_893 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1861 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_2129 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3201 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_2741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2544 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1810 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1843 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_18_993 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1794 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2337 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1973 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_429 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1525 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1113 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_889 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_333 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_417_ _765_/Q _764_/Q _425_/S GND GND VDD VDD _418_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_2613 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_348_ _516_/A GND GND VDD VDD _393_/A sky130_fd_sc_hd__buf_4
XFILLER_18_1068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_3093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1225 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1269 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2396 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1684 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1789 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_14_2101 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_421 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_498 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_14_1477 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3161 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_837 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_749 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_15_237 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3277 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3280 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2465 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1617 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_6_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_8_2909 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1033 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1077 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2265 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clk clkbuf_0_clk/X GND GND VDD VDD _791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_1105 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1285 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1149 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_601 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_751_ _775_/CLK _751_/D _642_/Y GND GND VDD VDD _751_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2121 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_1729 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_5_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_682_ _683_/A GND GND VDD VDD _682_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_513 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_557 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1130 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_2785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2605 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2373 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_973 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_3_461 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3217 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1561 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_11_1425 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1469 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2717 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2485 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2073 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_505 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2037 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2925 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2969 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1093 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_74 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_921 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_965 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1537 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_734_ _773_/CLK _734_/D _620_/Y GND GND VDD VDD _734_/Q sky130_fd_sc_hd__dfrtp_1
X_665_ _665_/A GND GND VDD VDD _690_/A sky130_fd_sc_hd__buf_4
XFILLER_17_844 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_596_ _596_/A GND GND VDD VDD _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_16_343 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_365 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1701 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_3 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_12_1745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_65 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_2181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1789 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_781 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_181 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_19 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_17_3025 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1681 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1233 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1813 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_450_ _750_/Q _749_/Q _458_/S GND GND VDD VDD _451_/A sky130_fd_sc_hd__mux2_1
X_381_ _381_/A GND GND VDD VDD _781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_825 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_869 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_317 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput5 _785_/Q GND GND VDD VDD COL_SEL[10] sky130_fd_sc_hd__clkbuf_1
Xoutput40 _717_/Q GND GND VDD VDD COL_SEL[42] sky130_fd_sc_hd__clkbuf_1
Xoutput51 _727_/Q GND GND VDD VDD COL_SEL[52] sky130_fd_sc_hd__clkbuf_1
Xoutput62 _737_/Q GND GND VDD VDD COL_SEL[62] sky130_fd_sc_hd__clkbuf_1
Xoutput73 _747_/Q GND GND VDD VDD COL_SEL[72] sky130_fd_sc_hd__clkbuf_1
Xoutput84 _757_/Q GND GND VDD VDD COL_SEL[82] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput95 _767_/Q GND GND VDD VDD COL_SEL[92] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_2737 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_717_ _791_/CLK _717_/D _599_/Y GND GND VDD VDD _717_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_641 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_648_ _652_/A GND GND VDD VDD _648_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_685 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_579_ _597_/A GND GND VDD VDD _584_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1553 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2801 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1597 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_2165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1442 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2029 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_309 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_3045 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1621 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_1665 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_416 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_502_ _502_/A GND GND VDD VDD _727_/D sky130_fd_sc_hd__clkbuf_1
X_433_ _433_/A GND GND VDD VDD _758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_364_ _364_/A GND GND VDD VDD _789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_861 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3297 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1873 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2753 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_1833 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2305 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2349 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1941 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1985 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1537 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_19_1548 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1261 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_629 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2894 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_12_53 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1169 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_12_97 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_389 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_953 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_416_ _449_/A GND GND VDD VDD _425_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_2625 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2669 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_1681 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_5_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_20_3065 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2353 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_3137 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_2293 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_2113 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1592 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_20_444 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_14_2157 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1309 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3173 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_205 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1301 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2981 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_249 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1345 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_2068 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_905 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2989 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2809 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1080 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_949 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_1821 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_665 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_153 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_197 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2881 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_566 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1009 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_3292 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_15_2433 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2477 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1001 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_1045 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_1089 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_1565 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_13_709 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_241 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_14_1253 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_1117 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1297 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_613 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_7_2409 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_750_ _775_/CLK _750_/D _640_/Y GND GND VDD VDD _750_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_657 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_2177 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_681_ _683_/A GND GND VDD VDD _681_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_525 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_18_85 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_569 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_19_1142 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2742 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_713 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_2617 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2797 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_757 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_10_3053 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_473 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_1229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1841 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_17_3229 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1885 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1805 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_1849 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_2241 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1437 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3121 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_2729 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3165 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2317 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2041 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1373 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_2085 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_517 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2937 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_14_1061 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_20 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_20_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_20_97 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_421 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_933 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1505 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_1_977 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_20_2908 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_7_1549 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_733_ _775_/CLK _733_/D _619_/Y GND GND VDD VDD _733_/Q sky130_fd_sc_hd__dfrtp_1
X_664_ _664_/A GND GND VDD VDD _664_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_856 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_595_ _596_/A GND GND VDD VDD _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_355 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_16_377 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_2561 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1757 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XANTENNA_4 input1/X GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_6_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_10_2193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_281 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_793 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3305 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_1037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_3073 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_19_193 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_3037 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_1693 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1201 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_15_1381 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1245 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_11_1289 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_2261 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_8_1869 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_2_2125 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_2169 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_380_ _781_/Q _780_/Q _380_/S GND GND VDD VDD _381_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_837 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_1101 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_13_347 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_13_2701 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_13_2745 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput6 _786_/Q GND GND VDD VDD COL_SEL[11] sky130_fd_sc_hd__clkbuf_1
Xoutput30 _708_/Q GND GND VDD VDD COL_SEL[33] sky130_fd_sc_hd__clkbuf_1
Xoutput41 _718_/Q GND GND VDD VDD COL_SEL[43] sky130_fd_sc_hd__clkbuf_1
Xoutput52 _728_/Q GND GND VDD VDD COL_SEL[53] sky130_fd_sc_hd__clkbuf_1
Xoutput63 _738_/Q GND GND VDD VDD COL_SEL[63] sky130_fd_sc_hd__clkbuf_1
Xoutput74 _748_/Q GND GND VDD VDD COL_SEL[73] sky130_fd_sc_hd__clkbuf_1
Xoutput85 _758_/Q GND GND VDD VDD COL_SEL[83] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_741 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput96 _768_/Q GND GND VDD VDD COL_SEL[93] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_785 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1313 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_7_1357 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_716_ _786_/CLK _716_/D _598_/Y GND GND VDD VDD _716_/Q sky130_fd_sc_hd__dfrtp_1
X_647_ _659_/A GND GND VDD VDD _652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_653 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_16_141 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_578_ _578_/A GND GND VDD VDD _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2645 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_17_697 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_18_1955 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_841 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1521 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_12_1565 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2813 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_2857 GND VDD VDD GND sky130_ef_sc_hd__decap_12
.ends

.subckt pixel_fill gring VDD GND VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT CSA_VREF
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=7.5 as=24.809025 ps=56.34 w=2 l=1.44
X1 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.995 ps=8.8 w=1 l=0.8
X2 a_5720_n730# a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.25 pd=1.5 as=0.35 ps=2.7 w=1 l=1
X3 a_4330_n30# a_3852_n32# a_3852_n32# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.23 pd=1.65 as=0.3927 ps=2.8 w=1 l=2
X4 VDD SF_IB a_5720_n730# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.25 ps=1.5 w=1 l=1
X5 a_5460_10# a_4330_n30# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X6 a_3852_n32# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.76 ps=8.8 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=1
X8 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=1.995 pd=8.8 as=1.4 ps=7.4 w=7 l=0.15
X9 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.119375 pd=7.15 as=0 ps=0 w=2 l=3.35
X10 a_4120_n520# a_3852_n32# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X11 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=3.1 as=0.42 ps=3.1 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=2.95 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# VREF a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=1.4 pd=7.4 as=1.76 ps=8.8 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1.15
X16 VDD a_4330_n30# a_4330_n30# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.23 ps=1.65 w=1 l=2
X17 VDD a_5720_n730# a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.6 ps=2.95 w=1 l=0.15
X18 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X19 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=10.715 pd=15.9 as=0 ps=0 w=2.6 l=0.35
.ends

.subckt marker_pixel gring VDD GND VREF ROW_SEL NB1 VBIAS NB2 AMP_IN SF_IB PIX_OUT
+ CSA_VREF
X0 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.5 pd=7.5 as=24.809025 ps=56.34 w=2 l=1.44
X1 a_4120_n520# VBIAS a_4120_n750# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.995 ps=8.8 w=1 l=0.8
X2 a_5720_n730# a_4600_n810# GND VDD sky130_fd_pr__pfet_01v8_lvt ad=0.25 pd=1.5 as=0.35 ps=2.7 w=1 l=1
X3 a_4330_n30# a_3852_n32# a_3852_n32# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.23 pd=1.65 as=0.3927 ps=2.8 w=1 l=2
X4 VDD SF_IB a_5720_n730# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.25 ps=1.5 w=1 l=1
X5 a_5460_10# a_4330_n30# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.175 pd=1.35 as=0.35 ps=2.7 w=1 l=2
X6 a_3852_n32# VBIAS a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=1.76 ps=8.8 w=1 l=0.8
X7 VDD a_4120_n520# a_4600_n810# GND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=1
X8 a_4120_n750# AMP_IN a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=1.995 pd=8.8 as=1.4 ps=7.4 w=7 l=0.15
X9 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=3.119375 pd=7.15 as=0 ps=0 w=2 l=3.35
X10 a_4120_n520# a_3852_n32# a_5460_10# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.175 ps=1.35 w=1 l=2
X11 AMP_IN a_4600_n810# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GND NB1 a_4050_n2590# GND sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=3.1 as=0.42 ps=3.1 w=1.2 l=1
X13 a_5750_n920# ROW_SEL PIX_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=2.95 as=5.4 ps=9.4 w=2 l=1
X14 a_4050_n2590# a_4020_n2270# a_3860_n1150# GND sky130_fd_pr__nfet_01v8_lvt ad=1.4 pd=7.4 as=1.76 ps=8.8 w=7 l=0.15
X15 a_4600_n810# NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1.15
X16 VDD a_4330_n30# a_4330_n30# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.35 pd=2.7 as=0.23 ps=1.65 w=1 l=2
X17 VDD a_5720_n730# a_5750_n920# GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.6 ps=2.95 w=1 l=0.15
X18 AMP_IN CSA_VREF a_4600_n810# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.294 pd=2.24 as=0.273 ps=2.14 w=0.42 l=8
X19 GND GND GND GND sky130_fd_pr__nfet_01v8_lvt ad=10.715 pd=15.9 as=0 ps=0 w=2.6 l=0.35
.ends

.subckt pixel_array100x100_fill VBIAS VREF NB2 VDD NB1 ROW_SEL[0] GRING ROW_SEL[1]
+ ROW_SEL[2] ROW_SEL[3] ROW_SEL[4] ROW_SEL[5] ROW_SEL[6] ROW_SEL[7] ROW_SEL[8] ROW_SEL[9]
+ ROW_SEL[10] ROW_SEL[11] ROW_SEL[12] ROW_SEL[13] ROW_SEL[14] ROW_SEL[15] ROW_SEL[16]
+ ROW_SEL[17] ROW_SEL[18] ROW_SEL[19] ROW_SEL[20] ROW_SEL[21] ROW_SEL[22] ROW_SEL[23]
+ ROW_SEL[24] ROW_SEL[25] ROW_SEL[26] ROW_SEL[27] ROW_SEL[28] ROW_SEL[29] ROW_SEL[30]
+ ROW_SEL[31] ROW_SEL[32] ROW_SEL[33] ROW_SEL[34] ROW_SEL[35] ROW_SEL[36] ROW_SEL[37]
+ ROW_SEL[38] ROW_SEL[39] ROW_SEL[40] ROW_SEL[41] ROW_SEL[42] ROW_SEL[43] ROW_SEL[44]
+ ROW_SEL[45] ROW_SEL[46] ROW_SEL[47] ROW_SEL[48] ROW_SEL[49] ROW_SEL[50] ROW_SEL[51]
+ ROW_SEL[52] ROW_SEL[53] ROW_SEL[54] ROW_SEL[55] ROW_SEL[56] ROW_SEL[57] ROW_SEL[58]
+ ROW_SEL[59] ROW_SEL[60] ROW_SEL[61] ROW_SEL[62] ROW_SEL[63] ROW_SEL[64] ROW_SEL[65]
+ ROW_SEL[66] ROW_SEL[67] ROW_SEL[68] ROW_SEL[69] ROW_SEL[70] ROW_SEL[71] ROW_SEL[72]
+ ROW_SEL[73] ROW_SEL[74] ROW_SEL[75] ROW_SEL[76] ROW_SEL[77] ROW_SEL[78] ROW_SEL[79]
+ ROW_SEL[80] ROW_SEL[81] ROW_SEL[82] ROW_SEL[83] ROW_SEL[84] ROW_SEL[85] ROW_SEL[86]
+ ROW_SEL[87] ROW_SEL[88] ROW_SEL[89] ROW_SEL[90] ROW_SEL[91] ROW_SEL[92] ROW_SEL[93]
+ ROW_SEL[94] ROW_SEL[95] ROW_SEL[96] ROW_SEL[97] ROW_SEL[98] COL_SEL[0] CSA_VREF
+ ROW_SEL[99] COL_SEL[1] COL_SEL[2] COL_SEL[3] COL_SEL[4] COL_SEL[5] COL_SEL[6] COL_SEL[7]
+ COL_SEL[8] COL_SEL[9] COL_SEL[10] COL_SEL[11] COL_SEL[12] COL_SEL[13] COL_SEL[14]
+ COL_SEL[15] COL_SEL[16] COL_SEL[17] COL_SEL[18] COL_SEL[19] COL_SEL[20] COL_SEL[21]
+ COL_SEL[22] COL_SEL[23] COL_SEL[24] COL_SEL[25] COL_SEL[26] COL_SEL[27] COL_SEL[28]
+ COL_SEL[29] COL_SEL[30] COL_SEL[31] COL_SEL[32] COL_SEL[33] COL_SEL[34] COL_SEL[35]
+ COL_SEL[36] COL_SEL[37] COL_SEL[38] COL_SEL[39] COL_SEL[40] COL_SEL[41] COL_SEL[42]
+ COL_SEL[43] COL_SEL[44] COL_SEL[45] COL_SEL[46] COL_SEL[47] COL_SEL[48] COL_SEL[49]
+ COL_SEL[50] COL_SEL[51] COL_SEL[52] COL_SEL[53] COL_SEL[54] COL_SEL[55] COL_SEL[56]
+ COL_SEL[57] COL_SEL[58] COL_SEL[59] COL_SEL[60] COL_SEL[61] COL_SEL[62] COL_SEL[63]
+ COL_SEL[64] COL_SEL[65] COL_SEL[66] COL_SEL[67] COL_SEL[68] COL_SEL[69] COL_SEL[70]
+ COL_SEL[71] COL_SEL[72] COL_SEL[73] COL_SEL[74] COL_SEL[75] COL_SEL[76] COL_SEL[77]
+ COL_SEL[78] COL_SEL[79] COL_SEL[80] COL_SEL[81] COL_SEL[82] COL_SEL[83] COL_SEL[84]
+ COL_SEL[85] COL_SEL[86] COL_SEL[87] COL_SEL[88] COL_SEL[89] COL_SEL[90] COL_SEL[91]
+ COL_SEL[92] COL_SEL[93] COL_SEL[94] COL_SEL[95] COL_SEL[96] COL_SEL[97] COL_SEL[98]
+ ARRAY_OUT COL_SEL[99] SF_IB GND
Xpixel_fill_8909 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_305 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_316 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_327 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_338 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_349 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3205 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3216 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3227 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3238 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2504 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2515 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2526 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3249 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1803 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1814 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1825 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2537 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2548 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2559 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1836 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1847 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1858 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1869 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5130 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_883 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_872 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_861 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_850 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5141 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5152 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5163 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_894 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4440 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4451 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4462 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5174 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5185 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5196 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3750 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4473 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4484 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4495 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3761 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3772 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3783 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3794 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9418 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9407 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9429 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8717 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8706 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8739 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8728 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_102 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_113 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_124 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_135 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_146 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_157 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_168 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_179 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3002 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3013 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2301 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3024 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3035 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3046 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1600 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2312 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2323 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2334 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2345 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3057 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3068 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3079 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1611 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1622 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1633 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2356 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2367 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2378 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1644 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1655 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1666 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2389 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1677 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1688 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1699 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9941 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9930 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9974 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9963 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9952 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9996 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9985 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_691 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_680 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4270 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4281 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4292 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3580 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3591 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2890 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9237 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9226 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9215 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9204 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9259 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9248 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8525 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8514 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8503 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8558 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8547 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8536 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7824 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7813 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7802 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8569 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7857 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7846 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7835 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7879 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7868 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2120 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2131 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2142 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2153 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1441 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1430 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2164 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2175 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2186 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1474 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1463 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1452 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2197 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1496 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1485 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9782 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9771 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9760 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9793 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7109 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6408 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6419 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5707 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5718 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5729 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9012 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9001 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9045 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9034 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9023 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8300 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9078 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9067 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9056 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8333 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8322 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8311 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9089 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8377 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8366 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8355 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8344 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7632 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7621 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7610 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8399 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8388 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7665 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7654 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7643 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6920 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7698 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7687 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7676 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6953 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6942 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6931 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6997 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6986 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6975 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6964 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1293 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1282 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1271 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1260 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9590 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6216 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6205 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6249 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6238 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6227 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5504 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4803 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5515 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5526 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5537 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5548 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4814 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4825 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4836 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5559 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4847 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4858 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4869 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8141 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8130 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8185 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8174 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8163 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8152 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7440 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8196 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7473 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7462 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7451 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7495 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7484 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6772 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6761 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6750 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6794 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6783 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1090 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_509 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3409 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2708 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2719 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6002 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6013 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6024 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5301 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5312 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6035 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6046 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6057 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4600 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4611 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5323 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5334 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5345 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5356 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6068 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6079 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4622 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4633 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4644 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5367 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5378 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5389 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3910 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3921 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3932 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3943 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4655 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4666 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4677 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4688 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3954 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3965 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3976 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4699 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3987 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3998 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7281 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7270 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7292 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6580 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6591 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5890 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_306 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_317 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_328 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_339 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3206 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3217 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3228 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2505 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2516 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2527 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3239 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1804 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1815 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2538 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2549 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1826 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1837 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1848 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1859 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_840 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5120 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5131 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_873 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_862 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_851 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5142 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5153 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5164 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_895 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_884 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4430 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4441 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4452 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5175 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5186 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5197 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3740 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3751 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4463 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4474 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4485 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4496 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3762 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3773 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3784 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3795 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9419 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9408 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8707 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8729 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8718 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_103 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_114 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_125 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_136 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_147 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_158 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_169 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3003 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2302 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3014 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3025 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3036 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3047 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2313 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2324 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2335 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3058 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3069 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1601 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1612 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1623 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2346 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2357 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2368 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1634 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1645 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1656 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1667 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2379 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1678 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1689 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9931 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9920 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9975 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9964 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9953 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9942 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9997 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9986 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_681 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_670 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_692 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4260 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4271 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4282 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4293 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3570 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3581 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3592 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2880 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2891 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9227 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9216 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9205 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9249 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9238 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8526 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8515 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8504 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8559 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8548 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8537 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7814 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7803 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7847 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7836 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7825 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7869 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7858 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2110 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2121 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2132 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2143 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1442 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1431 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1420 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2154 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2165 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2176 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2187 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1475 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1464 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1453 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2198 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1497 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1486 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9750 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9783 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9772 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9761 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9794 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4090 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6409 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5708 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5719 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9002 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9035 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9024 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9013 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9079 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9068 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9057 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9046 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8334 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8323 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8312 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8301 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8367 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8356 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8345 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7622 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7611 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7600 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8389 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8378 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7666 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7655 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7644 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7633 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6921 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6910 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7699 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7688 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7677 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6954 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6943 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6932 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6987 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6976 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6965 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6998 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1250 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1283 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1272 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1261 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1294 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9591 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9580 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8890 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6206 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6239 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6228 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6217 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5505 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5516 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5527 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5538 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4804 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4815 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4826 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4837 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5549 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4848 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4859 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8142 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8131 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8120 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8175 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8164 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8153 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7430 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8197 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8186 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7474 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7463 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7452 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7441 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7496 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7485 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6762 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6751 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6740 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6795 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6784 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6773 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1091 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1080 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2709 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6003 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6014 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6025 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5302 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5313 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6036 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6047 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6058 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4601 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5324 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5335 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5346 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6069 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3900 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4612 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4623 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4634 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4645 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5357 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5368 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5379 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3911 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3922 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3933 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4656 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4667 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4678 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3944 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3955 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3966 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4689 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3977 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3988 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3999 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7282 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7271 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7260 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7293 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6570 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6592 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6581 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5880 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5891 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_307 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_318 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_329 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3207 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3218 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3229 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2506 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2517 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1805 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1816 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2528 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2539 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1827 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1838 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1849 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_830 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5110 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5121 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_874 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_863 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_852 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_841 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4420 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5132 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5143 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5154 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_896 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_885 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4431 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4442 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4453 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5165 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5176 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5187 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5198 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3730 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3741 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4464 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4475 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4486 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3752 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3763 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3774 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3785 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4497 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3796 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7090 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9409 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8708 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8719 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_104 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_115 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_126 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_137 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_148 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_159 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3004 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3015 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3026 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3037 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2303 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2314 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2325 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2336 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3048 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3059 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1602 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1613 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1624 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2347 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2358 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2369 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1635 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1646 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1657 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1668 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1679 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9932 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9921 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9910 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9965 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9954 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9943 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9998 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9987 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9976 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_682 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_671 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_660 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_693 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4250 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4261 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3560 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4272 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4283 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4294 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3571 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3582 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3593 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2870 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2881 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2892 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9228 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9217 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9206 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9239 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8516 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8505 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8549 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8538 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8527 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7804 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7848 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7837 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7826 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7815 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7859 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2100 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2111 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2122 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2133 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2144 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1432 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1421 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1410 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2155 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2166 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2177 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1465 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1454 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1443 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2188 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2199 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1498 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1487 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1476 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9740 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9773 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9762 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9751 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9795 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9784 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_490 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4080 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4091 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3390 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5709 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9003 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9036 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9025 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9014 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9069 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9058 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9047 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8324 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8313 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8302 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8368 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8357 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8346 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8335 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7623 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7612 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7601 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8379 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7656 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7645 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7634 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6911 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6900 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7689 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7678 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7667 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6944 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6933 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6922 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6988 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6977 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6966 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6955 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6999 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1240 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1284 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1273 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1262 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1251 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1295 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9592 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9581 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9570 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8880 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8891 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6207 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6229 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6218 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5506 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5517 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5528 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5539 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4805 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4816 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4827 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4838 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4849 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8132 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8121 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8110 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8176 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8165 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8154 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8143 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7431 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7420 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8198 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8187 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7464 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7453 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7442 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7497 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7486 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7475 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6763 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6752 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6741 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6730 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6796 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6785 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6774 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1092 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1081 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1070 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6004 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6015 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5303 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6026 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6037 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6048 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4602 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5314 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5325 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5336 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5347 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6059 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4613 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4624 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4635 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5358 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5369 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3901 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3912 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3923 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3934 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4646 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4657 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4668 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4679 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3945 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3956 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3967 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3978 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3989 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7272 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7261 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7250 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7294 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7283 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6571 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6560 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6593 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6582 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5870 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5881 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5892 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_308 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_319 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3208 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3219 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2507 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2518 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1806 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2529 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1817 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1828 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1839 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_831 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_820 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5100 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5111 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5122 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_864 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_853 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_842 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4410 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5133 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5144 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5155 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_897 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_886 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_875 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4421 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4432 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4443 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5166 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5177 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5188 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3720 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3731 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3742 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4454 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4465 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4476 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4487 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5199 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3753 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3764 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3775 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4498 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3786 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3797 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7091 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7080 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6390 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8709 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_105 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_116 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_127 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_138 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_149 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3005 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3016 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3027 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3038 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2304 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2315 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2326 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3049 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1603 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1614 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2337 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2348 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2359 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1625 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1636 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1647 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1658 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1669 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9922 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9911 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9900 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9966 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9955 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9944 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9933 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9999 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9988 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9977 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_672 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_661 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_650 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_694 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_683 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4240 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4251 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4262 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3550 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4273 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4284 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4295 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3561 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3572 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3583 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2860 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2871 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2882 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3594 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2893 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9218 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9207 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9229 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8517 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8506 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8539 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8528 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7805 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7838 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7827 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7816 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7849 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2101 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2112 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2123 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2134 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1433 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1422 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1411 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1400 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2145 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2156 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2167 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1466 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1455 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1444 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2178 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2189 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1499 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1488 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1477 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9741 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9730 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9774 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9763 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9752 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9796 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9785 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_491 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_480 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4070 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4081 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4092 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3380 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3391 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2690 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9026 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9015 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9004 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9059 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9048 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9037 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8325 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8314 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8303 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8358 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8347 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8336 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7613 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7602 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8369 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7646 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7635 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7624 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6912 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6901 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7679 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7668 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7657 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6945 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6934 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6923 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6978 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6967 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6956 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6989 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1241 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1230 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1274 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1263 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1252 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1296 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1285 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9582 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9571 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9560 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9593 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8881 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8870 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8892 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6219 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6208 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5507 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5518 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5529 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4806 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4817 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4828 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4839 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8100 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8133 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8122 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8111 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8166 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8155 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8144 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7421 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7410 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8199 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8188 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8177 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7465 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7454 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7443 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7432 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6720 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7498 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7487 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7476 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6753 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6742 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6731 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6786 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6775 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6764 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6797 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1082 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1071 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1060 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1093 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9390 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6005 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6016 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5304 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6027 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6038 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6049 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5315 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5326 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5337 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4603 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4614 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4625 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4636 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5348 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5359 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3902 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3913 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3924 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4647 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4658 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4669 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3935 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3946 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3957 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3968 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3979 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7240 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7273 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7262 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7251 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7295 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7284 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6561 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6550 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6594 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6583 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6572 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5860 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5871 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5882 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5893 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_309 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3209 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2508 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1807 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2519 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1818 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1829 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_821 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_810 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5101 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5112 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_865 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_854 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_843 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_832 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4400 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4411 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5123 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5134 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5145 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_898 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_887 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_876 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4422 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4433 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4444 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5156 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5167 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5178 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5189 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3710 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3721 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3732 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4455 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4466 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4477 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3743 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3754 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3765 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3776 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4488 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4499 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3787 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3798 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7081 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7070 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7092 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6380 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6391 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5690 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_106 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_117 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_128 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_139 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3006 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3017 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3028 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2305 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2316 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3039 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1604 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1615 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2327 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2338 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2349 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1626 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1637 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1648 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1659 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9923 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9912 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9901 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9956 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9945 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9934 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9989 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9978 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9967 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_640 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_673 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_662 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_651 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_695 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_684 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4230 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4241 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4252 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3540 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3551 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4263 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4274 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4285 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3562 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3573 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3584 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4296 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2850 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2861 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2872 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3595 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2883 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2894 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9219 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9208 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8507 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8529 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8518 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7839 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7828 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7817 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7806 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2102 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2113 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2124 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2135 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1423 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1412 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1401 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2146 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2157 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2168 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1456 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1445 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1434 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2179 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1489 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1478 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1467 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9731 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9720 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9764 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9753 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9742 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9797 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9786 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9775 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_481 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_470 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_492 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4060 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4071 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4082 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4093 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3370 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3381 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3392 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2680 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2691 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1990 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9027 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9016 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9005 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9049 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9038 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8315 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8304 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8359 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8348 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8337 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8326 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7614 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7603 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7647 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7636 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7625 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6902 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7669 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7658 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6935 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6924 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6913 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6979 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6968 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6957 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6946 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1231 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1220 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1275 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1264 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1253 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1242 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1297 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1286 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9583 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9572 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9561 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9550 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9594 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8871 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8860 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8893 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8882 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6209 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5508 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5519 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4807 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4818 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4829 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8123 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8112 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8101 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8167 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8156 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8145 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8134 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7422 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7411 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7400 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8189 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8178 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7455 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7444 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7433 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6710 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7488 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7477 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7466 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6754 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6743 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6732 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6721 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7499 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6787 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6776 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6765 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6798 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1050 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1083 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1072 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1061 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1094 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9391 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9380 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8690 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6006 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6017 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6028 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6039 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5305 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5316 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5327 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5338 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4604 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4615 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4626 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5349 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3903 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3914 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3925 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4637 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4648 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4659 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3936 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3947 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3958 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3969 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7230 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7263 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7252 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7241 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7296 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7285 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7274 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6562 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6551 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6540 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6595 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6584 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6573 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5850 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5861 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5872 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5883 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5894 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2509 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1808 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1819 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_822 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_811 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_800 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5102 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5113 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_855 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_844 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_833 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4401 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5124 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5135 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5146 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_899 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_888 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_877 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_866 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3700 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4412 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4423 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4434 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5157 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5168 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5179 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3711 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3722 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3733 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4445 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4456 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4467 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4478 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3744 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3755 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3766 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4489 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3777 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3788 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3799 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7082 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7071 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7060 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7093 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6370 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6392 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6381 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5680 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5691 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4990 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_107 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_118 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_129 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3007 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3018 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3029 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2306 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2317 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1605 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2328 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2339 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1616 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1627 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1638 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1649 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9913 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9902 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9957 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9946 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9935 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9924 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9979 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9968 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_630 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_663 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_652 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_641 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_696 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_685 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_674 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4220 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4231 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4242 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4253 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3530 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3541 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4264 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4275 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4286 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2840 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3552 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3563 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3574 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4297 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2851 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2862 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2873 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3585 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3596 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2884 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2895 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9209 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8508 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8519 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7829 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7818 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7807 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2103 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2114 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2125 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1424 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1413 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1402 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2136 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2147 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2158 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1457 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1446 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1435 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2169 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1479 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1468 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9732 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9721 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9710 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9765 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9754 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9743 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9798 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9787 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9776 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_482 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_471 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_460 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_493 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4050 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4061 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4072 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4083 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4094 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3360 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3371 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3382 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3393 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2670 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2681 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2692 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1980 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1991 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9017 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9006 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9039 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9028 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8316 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8305 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8349 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8338 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8327 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7604 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7637 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7626 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7615 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6903 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7659 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7648 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6936 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6925 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6914 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6969 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6958 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6947 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1232 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1221 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1210 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1265 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1254 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1243 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1298 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1287 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1276 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9540 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9573 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9562 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9551 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9595 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9584 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8872 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8861 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8850 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8894 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8883 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_290 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3190 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5509 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4808 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4819 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8124 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8113 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8102 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8157 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8146 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8135 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7412 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7401 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8179 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8168 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7456 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7445 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7434 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7423 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6711 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6700 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7489 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7478 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7467 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6744 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6733 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6722 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6777 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6766 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6755 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6799 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6788 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1040 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1073 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1062 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1051 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1095 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1084 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9381 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9370 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9392 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8680 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8691 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7990 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6007 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6018 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6029 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5306 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5317 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5328 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4605 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4616 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4627 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5339 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3904 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3915 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4638 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4649 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3926 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3937 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3948 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3959 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7231 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7220 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7264 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7253 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7242 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7297 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7286 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7275 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6552 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6541 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6530 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6596 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6585 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6574 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6563 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5840 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5851 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5862 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5873 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5884 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5895 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1809 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_812 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_801 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5103 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_856 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_845 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_834 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_823 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4402 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5114 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5125 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5136 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_889 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_878 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_867 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4413 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4424 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4435 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5147 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5158 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5169 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3701 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3712 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3723 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4446 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4457 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4468 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3734 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3745 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3756 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3767 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4479 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3778 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3789 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7072 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7061 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7050 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7094 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7083 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6371 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6360 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6393 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6382 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5670 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5681 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5692 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4980 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4991 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_108 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_119 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3008 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3019 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2307 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1606 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2318 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2329 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1617 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1628 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1639 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9914 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9903 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9947 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9936 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9925 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9969 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9958 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_631 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_620 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_664 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_653 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_642 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4210 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_697 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_686 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_675 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4221 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4232 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4243 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3520 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3531 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3542 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4254 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4265 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4276 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2830 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3553 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3564 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3575 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4287 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4298 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2841 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2852 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2863 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3586 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3597 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2874 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2885 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2896 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6190 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8509 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7819 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7808 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2104 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2115 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2126 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1414 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1403 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2137 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2148 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2159 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1447 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1436 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1425 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1469 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1458 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9722 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9711 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9700 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9755 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9744 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9733 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9799 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9788 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9777 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9766 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_472 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_461 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_450 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_494 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_483 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4040 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4051 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3350 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4062 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4073 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4084 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4095 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3361 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3372 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3383 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2660 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2671 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2682 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3394 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1970 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2693 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1981 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1992 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9018 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9007 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9029 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8306 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8339 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8328 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8317 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7605 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7638 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7627 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7616 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7649 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6926 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6915 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6904 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6959 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6948 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6937 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1222 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1211 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1200 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1266 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1255 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1244 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1233 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1299 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1288 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1277 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9530 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9574 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9563 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9552 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9541 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9596 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9585 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8862 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8851 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8840 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8895 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8884 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8873 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_280 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_291 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3180 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3191 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2490 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4809 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8114 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8103 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8158 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8147 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8136 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8125 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7413 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7402 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8169 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7446 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7435 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7424 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6701 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7479 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7468 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7457 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6745 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6734 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6723 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6712 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6778 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6767 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6756 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6789 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1041 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1030 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1074 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1063 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1052 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1096 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1085 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9382 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9371 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9360 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9393 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8670 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8692 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8681 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7991 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7980 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6008 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6019 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5307 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5318 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5329 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4606 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4617 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3905 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3916 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4628 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4639 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3927 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3938 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3949 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7221 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7210 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7254 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7243 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7232 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6520 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7298 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7287 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7276 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7265 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6553 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6542 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6531 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6586 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6575 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6564 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5830 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5841 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6597 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5852 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5863 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5874 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5885 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5896 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9190 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_813 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_802 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5104 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_846 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_835 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_824 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5115 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5126 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5137 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_879 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_868 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_857 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4403 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4414 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4425 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5148 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5159 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3702 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3713 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3724 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4436 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4447 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4458 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4469 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3735 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3746 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3757 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3768 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3779 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7073 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7062 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7051 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7040 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7095 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7084 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6361 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6350 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6394 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6383 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6372 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5660 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5671 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5682 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5693 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4970 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4981 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4992 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_109 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3009 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2308 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2319 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1607 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1618 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1629 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9904 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9948 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9937 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9926 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9915 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9959 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_621 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_610 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_654 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_643 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_632 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4200 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_698 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_687 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_676 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_665 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4211 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4222 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4233 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4244 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3510 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3521 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3532 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4255 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4266 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4277 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2820 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2831 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3543 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3554 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3565 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4288 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4299 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2842 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2853 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2864 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3576 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3587 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3598 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2875 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2886 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2897 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6191 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6180 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5490 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7809 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2105 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2116 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1415 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1404 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2127 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2138 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2149 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1448 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1437 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1426 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1459 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9723 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9712 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9701 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9756 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9745 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9734 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9789 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9778 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9767 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_473 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_462 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_451 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_440 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_495 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_484 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4030 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4041 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4052 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3340 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4063 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4074 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4085 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3351 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3362 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3373 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3384 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4096 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2650 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2661 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2672 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3395 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1960 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2683 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2694 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1971 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1982 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1993 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9008 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9019 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8307 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8329 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8318 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7628 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7617 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7606 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7639 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6927 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6916 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6905 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6949 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6938 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1223 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1212 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1201 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1256 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1245 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1234 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1289 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1278 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1267 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9531 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9520 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9564 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9553 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9542 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9597 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9586 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9575 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8863 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8852 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8841 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8830 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8896 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8885 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8874 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_270 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_281 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_292 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3170 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3181 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3192 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2480 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2491 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1790 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xmarker_pixel_0 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 marker_pixel_0/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF marker_pixel
Xpixel_fill_8115 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8104 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8148 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8137 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8126 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7403 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8159 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7447 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7436 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7425 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7414 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6702 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7469 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7458 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6735 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6724 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6713 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6768 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6757 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6746 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6779 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1031 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1020 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1064 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1053 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1042 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1097 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1086 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1075 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9372 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9361 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9350 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9394 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9383 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8671 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8660 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8693 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8682 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7992 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7981 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7970 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6009 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5308 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5319 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4607 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4618 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3906 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4629 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3917 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3928 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3939 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7222 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7211 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7200 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7255 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7244 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7233 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6510 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7288 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7277 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7266 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6543 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6532 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6521 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7299 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6587 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6576 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6565 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6554 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5820 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5831 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5842 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6598 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5853 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5864 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5875 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5886 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5897 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9191 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9180 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8490 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_803 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_847 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_836 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_825 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_814 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5105 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5116 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5127 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_869 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_858 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4404 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4415 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4426 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5138 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5149 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3703 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3714 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4437 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4448 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4459 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3725 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3736 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3747 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3758 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3769 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7030 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7063 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7052 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7041 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7096 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7085 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7074 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6362 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6351 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6340 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6395 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6384 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6373 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5650 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5661 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5672 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5683 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4960 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4971 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4982 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5694 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4993 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2309 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1608 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1619 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9905 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9938 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9927 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9916 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9949 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_622 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_611 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_600 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_655 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_644 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_633 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4201 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_688 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_677 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_666 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4212 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4223 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4234 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_699 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3500 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3511 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3522 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3533 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4245 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4256 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4267 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2810 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2821 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3544 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3555 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3566 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4278 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4289 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2832 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2843 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2854 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3577 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3588 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3599 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2865 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2876 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2887 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2898 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6170 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6192 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6181 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5480 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5491 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4790 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2106 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2117 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1405 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2128 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2139 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1438 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1427 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1416 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1449 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9713 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9702 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9746 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9735 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9724 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9779 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9768 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9757 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_430 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_463 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_452 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_441 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_496 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_485 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_474 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4020 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4031 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4042 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3330 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3341 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4053 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4064 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4075 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4086 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3352 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3363 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3374 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4097 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2640 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2651 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2662 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2673 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3385 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3396 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1950 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1961 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2684 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2695 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1972 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1983 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1994 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9009 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8319 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8308 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7629 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7618 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7607 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6917 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6906 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6939 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6928 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1213 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1202 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1257 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1246 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1235 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1224 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1279 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1268 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9521 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9510 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9565 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9554 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9543 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9532 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8820 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9598 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9587 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9576 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8853 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8842 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8831 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8886 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8875 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8864 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8897 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_260 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_271 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_282 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_293 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3160 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3171 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3182 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2470 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2481 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3193 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2492 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1780 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1791 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xmarker_pixel_1 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 marker_pixel_1/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF marker_pixel
Xpixel_fill_8105 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8149 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8138 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8127 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8116 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7404 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7437 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7426 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7415 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7459 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7448 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6736 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6725 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6714 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6703 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6769 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6758 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6747 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1032 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1021 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1010 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1065 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1054 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1043 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1098 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1087 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1076 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9340 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9373 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9362 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9351 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9395 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9384 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8661 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8650 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8694 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8683 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8672 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7960 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7993 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7982 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7971 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5309 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4608 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3907 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4619 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3918 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3929 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7212 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7201 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7245 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7234 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7223 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6511 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6500 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7289 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7278 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7267 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7256 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6544 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6533 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6522 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6577 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6566 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6555 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5810 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5821 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5832 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6599 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6588 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5843 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5854 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5865 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5876 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5887 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5898 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9181 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9170 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9192 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8491 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8480 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7790 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_804 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_837 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_826 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_815 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5106 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5117 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5128 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_859 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_848 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4405 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4416 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5139 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3704 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3715 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4427 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4438 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4449 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3726 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3737 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3748 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3759 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7020 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7064 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7053 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7042 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7031 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7097 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7086 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7075 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6352 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6341 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6330 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6385 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6374 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6363 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5640 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6396 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5651 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5662 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5673 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5684 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4950 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4961 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4972 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5695 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4983 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4994 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1609 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9939 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9928 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9917 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9906 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_612 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_601 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_645 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_634 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_623 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_689 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_678 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_667 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_656 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4202 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4213 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4224 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4235 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3501 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3512 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3523 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4246 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4257 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4268 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2800 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2811 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3534 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3545 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3556 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4279 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2822 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2833 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2844 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2855 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3567 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3578 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3589 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2866 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2877 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2888 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2899 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6160 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6193 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6182 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6171 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5470 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5481 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5492 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4780 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4791 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2107 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1406 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2118 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2129 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1439 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1428 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1417 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9714 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9703 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9747 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9736 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9725 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9769 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9758 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_420 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_464 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_453 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_442 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_431 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4010 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_497 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_486 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_475 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4021 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4032 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4043 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3320 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3331 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4054 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4065 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4076 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2630 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3342 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3353 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3364 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3375 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4087 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4098 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2641 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2652 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2663 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3386 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3397 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1940 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1951 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2674 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2685 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2696 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1962 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1973 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1984 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1995 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8309 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7619 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7608 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6918 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6907 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6929 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1214 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1203 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1247 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1236 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1225 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1269 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1258 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9522 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9511 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9500 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9555 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9544 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9533 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8810 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9588 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9577 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9566 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8854 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8843 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8832 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8821 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9599 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8887 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8876 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8865 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8898 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_250 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_261 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_272 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_283 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_294 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3150 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3161 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3172 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3183 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2460 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2471 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3194 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1770 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2482 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2493 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1781 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1792 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8106 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8139 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8128 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8117 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7438 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7427 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7416 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7405 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7449 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6726 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6715 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6704 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6759 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6748 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6737 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1022 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1011 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1000 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1055 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1044 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1033 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1099 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1088 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1077 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1066 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9330 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9363 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9352 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9341 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9396 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9385 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9374 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8662 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8651 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8640 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8695 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8684 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8673 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7950 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7983 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7972 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7961 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7994 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2290 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4609 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3908 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3919 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7213 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7202 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7246 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7235 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7224 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6501 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7279 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7268 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7257 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6534 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6523 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6512 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6578 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6567 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6556 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6545 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5800 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5811 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5822 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5833 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6589 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5844 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5855 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5866 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5877 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5888 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5899 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9182 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9171 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9160 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9193 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8470 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8492 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8481 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7791 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7780 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_838 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_827 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_816 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_805 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5107 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5118 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_849 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4406 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4417 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5129 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3705 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4428 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4439 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3716 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3727 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3738 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3749 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7021 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7010 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7054 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7043 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7032 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7087 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7076 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7065 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6353 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6342 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6331 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6320 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7098 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6386 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6375 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6364 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5630 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5641 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6397 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5652 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5663 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5674 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4940 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4951 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4962 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4973 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5685 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5696 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4984 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4995 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9929 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9918 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9907 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_613 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_602 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_646 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_635 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_624 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_679 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_668 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_657 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4203 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4214 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4225 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3502 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3513 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3524 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4236 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4247 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4258 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2801 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2812 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3535 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3546 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3557 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4269 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2823 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2834 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2845 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3568 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3579 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2856 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2867 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2878 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2889 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6161 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6150 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6194 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6183 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6172 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5460 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5471 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5482 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4770 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4781 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5493 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4792 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2108 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2119 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1429 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1418 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1407 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9704 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9737 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9726 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9715 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9759 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9748 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_421 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_410 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_454 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_443 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_432 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4000 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_487 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_476 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_465 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4011 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4022 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4033 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_498 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3310 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3321 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3332 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4044 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4055 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4066 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4077 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2620 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3343 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3354 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3365 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4088 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4099 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2631 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2642 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2653 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3376 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3387 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3398 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1930 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1941 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1952 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2664 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2675 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2686 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2697 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1963 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1974 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1985 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1996 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5290 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7609 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6908 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6919 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1204 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1248 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1237 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1226 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1215 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1259 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9512 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9501 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9556 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9545 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9534 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9523 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8811 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8800 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9589 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9578 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9567 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8844 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8833 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8822 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8877 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8866 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8855 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8899 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8888 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_240 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_251 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_262 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_273 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_284 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_295 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3140 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3151 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3162 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3173 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2450 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2461 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2472 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3184 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3195 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1760 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2483 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2494 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1771 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1782 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1793 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8129 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8118 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8107 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7428 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7417 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7406 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7439 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6727 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6716 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6705 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6749 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6738 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1023 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1012 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1001 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1056 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1045 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1034 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1089 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1078 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1067 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9331 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9320 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9364 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9353 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9342 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9397 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9386 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9375 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8652 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8641 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8630 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8696 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8685 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8674 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8663 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7951 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7940 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7984 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7973 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7962 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7995 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2280 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2291 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1590 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3909 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7203 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7236 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7225 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7214 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6502 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7269 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7258 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7247 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6535 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6524 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6513 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6568 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6557 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6546 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5801 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5812 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5823 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6579 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5834 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5845 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5856 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5867 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5878 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5889 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9172 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9161 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9150 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9194 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9183 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8460 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8493 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8482 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8471 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7792 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7781 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7770 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_828 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_817 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_806 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5108 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5119 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_839 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4407 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3706 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4418 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4429 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3717 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3728 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3739 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7011 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7000 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7055 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7044 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7033 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7022 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6310 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7088 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7077 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7066 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6343 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6332 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6321 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7099 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6376 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6365 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6354 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5620 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5631 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6398 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6387 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4930 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5642 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5653 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5664 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5675 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4941 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4952 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4963 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5686 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5697 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4974 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4985 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4996 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8290 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9919 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9908 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_603 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_636 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_625 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_614 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_669 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_658 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_647 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4204 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4215 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4226 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3503 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3514 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4237 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4248 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4259 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2802 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3525 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3536 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3547 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2813 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2824 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2835 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2846 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3558 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3569 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2857 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2868 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2879 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6151 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6140 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6195 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6184 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6173 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6162 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5450 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5461 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5472 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5483 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4760 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4771 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5494 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4782 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4793 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2109 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1419 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1408 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9705 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9738 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9727 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9716 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9749 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_411 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_400 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_455 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_444 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_433 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_422 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_488 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_477 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_466 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4001 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4012 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4023 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4034 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_499 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3300 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3311 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3322 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4045 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4056 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4067 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2610 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2621 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3333 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3344 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3355 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3366 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4078 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4089 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2632 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2643 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2654 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3377 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3388 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3399 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1920 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1931 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1942 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2665 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2676 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2687 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1953 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1964 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1975 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1986 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2698 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1997 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5280 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5291 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4590 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6909 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1205 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1238 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1227 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1216 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1249 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9513 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9502 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9546 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9535 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9524 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8801 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9579 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9568 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9557 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8845 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8834 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8823 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8812 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8878 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8867 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8856 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8889 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_230 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_241 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_252 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_263 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_274 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_285 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_296 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3130 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3141 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3152 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3163 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3174 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2440 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2451 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2462 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3185 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3196 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1750 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1761 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2473 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2484 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2495 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1772 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1783 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1794 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8119 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8108 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7429 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7418 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7407 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6717 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6706 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6739 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6728 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1013 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1002 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1046 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1035 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1024 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1079 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1068 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1057 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9321 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9310 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9354 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9343 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9332 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9398 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9387 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9376 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9365 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8653 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8642 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8631 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8620 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8686 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8675 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8664 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7941 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7930 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8697 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7974 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7963 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7952 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7996 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7985 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2270 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2281 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2292 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1580 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1591 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7204 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7237 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7226 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7215 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7259 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7248 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6525 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6514 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6503 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6569 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6558 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6547 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6536 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5802 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5813 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5824 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5835 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5846 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5857 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5868 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5879 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9173 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9162 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9151 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9140 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9195 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9184 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8461 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8450 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8494 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8483 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8472 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7793 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7782 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7771 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7760 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_829 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_818 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_807 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5109 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4408 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4419 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3707 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3718 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3729 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7012 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7001 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7045 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7034 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7023 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6300 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7078 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7067 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7056 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6344 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6333 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6322 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6311 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7089 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6377 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6366 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6355 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5610 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5621 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5632 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6399 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6388 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4920 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5643 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5654 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5665 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4931 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4942 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4953 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4964 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5676 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5687 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5698 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4975 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4986 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4997 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8291 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8280 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7590 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9909 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_604 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_637 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_626 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_615 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_659 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_648 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4205 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4216 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3504 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3515 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4227 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4238 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4249 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2803 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3526 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3537 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3548 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2814 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2825 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2836 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3559 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2847 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2858 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2869 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6152 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6130 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6141 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6185 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6174 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6163 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5440 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6196 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5451 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5462 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5473 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4750 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4761 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4772 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5484 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5495 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4783 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4794 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1409 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9728 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9717 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9706 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9739 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_412 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_401 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_445 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_434 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_423 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_478 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_467 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_456 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4002 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4013 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4024 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_489 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3301 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3312 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3323 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4035 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4046 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4057 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4068 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2600 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2611 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3334 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3345 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3356 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4079 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1910 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2622 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2633 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2644 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3367 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3378 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3389 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1921 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1932 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1943 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2655 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2666 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2677 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2688 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1954 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1965 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1976 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2699 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1987 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1998 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_990 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5270 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5281 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5292 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4580 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4591 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3890 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1239 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1228 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1217 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1206 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9503 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9547 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9536 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9525 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9514 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8802 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9569 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9558 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8835 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8824 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8813 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8868 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8857 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8846 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8879 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_220 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_231 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_242 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_253 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_264 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_275 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_286 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_297 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3120 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3131 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3142 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3153 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3164 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2430 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2441 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2452 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2463 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3175 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3186 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3197 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1740 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1751 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2474 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2485 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2496 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1762 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1773 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1784 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1795 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8109 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7419 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7408 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6718 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6707 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6729 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1014 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1003 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1047 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1036 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1025 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1069 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1058 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9311 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9300 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9355 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9344 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9333 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9322 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8610 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9388 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9377 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9366 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8643 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8632 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8621 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9399 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8687 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8676 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8665 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8654 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7942 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7931 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7920 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8698 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7975 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7964 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7953 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7997 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7986 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2260 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2271 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2282 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2293 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1570 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1581 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1592 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7227 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7216 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7205 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7249 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7238 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6526 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6515 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6504 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6559 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6548 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6537 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5803 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5814 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5825 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5836 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5847 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5858 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5869 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9130 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9163 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9152 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9141 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9196 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9185 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9174 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8451 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8440 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8495 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8484 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8473 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8462 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7750 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7783 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7772 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7761 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7794 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2090 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_819 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_808 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4409 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3708 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3719 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7002 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7046 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7035 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7024 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7013 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6301 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7079 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7068 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7057 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6334 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6323 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6312 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6367 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6356 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6345 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5600 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5611 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5622 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6389 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6378 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4910 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4921 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5633 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5644 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5655 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5666 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4932 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4943 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4954 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5677 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5688 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5699 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4965 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4976 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4987 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4998 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8270 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8292 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8281 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7591 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7580 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6890 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_627 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_616 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_605 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_649 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_638 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4206 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4217 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3505 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4228 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4239 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3516 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3527 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3538 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2804 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2815 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2826 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2837 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3549 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2848 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2859 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6120 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6131 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6142 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6186 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6175 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6164 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6153 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5430 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5441 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6197 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5452 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5463 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5474 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4740 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4751 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4762 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5485 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5496 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4773 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4784 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4795 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9729 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9718 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9707 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_402 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_446 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_435 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_424 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_413 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_479 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_468 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_457 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4003 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4014 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4025 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3302 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3313 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4036 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4047 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4058 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2601 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2612 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3324 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3335 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3346 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3357 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4069 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1900 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2623 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2634 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2645 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3368 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3379 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1911 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1922 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1933 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2656 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2667 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2678 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1944 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1955 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1966 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1977 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2689 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1988 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1999 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_991 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_980 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5260 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5271 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5282 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4570 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4581 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5293 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4592 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3880 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3891 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1229 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1218 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1207 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9504 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9537 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9526 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9515 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9559 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9548 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8836 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8825 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8814 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8803 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8869 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8858 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8847 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_210 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_221 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_232 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_243 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_254 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_265 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_276 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_287 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_298 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3110 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3121 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2420 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3132 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3143 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3154 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3165 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2431 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2442 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2453 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3176 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3187 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3198 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1730 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1741 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1752 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2464 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2475 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2486 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1763 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1774 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1785 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2497 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1796 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5090 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7409 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6708 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6719 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1004 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1037 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1026 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1015 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1059 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1048 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9312 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9301 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9345 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9334 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9323 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8600 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9389 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9378 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9367 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9356 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8644 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8633 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8622 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8611 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8677 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8666 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8655 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7932 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7921 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7910 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8699 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8688 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7965 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7954 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7943 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7998 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7987 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7976 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2250 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2261 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1560 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2272 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2283 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2294 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1571 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1582 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1593 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9890 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7228 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7217 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7206 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7239 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6516 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6505 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6549 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6538 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6527 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5804 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5815 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5826 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5837 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5848 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5859 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9120 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9153 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9142 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9131 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9197 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9186 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9175 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9164 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8452 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8441 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8430 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8485 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8474 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8463 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7740 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8496 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7784 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7773 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7762 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7751 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7795 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2080 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2091 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1390 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_809 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3709 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7003 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7036 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7025 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7014 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7069 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7058 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7047 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6335 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6324 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6313 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6302 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6368 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6357 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6346 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5601 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5612 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5623 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6379 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4900 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4911 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5634 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5645 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5656 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4922 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4933 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4944 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4955 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5667 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5678 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5689 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4966 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4977 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4988 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4999 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8260 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8293 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8282 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8271 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7592 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7581 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7570 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6880 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6891 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_628 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_617 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_606 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_639 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4207 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3506 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4218 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4229 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3517 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3528 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3539 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2805 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2816 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2827 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2838 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2849 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6110 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6121 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6132 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6143 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6176 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6165 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6154 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5420 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5431 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6198 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6187 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4730 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5442 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5453 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5464 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4741 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4752 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4763 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5475 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5486 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5497 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4774 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4785 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4796 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8090 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9719 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9708 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_403 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_436 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_425 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_414 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_2/AMP_IN SF_IB
+ pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_469 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_458 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_447 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4004 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4015 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3303 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3314 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4026 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4037 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4048 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4059 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2602 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3325 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3336 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3347 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1901 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2613 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2624 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2635 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3358 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3369 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1912 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1923 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1934 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2646 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2657 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2668 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2679 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1945 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1956 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1967 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1978 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1989 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_992 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_981 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_970 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5250 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5261 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5272 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5283 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4560 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4571 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5294 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3870 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4582 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4593 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3881 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3892 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1219 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1208 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9538 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9527 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9516 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9505 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9549 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8826 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8815 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8804 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8859 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8848 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8837 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_200 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_211 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_222 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_233 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_244 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_255 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_266 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_277 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_288 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_299 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3100 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3111 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3122 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2410 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3133 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3144 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3155 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2421 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2432 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2443 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2454 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3166 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3177 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3188 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3199 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1720 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1731 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1742 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2465 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2476 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2487 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1753 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1764 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1775 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2498 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1786 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1797 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5080 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5091 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4390 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6709 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1005 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1038 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1027 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1016 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1049 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9302 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9346 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9335 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9324 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9313 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8601 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9379 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9368 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9357 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8634 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8623 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8612 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8678 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8667 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8656 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8645 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7933 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7922 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7911 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7900 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8689 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7966 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7955 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7944 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7999 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7988 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7977 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2240 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2251 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2262 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1550 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2273 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2284 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2295 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1561 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1572 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1583 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1594 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9891 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9880 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7218 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7207 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7229 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6517 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6506 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6539 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6528 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5805 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5816 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5827 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5838 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5849 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9121 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9110 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9154 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9143 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9132 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9187 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9176 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9165 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8442 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8431 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8420 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9198 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8486 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8475 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8464 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8453 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7741 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7730 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8497 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7774 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7763 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7752 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7796 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7785 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2070 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2081 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2092 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1391 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1380 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7037 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7026 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7015 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7004 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7059 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7048 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6325 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6314 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6303 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6358 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6347 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6336 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5602 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5613 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6369 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4901 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4912 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5624 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5635 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5646 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5657 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4923 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4934 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4945 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5668 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5679 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4956 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4967 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4978 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4989 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8261 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8250 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8294 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8283 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8272 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7582 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7571 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7560 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7593 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6881 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6870 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6892 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_618 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_607 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_629 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4208 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4219 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3507 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3518 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3529 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2806 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2817 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2828 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2839 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6100 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6111 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6122 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6133 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6177 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6166 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6155 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5410 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5421 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5432 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6144 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6199 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6188 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4720 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5443 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5454 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5465 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4731 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4742 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4753 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5476 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5487 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5498 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4764 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4775 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4786 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4797 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8091 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8080 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7390 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9709 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_437 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_426 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_415 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_404 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_3/AMP_IN SF_IB
+ pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_459 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_448 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4005 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4016 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3304 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4027 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4038 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4049 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2603 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3315 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3326 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3337 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3348 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2614 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2625 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2636 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3359 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1902 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1913 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1924 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2647 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2658 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2669 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1935 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1946 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1957 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1968 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1979 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5240 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_982 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_971 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_960 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5251 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5262 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5273 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_993 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4550 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4561 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4572 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5284 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5295 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3860 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4583 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4594 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3871 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3882 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3893 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_90 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_90/AMP_IN SF_IB
+ pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1209 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9528 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9517 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9506 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9539 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8827 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8816 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8805 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8849 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8838 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_201 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_212 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_223 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_234 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_245 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_256 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_267 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_278 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_289 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3101 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3112 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2400 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2411 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3123 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3134 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3145 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3156 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2422 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2433 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2444 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3167 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3178 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3189 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1710 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1721 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1732 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1743 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2455 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2466 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2477 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1754 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1765 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1776 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2488 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2499 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1787 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1798 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_790 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5070 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5081 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4380 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5092 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4391 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3690 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1028 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1017 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1006 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1039 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9303 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9336 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9325 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9314 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9369 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9358 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9347 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8635 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8624 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8613 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8602 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8668 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8657 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8646 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7923 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7912 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7901 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8679 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7956 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7945 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7934 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7989 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7978 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7967 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2230 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2241 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2252 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1540 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1551 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2263 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2274 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2285 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2296 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1562 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1573 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1584 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1595 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9892 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9881 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9870 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7219 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7208 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6507 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6529 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6518 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5806 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5817 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5828 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5839 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9111 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9100 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9144 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9133 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9122 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8410 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9188 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9177 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9166 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9155 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8443 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8432 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8421 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9199 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8476 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8465 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8454 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7731 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7720 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8498 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8487 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7775 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7764 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7753 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7742 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7797 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7786 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2060 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2071 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2082 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2093 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1392 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1381 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1370 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7027 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7016 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7005 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7049 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7038 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6315 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6304 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6359 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6348 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6337 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6326 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5603 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5614 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4902 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5625 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5636 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5647 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4913 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4924 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4935 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4946 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5658 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5669 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4957 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4968 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4979 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8251 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8240 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8284 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8273 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8262 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7550 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8295 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7583 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7572 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7561 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7594 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6871 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6860 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6893 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6882 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_619 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_608 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4209 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3508 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3519 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2807 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2818 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2829 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6101 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6112 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6123 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6134 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6167 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6156 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5400 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5411 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5422 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6145 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6189 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6178 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4710 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4721 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5433 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5444 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5455 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4732 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4743 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4754 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5466 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5477 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5488 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5499 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4765 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4776 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4787 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4798 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8092 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8081 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8070 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7391 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7380 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6690 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_427 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_416 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_405 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_449 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_438 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_4/AMP_IN SF_IB
+ pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4006 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3305 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4017 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4028 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4039 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3316 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3327 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3338 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2604 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2615 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2626 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3349 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1903 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1914 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1925 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2637 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2648 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2659 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1936 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1947 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1958 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1969 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_950 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5230 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_983 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_972 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_961 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5241 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5252 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5263 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5274 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_994 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4540 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4551 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4562 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5285 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5296 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3850 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3861 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4573 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4584 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4595 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3872 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3883 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3894 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_91 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_91/AMP_IN SF_IB
+ pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_80 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_80/AMP_IN SF_IB
+ pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9529 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9518 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9507 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8817 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8806 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8839 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8828 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_202 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_213 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_224 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_235 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_246 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_257 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_268 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_279 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3102 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3113 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2401 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3124 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3135 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3146 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1700 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2412 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2423 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2434 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2445 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3157 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3168 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3179 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1711 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1722 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1733 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2456 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2467 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2478 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1744 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1755 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1766 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2489 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1777 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1788 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1799 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_791 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_780 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5060 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5071 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5082 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4370 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5093 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4381 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4392 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3680 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3691 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2990 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1029 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1018 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1007 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9337 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9326 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9315 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9304 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9359 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9348 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8625 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8614 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8603 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8669 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8658 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8647 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8636 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7924 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7913 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7902 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7957 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7946 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7935 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7979 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7968 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2220 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2231 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2242 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2253 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1530 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1541 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2264 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2275 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2286 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1552 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1563 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1574 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1585 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2297 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1596 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9893 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9882 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9871 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9860 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7209 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6508 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6519 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5807 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5818 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5829 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9112 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9101 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9145 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9134 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9123 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8400 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9178 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9167 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9156 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8433 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8422 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8411 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9189 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8477 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8466 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8455 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8444 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7732 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7721 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7710 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8499 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8488 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7765 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7754 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7743 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7798 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7787 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7776 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2050 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2061 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1360 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2072 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2083 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2094 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1393 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1382 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1371 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9690 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7028 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7017 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7006 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7039 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6316 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6305 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6349 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6338 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6327 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5604 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4903 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5615 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5626 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5637 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5648 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4914 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4925 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4936 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5659 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4947 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4958 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4969 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8252 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8241 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8230 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8285 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8274 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8263 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7540 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8296 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7573 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7562 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7551 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7595 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7584 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6872 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6861 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6850 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6894 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6883 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1190 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_609 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3509 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2808 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2819 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6102 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6113 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6124 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6157 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6146 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5401 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5412 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5423 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6135 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6179 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6168 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4700 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4711 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5434 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5445 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5456 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4722 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4733 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4744 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5467 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5478 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5489 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4755 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4766 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4777 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4788 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4799 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8060 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8093 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8082 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8071 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7392 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7381 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7370 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6680 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6691 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5990 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_428 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_417 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_406 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_439 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_5/AMP_IN SF_IB
+ pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4007 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4018 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4029 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3306 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3317 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3328 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3339 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2605 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2616 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2627 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1904 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1915 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2638 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2649 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1926 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1937 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1948 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1959 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_940 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5220 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5231 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_973 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_962 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_951 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5242 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5253 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5264 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_995 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_984 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4530 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4541 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4552 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4563 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5275 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5286 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5297 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3840 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3851 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4574 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4585 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4596 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3862 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3873 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3884 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3895 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_70 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_70/AMP_IN SF_IB
+ pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_92 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_92/AMP_IN SF_IB
+ pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_81 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_81/AMP_IN SF_IB
+ pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9519 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9508 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8818 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8807 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8829 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_203 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_214 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_225 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_236 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_247 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_258 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_269 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3103 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2402 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3114 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3125 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3136 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3147 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2413 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2424 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2435 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3158 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3169 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1701 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1712 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1723 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1734 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2446 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2457 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2468 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1745 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1756 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1767 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2479 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1778 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1789 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_792 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_781 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_770 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5050 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5061 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5072 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4360 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4371 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5083 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5094 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4382 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4393 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3670 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3681 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3692 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2980 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2991 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1019 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1008 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9327 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9316 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9305 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9349 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9338 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8626 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8615 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8604 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8659 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8648 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8637 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7914 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7903 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7947 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7936 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7925 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7969 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7958 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2210 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2221 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2232 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2243 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1531 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1520 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1542 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2254 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2265 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2276 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2287 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1553 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1564 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1575 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2298 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1586 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1597 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9850 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9883 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9872 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9861 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9894 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4190 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6509 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5808 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5819 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9102 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9135 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9124 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9113 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8401 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9179 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9168 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9157 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9146 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8434 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8423 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8412 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8467 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8456 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8445 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7722 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7711 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7700 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8489 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8478 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7766 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7755 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7744 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7733 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7799 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7788 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7777 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2040 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2051 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2062 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1350 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2073 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2084 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2095 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1383 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1372 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1361 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1394 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9691 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9680 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8990 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7018 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7007 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7029 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6306 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6339 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6328 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6317 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5605 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5616 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5627 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5638 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4904 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4915 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4926 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4937 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5649 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4948 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4959 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8242 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8231 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8220 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8275 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8264 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8253 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7541 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7530 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8297 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8286 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7574 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7563 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7552 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7596 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7585 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6862 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6851 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6840 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6895 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6884 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6873 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1191 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1180 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2809 GRING VDD GND VREF ROW_SEL[28] NB1 VBIAS NB2 pixel_fill_2809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6103 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6114 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6125 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6158 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6147 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5402 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5413 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6136 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6169 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4701 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4712 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5424 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5435 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5446 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4723 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4734 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4745 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5457 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5468 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5479 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4756 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4767 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4778 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4789 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8050 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8094 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8083 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8072 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8061 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7382 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7371 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7360 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7393 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6681 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6670 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6692 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5980 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5991 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_418 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_407 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_429 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_6/AMP_IN SF_IB
+ pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4008 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4019 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3307 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3318 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3329 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2606 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2617 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1905 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1916 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2628 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2639 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1927 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1938 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1949 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_941 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_930 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5210 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5221 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_974 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_963 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_952 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4520 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5232 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5243 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5254 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5265 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_996 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_985 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4531 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4542 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4553 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5276 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5287 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5298 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3830 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3841 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3852 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4564 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4575 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4586 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3863 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3874 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3885 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4597 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3896 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7190 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_60 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_60/AMP_IN SF_IB
+ pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_93 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_93/AMP_IN SF_IB
+ pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_82 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_82/AMP_IN SF_IB
+ pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_71 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_71/AMP_IN SF_IB
+ pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9509 GRING VDD GND VREF ROW_SEL[95] NB1 VBIAS NB2 pixel_fill_9509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8808 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8819 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_204 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_215 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_226 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_237 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_248 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_259 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3104 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3115 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3126 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3137 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2403 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2414 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2425 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2436 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3148 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3159 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1702 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1713 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1724 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2447 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2458 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2469 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1735 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1746 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1757 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1768 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1779 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5040 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_782 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_771 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_760 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5051 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5062 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5073 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_793 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4350 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4361 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5084 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5095 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3660 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4372 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4383 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4394 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3671 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3682 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3693 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2970 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2981 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2992 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1009 GRING VDD GND VREF ROW_SEL[10] NB1 VBIAS NB2 pixel_fill_1009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9328 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9317 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9306 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9339 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8616 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8605 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8649 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8638 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8627 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7915 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7904 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7948 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7937 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7926 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7959 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2200 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2211 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2222 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2233 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2244 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1532 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1521 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1510 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2255 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2266 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2277 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1543 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1554 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1565 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1576 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2288 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2299 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1587 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1598 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9840 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9884 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9873 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9862 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9851 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9895 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_590 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4180 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4191 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3490 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5809 GRING VDD GND VREF ROW_SEL[58] NB1 VBIAS NB2 pixel_fill_5809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9103 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9136 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9125 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9114 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9169 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9158 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9147 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8424 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8413 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8402 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8468 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8457 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8446 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8435 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7723 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7712 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7701 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8479 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7756 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7745 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7734 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7789 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7778 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7767 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2030 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2041 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2052 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1351 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1340 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2063 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2074 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2085 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1384 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1373 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1362 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2096 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1395 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9692 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9681 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9670 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8980 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8991 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7019 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7008 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6307 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6329 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6318 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5606 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5617 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5628 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5639 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4905 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4916 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4927 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4938 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4949 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8243 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8232 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8221 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8210 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8276 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8265 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8254 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7531 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7520 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8298 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8287 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7564 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7553 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7542 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6830 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7597 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7586 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7575 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6863 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6852 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6841 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6896 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6885 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6874 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1192 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1181 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1170 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6104 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6115 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6148 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5403 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5414 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6126 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6137 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6159 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4702 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5425 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5436 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5447 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4713 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4724 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4735 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5458 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5469 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4746 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4757 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4768 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4779 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8051 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8040 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8084 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8073 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8062 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8095 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7383 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7372 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7361 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7350 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7394 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6671 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6660 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6693 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6682 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5970 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5981 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5992 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_419 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_408 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_7/AMP_IN SF_IB
+ pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4009 GRING VDD GND VREF ROW_SEL[40] NB1 VBIAS NB2 pixel_fill_4009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3308 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3319 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2607 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2618 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1906 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2629 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1917 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1928 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1939 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_931 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_920 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5200 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5211 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5222 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_964 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_953 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_942 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4510 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5233 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5244 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5255 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_997 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_986 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_975 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4521 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4532 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4543 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4554 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5266 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5277 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5288 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3820 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3831 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3842 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4565 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4576 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4587 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5299 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3853 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3864 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3875 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4598 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3886 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3897 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7191 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7180 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_61 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_61/AMP_IN SF_IB
+ pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_50 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_50/AMP_IN SF_IB
+ pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6490 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_94 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_94/AMP_IN SF_IB
+ pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_83 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_83/AMP_IN SF_IB
+ pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_72 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_72/AMP_IN SF_IB
+ pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8809 GRING VDD GND VREF ROW_SEL[88] NB1 VBIAS NB2 pixel_fill_8809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_205 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_216 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_227 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_238 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_249 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3105 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3116 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3127 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3138 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2404 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2415 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2426 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3149 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1703 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1714 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1725 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2437 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2448 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2459 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1736 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1747 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1758 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1769 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5030 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_783 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_772 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_761 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_750 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5041 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5052 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5063 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_794 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4340 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4351 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4362 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5074 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5085 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5096 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3650 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4373 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4384 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4395 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3661 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3672 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3683 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3694 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2960 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2971 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2982 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2993 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9318 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9307 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9329 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8617 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8606 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8639 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8628 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7905 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7938 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7927 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7916 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7949 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2201 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1500 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2212 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2223 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2234 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1533 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1522 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1511 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2245 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2256 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2267 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2278 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1544 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1555 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1566 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2289 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1577 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1588 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1599 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9841 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9830 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9874 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9863 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9852 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9896 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9885 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_591 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_580 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4170 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4181 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4192 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3480 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3491 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2790 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9126 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9115 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9104 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9159 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9148 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9137 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8425 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8414 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8403 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8458 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8447 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8436 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7713 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7702 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8469 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7757 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7746 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7735 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7724 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7779 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7768 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2020 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2031 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2042 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2053 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1341 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1330 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2064 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2075 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2086 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1374 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1363 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1352 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2097 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1396 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1385 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9682 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9671 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9660 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9693 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8981 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8970 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8992 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7009 GRING VDD GND VREF ROW_SEL[70] NB1 VBIAS NB2 pixel_fill_7009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6319 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6308 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5607 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5618 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5629 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4906 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4917 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4928 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4939 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8200 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8233 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8222 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8211 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8266 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8255 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8244 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7532 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7521 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7510 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8299 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8288 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8277 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7565 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7554 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7543 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6820 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7598 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7587 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7576 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6853 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6842 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6831 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6897 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6886 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6875 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6864 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1193 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1182 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1171 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1160 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9490 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6105 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6116 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6149 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5404 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6127 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6138 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4703 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5415 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5426 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5437 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4714 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4725 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4736 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5448 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5459 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4747 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4758 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4769 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8041 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8030 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8085 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8074 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8063 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8052 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7340 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8096 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7373 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7362 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7351 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7395 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7384 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6672 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6661 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6650 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6694 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6683 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5960 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5971 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5982 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5993 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_409 GRING VDD GND VREF ROW_SEL[4] NB1 VBIAS NB2 pixel_fill_409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_8/AMP_IN SF_IB
+ pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3309 GRING VDD GND VREF ROW_SEL[33] NB1 VBIAS NB2 pixel_fill_3309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2608 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1907 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2619 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1918 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1929 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_932 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_921 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_910 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5201 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5212 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_965 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_954 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_943 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4500 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4511 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5223 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5234 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5245 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5256 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_998 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_987 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_976 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4522 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4533 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4544 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5267 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5278 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5289 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3810 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3821 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3832 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3843 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4555 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4566 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4577 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3854 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3865 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3876 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4588 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4599 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3887 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3898 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7181 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7170 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7192 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6480 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_51 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_51/AMP_IN SF_IB
+ pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_40 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_40/AMP_IN SF_IB
+ pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6491 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_95 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_95/AMP_IN SF_IB
+ pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_84 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_84/AMP_IN SF_IB
+ pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_73 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_73/AMP_IN SF_IB
+ pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_62 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_62/AMP_IN SF_IB
+ pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5790 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_206 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_217 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_228 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_239 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3106 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3117 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3128 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2405 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2416 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2427 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3139 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1704 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1715 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2438 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2449 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1726 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1737 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1748 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1759 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_740 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5020 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5031 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_773 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_762 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_751 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5042 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5053 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5064 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_795 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_784 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4330 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4341 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4352 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5075 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5086 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5097 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3640 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3651 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4363 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4374 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4385 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4396 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3662 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3673 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3684 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2950 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2961 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2972 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3695 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2983 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2994 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9319 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9308 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8607 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8629 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8618 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7906 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7939 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7928 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7917 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2202 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2213 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2224 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2235 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1523 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1512 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1501 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2246 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2257 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2268 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1534 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1545 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1556 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1567 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2279 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1578 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1589 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9831 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9820 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9875 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9864 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9853 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9842 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9897 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9886 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_581 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_570 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_592 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4160 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4171 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4182 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4193 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3470 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3481 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3492 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2780 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2791 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9127 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9116 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9105 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9149 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9138 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8415 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8404 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8459 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8448 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8437 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8426 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7714 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7703 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7747 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7736 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7725 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7769 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7758 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2010 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2021 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2032 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2043 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1342 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1331 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1320 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2054 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2065 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2076 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1375 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1364 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1353 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2087 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2098 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1397 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1386 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9683 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9672 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9661 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9650 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9694 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8971 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8960 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8993 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8982 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6309 GRING VDD GND VREF ROW_SEL[63] NB1 VBIAS NB2 pixel_fill_6309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5608 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5619 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4907 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4918 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4929 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8234 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8223 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8212 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8201 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8267 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8256 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8245 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7522 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7511 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7500 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8289 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8278 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7555 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7544 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7533 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6821 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6810 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7599 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7588 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7577 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7566 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6854 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6843 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6832 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6887 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6876 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6865 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6898 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1150 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1183 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1172 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1161 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1194 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9491 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9480 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8790 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6106 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5405 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6117 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6128 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6139 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5416 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5427 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5438 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4704 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4715 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4726 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5449 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4737 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4748 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4759 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8042 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8031 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8020 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8075 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8064 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8053 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7330 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8097 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8086 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7374 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7363 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7352 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7341 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7396 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7385 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6662 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6651 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6640 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6695 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6684 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6673 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5950 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5961 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5972 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5983 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5994 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_9/AMP_IN SF_IB
+ pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2609 GRING VDD GND VREF ROW_SEL[26] NB1 VBIAS NB2 pixel_fill_2609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1908 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1919 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_922 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_911 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_900 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5202 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5213 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_955 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_944 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_933 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4501 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5224 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5235 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5246 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_999 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_988 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_977 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_966 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3800 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4512 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4523 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4534 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4545 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5257 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5268 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5279 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3811 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3822 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3833 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4556 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4567 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4578 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3844 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3855 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3866 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4589 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3877 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3888 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3899 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7182 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7171 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7160 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7193 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6470 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_52 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_52/AMP_IN SF_IB
+ pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_41 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_41/AMP_IN SF_IB
+ pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_30 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_30/AMP_IN SF_IB
+ pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6492 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6481 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_85 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_85/AMP_IN SF_IB
+ pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_74 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_74/AMP_IN SF_IB
+ pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_63 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_63/AMP_IN SF_IB
+ pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_96 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_96/AMP_IN SF_IB
+ pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5780 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5791 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_207 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_218 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_229 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3107 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3118 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3129 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2406 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2417 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1705 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1716 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2428 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2439 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1727 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1738 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1749 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_730 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5010 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5021 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_774 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_763 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_752 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_741 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5032 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5043 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5054 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_796 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_785 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4320 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4331 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4342 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4353 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5065 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5076 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5087 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5098 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3630 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3641 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4364 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4375 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4386 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2940 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3652 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3663 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3674 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3685 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4397 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2951 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2962 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2973 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3696 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2984 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2995 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9309 GRING VDD GND VREF ROW_SEL[93] NB1 VBIAS NB2 pixel_fill_9309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8608 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8619 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7929 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7918 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7907 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2203 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2214 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2225 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1524 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1513 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1502 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2236 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2247 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2258 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2269 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1535 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1546 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1557 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1568 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1579 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9832 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9821 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9810 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9865 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9854 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9843 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9898 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9887 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9876 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_582 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_571 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_560 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_593 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4150 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4161 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4172 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4183 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4194 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3460 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3471 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3482 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3493 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2770 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2781 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2792 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9117 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9106 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9139 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9128 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8416 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8405 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8449 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8438 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8427 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7704 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7748 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7737 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7726 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7715 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7759 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2000 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2011 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2022 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2033 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2044 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1332 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1321 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1310 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2055 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2066 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2077 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1365 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1354 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1343 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2088 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2099 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1398 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1387 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1376 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9640 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9673 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9662 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9651 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9695 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9684 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8972 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8961 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8950 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8994 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8983 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_390 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3290 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5609 GRING VDD GND VREF ROW_SEL[56] NB1 VBIAS NB2 pixel_fill_5609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4908 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4919 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8224 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8213 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8202 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8257 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8246 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8235 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7523 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7512 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7501 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8279 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8268 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7556 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7545 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7534 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6811 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6800 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7589 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7578 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7567 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6844 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6833 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6822 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6888 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6877 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6866 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6855 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6899 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1140 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1173 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1162 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1151 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1195 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1184 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9481 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9470 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9492 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8780 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8791 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6107 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6118 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6129 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5406 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5417 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5428 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4705 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4716 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4727 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5439 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4738 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4749 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8032 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8021 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8010 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8076 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8065 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8054 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8043 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7331 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7320 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8098 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8087 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7364 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7353 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7342 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7397 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7386 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7375 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6652 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6641 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6630 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6696 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6685 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6674 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6663 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5940 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5951 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5962 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5973 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5984 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5995 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1909 GRING VDD GND VREF ROW_SEL[19] NB1 VBIAS NB2 pixel_fill_1909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_923 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_912 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_901 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5203 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_956 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_945 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_934 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4502 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5214 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5225 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5236 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5247 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_989 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_978 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_967 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4513 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4524 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4535 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5258 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5269 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3801 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3812 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3823 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3834 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4546 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4557 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4568 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3845 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3856 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3867 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4579 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3878 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3889 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7172 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7161 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7150 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7194 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7183 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6471 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6460 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_42 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_42/AMP_IN SF_IB
+ pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_31 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_31/AMP_IN SF_IB
+ pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_20 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_20/AMP_IN SF_IB
+ pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6493 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6482 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_86 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_86/AMP_IN SF_IB
+ pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_75 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_75/AMP_IN SF_IB
+ pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_64 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_64/AMP_IN SF_IB
+ pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_53 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_53/AMP_IN SF_IB
+ pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_97 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_97/AMP_IN SF_IB
+ pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5770 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5781 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5792 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_208 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_219 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3108 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3119 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2407 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2418 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1706 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2429 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1717 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1728 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1739 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_731 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_720 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5000 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5011 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5022 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_764 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_753 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_742 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4310 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5033 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5044 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5055 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_797 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_786 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_775 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4321 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4332 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4343 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5066 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5077 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5088 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3620 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3631 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3642 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4354 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4365 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4376 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4387 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5099 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2930 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3653 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3664 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3675 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4398 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2941 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2952 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2963 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3686 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3697 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2974 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2985 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2996 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6290 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8609 GRING VDD GND VREF ROW_SEL[86] NB1 VBIAS NB2 pixel_fill_8609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7919 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7908 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2204 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2215 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2226 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1514 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1503 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2237 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2248 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2259 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1536 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1525 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1547 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1558 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1569 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9822 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9811 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9800 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9866 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9855 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9844 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9833 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9899 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9888 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9877 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_572 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_561 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_550 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_594 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_583 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4140 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4151 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3450 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4162 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4173 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4184 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4195 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3461 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3472 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3483 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2760 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2771 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2782 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3494 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2793 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9118 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9107 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9129 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8406 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8439 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8428 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8417 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7705 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7738 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7727 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7716 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7749 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2001 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2012 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2023 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2034 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1322 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1311 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1300 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2045 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2056 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2067 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1366 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1355 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1344 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1333 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2078 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2089 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1399 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1388 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1377 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9630 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9674 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9663 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9652 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9641 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9696 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9685 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8962 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8951 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8940 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8995 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8984 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8973 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_380 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_391 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3280 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3291 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2590 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4909 GRING VDD GND VREF ROW_SEL[49] NB1 VBIAS NB2 pixel_fill_4909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8225 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8214 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8203 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8258 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8247 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8236 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7513 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7502 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8269 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7546 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7535 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7524 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6801 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7579 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7568 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7557 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6845 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6834 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6823 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6812 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6878 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6867 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6856 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6889 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1141 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1130 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1174 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1163 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1152 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1196 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1185 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9482 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9471 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9460 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9493 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8770 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8792 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8781 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6108 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6119 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5407 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5418 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5429 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4706 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4717 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4728 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4739 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8000 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8033 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8022 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8011 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8066 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8055 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8044 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7321 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7310 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8099 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8088 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8077 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7365 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7354 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7343 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7332 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6620 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7398 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7387 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7376 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6653 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6642 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6631 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6686 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6675 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6664 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5930 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5941 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6697 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5952 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5963 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5974 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5985 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5996 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9290 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_913 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_902 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5204 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_946 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_935 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_924 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5215 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5226 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5237 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_979 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_968 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_957 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4503 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4514 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4525 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4536 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5248 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5259 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3802 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3813 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3824 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4547 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4558 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4569 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3835 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3846 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3857 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3868 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3879 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7173 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7162 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7151 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7140 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7195 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7184 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6461 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6450 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_43 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_43/AMP_IN SF_IB
+ pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_32 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_32/AMP_IN SF_IB
+ pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_21 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_21/AMP_IN SF_IB
+ pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_10 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_10/AMP_IN SF_IB
+ pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6494 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6483 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6472 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_76 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_76/AMP_IN SF_IB
+ pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_65 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_65/AMP_IN SF_IB
+ pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_54 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_54/AMP_IN SF_IB
+ pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5760 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_87 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_87/AMP_IN SF_IB
+ pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_98 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_98/AMP_IN SF_IB
+ pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5771 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5782 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5793 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_209 GRING VDD GND VREF ROW_SEL[2] NB1 VBIAS NB2 pixel_fill_209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3109 GRING VDD GND VREF ROW_SEL[31] NB1 VBIAS NB2 pixel_fill_3109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2408 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1707 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2419 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1718 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1729 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_721 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_710 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5001 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5012 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_765 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_754 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_743 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_732 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4300 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5023 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5034 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5045 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_798 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_787 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_776 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4311 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4322 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4333 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4344 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5056 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5067 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5078 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5089 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3610 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3621 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3632 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4355 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4366 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4377 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2920 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2931 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3643 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3654 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3665 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3676 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4388 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4399 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2942 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2953 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2964 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3687 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3698 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2975 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2986 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2997 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6291 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6280 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5590 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7909 GRING VDD GND VREF ROW_SEL[79] NB1 VBIAS NB2 pixel_fill_7909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2205 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2216 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1515 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1504 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2227 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2238 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2249 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1537 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1526 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1548 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1559 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9823 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9812 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9801 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9856 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9845 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9834 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9889 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9878 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9867 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_573 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_562 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_551 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_540 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_595 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_584 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4130 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4141 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4152 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3440 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4163 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4174 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4185 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3451 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3462 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3473 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3484 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4196 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2750 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2761 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2772 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3495 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2783 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2794 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9108 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9119 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8407 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8429 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8418 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7739 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7728 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7717 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7706 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2002 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2013 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2024 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2035 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1323 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1312 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1301 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2046 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2057 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2068 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1356 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1345 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1334 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2079 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1389 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1378 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1367 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9631 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9620 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9664 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9653 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9642 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9697 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9686 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9675 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8963 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8952 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8941 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8930 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8996 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8985 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8974 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_370 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_381 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_392 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3270 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3281 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3292 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2580 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2591 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1890 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8215 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8204 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8248 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8237 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8226 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7514 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7503 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8259 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7547 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7536 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7525 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6802 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7569 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7558 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6835 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6824 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6813 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6879 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6868 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6857 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6846 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1131 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1120 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1164 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1153 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1142 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1197 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1186 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1175 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9472 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9461 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9450 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9494 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9483 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8771 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8760 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8793 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8782 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6109 GRING VDD GND VREF ROW_SEL[61] NB1 VBIAS NB2 pixel_fill_6109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5408 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5419 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4707 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4718 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4729 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8023 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8012 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8001 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8067 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8056 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8045 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8034 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7322 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7311 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7300 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8089 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8078 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7355 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7344 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7333 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6610 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7388 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7377 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7366 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6643 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6632 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6621 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7399 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6687 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6676 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6665 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6654 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5920 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5931 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5942 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6698 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5953 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5964 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5975 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5986 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5997 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9291 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9280 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8590 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_914 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_903 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_947 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_936 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_925 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5205 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5216 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5227 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5238 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_969 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_958 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4504 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4515 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4526 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5249 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3803 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3814 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3825 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4537 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4548 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4559 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3836 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3847 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3858 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3869 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7130 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7163 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7152 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7141 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7196 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7185 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7174 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6462 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6451 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6440 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_33 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_33/AMP_IN SF_IB
+ pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_22 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_22/AMP_IN SF_IB
+ pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_11 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_11/AMP_IN SF_IB
+ pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6495 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6484 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6473 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_77 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_77/AMP_IN SF_IB
+ pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_66 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_66/AMP_IN SF_IB
+ pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_55 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_55/AMP_IN SF_IB
+ pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_44 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_44/AMP_IN SF_IB
+ pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5750 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_88 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_88/AMP_IN SF_IB
+ pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_99 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_99/AMP_IN SF_IB
+ pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5761 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5772 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5783 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5794 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2409 GRING VDD GND VREF ROW_SEL[24] NB1 VBIAS NB2 pixel_fill_2409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1708 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1719 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_722 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_711 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_700 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5002 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5013 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_755 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_744 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_733 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4301 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5024 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5035 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5046 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_788 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_777 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_766 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4312 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4323 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4334 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5057 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5068 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5079 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_799 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3600 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3611 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3622 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3633 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4345 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4356 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4367 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4378 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2910 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2921 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3644 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3655 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3666 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4389 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2932 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2943 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2954 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3677 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3688 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3699 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2965 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2976 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2987 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2998 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6270 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6292 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6281 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5580 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5591 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4890 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2206 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2217 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1505 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2228 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2239 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1527 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1516 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1538 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1549 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9813 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9802 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9857 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9846 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9835 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9824 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9879 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9868 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_530 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_563 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_552 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_541 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_596 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_585 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_574 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4120 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4131 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4142 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3430 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3441 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4153 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4164 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4175 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4186 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3452 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3463 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3474 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4197 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2740 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2751 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2762 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2773 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3485 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3496 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2784 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2795 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9109 GRING VDD GND VREF ROW_SEL[91] NB1 VBIAS NB2 pixel_fill_9109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8419 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8408 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7729 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7718 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7707 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2003 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2014 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2025 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1313 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1302 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2036 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2047 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2058 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1357 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1346 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1335 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1324 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2069 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1379 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1368 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9621 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9610 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9665 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9654 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9643 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9632 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8920 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9698 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9687 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9676 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8953 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8942 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8931 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8997 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8986 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8975 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8964 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_360 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_371 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_393 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_382 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3260 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3271 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3282 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2570 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2581 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3293 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2592 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1880 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1891 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8216 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8216/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8205 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8205/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8249 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8249/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8238 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8238/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8227 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8227/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7504 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7537 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7526 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7515 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7559 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7548 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6836 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6825 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6814 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6803 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6869 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6858 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6847 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1132 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1121 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1110 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1165 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1154 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1143 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1198 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1187 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1176 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9440 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9473 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9462 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9451 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9495 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9484 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8761 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8761/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8750 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8750/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8794 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8794/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8783 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8783/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8772 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8772/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_190 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3090 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5409 GRING VDD GND VREF ROW_SEL[54] NB1 VBIAS NB2 pixel_fill_5409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4708 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4719 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8024 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8024/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8013 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8013/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8002 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8002/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8057 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8057/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8046 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8046/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8035 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8035/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7312 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7301 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8079 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8079/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8068 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8068/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7356 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7345 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7334 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7323 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6611 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6600 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7389 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7378 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7367 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6644 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6633 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6622 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6677 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6666 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6655 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5910 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5921 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5932 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6699 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6688 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5943 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5954 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5965 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5976 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5987 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5998 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9281 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9270 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9292 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8580 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8580/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8591 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8591/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7890 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_904 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_937 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_926 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_915 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5206 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5217 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5228 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_959 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_948 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4505 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4516 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4527 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5239 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3804 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3815 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4538 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4549 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3826 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3837 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3848 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3859 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7120 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7164 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7153 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7142 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7131 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7197 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7186 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7175 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6452 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6441 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6430 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_34 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_34/AMP_IN SF_IB
+ pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_23 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_23/AMP_IN SF_IB
+ pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_12 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_12/AMP_IN SF_IB
+ pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6485 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6474 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6463 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_67 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_67/AMP_IN SF_IB
+ pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_56 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_56/AMP_IN SF_IB
+ pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_45 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_45/AMP_IN SF_IB
+ pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5740 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5751 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6496 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_89 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_89/AMP_IN SF_IB
+ pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_78 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_78/AMP_IN SF_IB
+ pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5762 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5773 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5784 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5795 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1709 GRING VDD GND VREF ROW_SEL[17] NB1 VBIAS NB2 pixel_fill_1709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_712 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_701 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5003 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_756 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_745 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_734 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_723 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5014 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5025 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5036 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_789 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_778 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_767 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4302 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4313 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4324 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4335 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5047 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5058 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5069 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3601 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3612 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3623 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4346 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4357 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4368 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2900 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2911 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2922 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3634 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3645 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3656 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3667 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4379 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2933 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2944 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2955 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3678 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3689 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2966 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2977 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2988 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2999 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6260 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6293 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6282 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6271 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5570 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5581 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5592 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4880 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4891 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2207 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1506 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2218 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2229 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1528 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1517 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1539 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9814 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9814/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9803 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9803/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9847 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9847/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9836 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9836/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9825 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9825/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9869 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9869/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9858 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9858/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_520 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_564 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_553 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_542 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_531 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4110 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_597 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_586 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_575 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4121 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4132 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4143 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3420 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3431 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4154 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4165 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4176 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2730 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3442 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3453 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3464 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3475 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4187 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4198 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2741 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2752 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2763 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3486 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3497 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2774 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2785 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2796 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6090 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8409 GRING VDD GND VREF ROW_SEL[84] NB1 VBIAS NB2 pixel_fill_8409/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7719 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7708 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2004 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2015 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2026 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1314 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1303 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2037 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2048 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2059 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1347 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1336 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1325 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1369 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1358 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9622 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9622/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9611 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9611/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9600 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9600/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9655 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9655/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9644 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9644/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9633 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9633/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8910 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8910/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9699 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9699/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9688 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9688/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9677 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9677/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9666 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9666/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8954 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8954/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8943 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8943/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8932 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8932/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8921 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8921/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8987 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8987/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8976 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8976/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8965 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8965/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8998 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8998/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_350 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_361 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_372 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_394 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_383 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3250 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3261 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3272 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3283 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2560 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2571 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3294 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1870 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2582 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2593 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1881 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1892 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8206 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8206/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8239 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8239/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8228 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8228/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8217 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8217/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7505 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7538 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7527 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7516 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7549 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6826 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6815 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6804 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6859 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6848 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6837 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1122 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1111 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1100 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1155 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1144 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1133 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1199 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1188 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1177 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1166 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9430 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9430/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9463 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9463/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9452 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9452/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9441 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9441/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9496 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9496/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9485 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9485/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9474 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9474/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8762 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8762/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8751 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8751/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8740 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8740/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8795 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8795/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8784 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8784/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8773 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8773/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_180 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_191 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3080 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3091 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2390 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4709 GRING VDD GND VREF ROW_SEL[47] NB1 VBIAS NB2 pixel_fill_4709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8014 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8014/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8003 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8003/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8058 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8058/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8047 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8047/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8036 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8036/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8025 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8025/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7313 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7302 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8069 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8069/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7346 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7335 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7324 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6601 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7379 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7368 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7357 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6634 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6623 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6612 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5900 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6678 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6667 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6656 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6645 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5911 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5922 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5933 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6689 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5944 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5955 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5966 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5977 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5988 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5999 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9282 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9282/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9271 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9271/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9260 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9260/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9293 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9293/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8570 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8570/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8592 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8592/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8581 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8581/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7891 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7880 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_905 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_938 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_927 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_916 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5207 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5218 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5229 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_949 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4506 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4517 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3805 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4528 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4539 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3816 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3827 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3838 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3849 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7121 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7110 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7154 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7143 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7132 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7198 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7187 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7176 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7165 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6453 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6442 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6431 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6420 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_24 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_24/AMP_IN SF_IB
+ pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_13 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_13/AMP_IN SF_IB
+ pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6486 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6475 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6464 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_68 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_68/AMP_IN SF_IB
+ pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_57 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_57/AMP_IN SF_IB
+ pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_46 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_46/AMP_IN SF_IB
+ pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_35 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_35/AMP_IN SF_IB
+ pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5730 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5741 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6497 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_79 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_79/AMP_IN SF_IB
+ pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5752 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5763 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5774 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5785 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5796 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9090 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9090/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_713 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_702 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5004 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_746 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_735 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_724 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5015 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5026 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5037 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_779 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_768 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_757 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4303 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4314 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4325 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5048 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5059 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3602 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3613 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3624 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4336 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4347 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4358 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4369 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2901 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2912 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3635 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3646 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3657 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2923 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2934 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2945 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3668 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3679 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2956 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2967 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2978 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2989 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6261 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6250 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6294 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6283 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6272 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5560 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5571 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5582 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5593 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4870 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4881 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4892 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2208 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2219 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1529 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1518 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1507 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9804 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9804/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9848 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9848/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9837 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9837/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9826 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9826/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9815 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9815/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9859 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9859/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_521 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_510 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_554 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_543 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_532 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4100 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_598 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_587 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_576 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_565 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4111 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4122 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4133 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3410 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3421 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3432 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4144 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4155 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4166 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4177 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2720 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3443 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3454 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3465 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4188 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4199 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2731 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2742 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2753 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2764 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3476 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3487 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3498 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2775 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2786 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2797 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6080 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6091 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5390 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7709 GRING VDD GND VREF ROW_SEL[77] NB1 VBIAS NB2 pixel_fill_7709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2005 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2016 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1304 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2027 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2038 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2049 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1348 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1337 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1326 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1315 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1359 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9612 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9612/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9601 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9601/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9656 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9656/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9645 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9645/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9634 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9634/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9623 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9623/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8911 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8911/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8900 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8900/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9689 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9689/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9678 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9678/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9667 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9667/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8944 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8944/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8933 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8933/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8922 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8922/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8977 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8977/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8966 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8966/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8955 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8955/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8999 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8999/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8988 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8988/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_340 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_351 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_362 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_395 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_373 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_384 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3240 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3251 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3262 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3273 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2550 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2561 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2572 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3284 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3295 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1860 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2583 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2594 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1871 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1882 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1893 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8207 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8207/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8229 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8229/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8218 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8218/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7528 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7517 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7506 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7539 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6827 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6816 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6805 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6849 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6838 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1123 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1112 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1101 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1156 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1145 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1134 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1189 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1178 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1167 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9431 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9431/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9420 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9420/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9464 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9464/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9453 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9453/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9442 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9442/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9497 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9497/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9486 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9486/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9475 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9475/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8752 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8752/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8741 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8741/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8730 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8730/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8796 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8796/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8785 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8785/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8774 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8774/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8763 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8763/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_170 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_181 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_192 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3070 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3081 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3092 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2380 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2391 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1690 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8015 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8015/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8004 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8004/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8048 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8048/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8037 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8037/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8026 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8026/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7303 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8059 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8059/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7347 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7336 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7325 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7314 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6602 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7369 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7358 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6635 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6624 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6613 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6668 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6657 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6646 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5901 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5912 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5923 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6679 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5934 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5945 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5956 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5967 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5978 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5989 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9272 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9272/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9261 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9261/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9250 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9250/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9294 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9294/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9283 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9283/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8571 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8571/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8560 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8560/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8593 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8593/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8582 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8582/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7892 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7881 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7870 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_928 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_917 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_906 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5208 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5219 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_939 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4507 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4518 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3806 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4529 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3817 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3828 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3839 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7111 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7100 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7155 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7144 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7133 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7122 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6410 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7188 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7177 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7166 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6443 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6432 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6421 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_25 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_25/AMP_IN SF_IB
+ pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_14 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_14/AMP_IN SF_IB
+ pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7199 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6476 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6465 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6454 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_58 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_58/AMP_IN SF_IB
+ pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_47 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_47/AMP_IN SF_IB
+ pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_36 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_36/AMP_IN SF_IB
+ pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5720 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5731 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5742 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6498 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6487 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_69 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_69/AMP_IN SF_IB
+ pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5753 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5764 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5775 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5786 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5797 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9080 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9080/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9091 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9091/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8390 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8390/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_703 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_747 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_736 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_725 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_714 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5005 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5016 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5027 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_769 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_758 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4304 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4315 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4326 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5038 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5049 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3603 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3614 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4337 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4348 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4359 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2902 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2913 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3625 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3636 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3647 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2924 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2935 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2946 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3658 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3669 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2957 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2968 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2979 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6251 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6240 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6295 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6284 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6273 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6262 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5550 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5561 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5572 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5583 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4860 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4871 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4882 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5594 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4893 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2209 GRING VDD GND VREF ROW_SEL[22] NB1 VBIAS NB2 pixel_fill_2209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1519 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1508 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9805 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9805/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9838 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9838/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9827 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9827/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9816 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9816/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9849 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9849/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_511 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_500 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_555 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_544 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_533 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_522 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4101 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_588 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_577 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_566 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4112 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4123 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4134 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_599 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3400 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3411 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3422 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4145 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4156 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4167 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2710 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2721 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3433 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3444 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3455 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3466 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4178 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4189 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2732 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2743 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2754 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3477 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3488 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3499 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2765 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2776 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2787 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2798 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6070 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6081 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6092 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5380 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5391 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4690 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2006 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2017 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1305 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2028 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2039 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1338 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1327 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1316 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1349 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9613 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9613/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9602 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9602/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9646 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9646/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9635 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9635/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9624 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9624/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8901 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8901/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9679 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9679/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9668 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9668/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9657 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9657/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8945 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8945/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8934 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8934/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8923 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8923/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8912 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8912/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8978 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8978/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8967 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8967/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8956 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8956/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8989 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8989/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_330 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_341 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_352 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_363 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_396 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_374 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_385 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3230 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3241 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3252 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3263 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3274 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2540 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2551 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2562 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3285 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3296 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1850 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1861 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2573 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2584 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2595 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1872 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1883 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1894 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8219 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8219/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8208 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8208/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7529 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7518 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7507 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6817 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6806 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6839 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6828 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1113 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1102 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1146 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1135 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1124 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1179 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1168 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1157 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9421 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9421/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9410 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9410/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9454 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9454/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9443 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9443/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9432 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9432/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8720 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8720/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9498 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9498/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9487 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9487/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9476 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9476/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9465 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9465/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8753 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8753/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8742 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8742/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8731 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8731/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8786 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8786/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8775 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8775/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8764 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8764/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8797 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8797/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_160 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_171 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_182 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_193 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3060 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3071 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3082 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2370 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2381 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3093 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2392 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1680 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1691 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8005 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8005/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8049 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8049/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8038 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8038/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8027 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8027/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8016 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8016/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7304 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7337 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7326 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7315 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7359 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7348 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6625 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6614 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6603 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6669 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6658 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6647 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6636 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5902 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5913 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5924 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5935 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5946 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5957 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5968 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5979 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9273 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9273/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9262 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9262/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9251 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9251/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9240 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9240/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9295 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9295/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9284 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9284/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8561 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8561/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8550 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8550/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8594 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8594/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8583 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8583/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8572 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8572/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7860 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7893 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7882 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7871 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_929 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_918 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_907 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5209 GRING VDD GND VREF ROW_SEL[52] NB1 VBIAS NB2 pixel_fill_5209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4508 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4519 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3807 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3818 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3829 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7112 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7101 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7145 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7134 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7123 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6400 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7189 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7178 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7167 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7156 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6444 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6433 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6422 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6411 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_15 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_15/AMP_IN SF_IB
+ pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6477 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6466 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6455 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_59 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_59/AMP_IN SF_IB
+ pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_48 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_48/AMP_IN SF_IB
+ pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_37 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_37/AMP_IN SF_IB
+ pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_26 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_26/AMP_IN SF_IB
+ pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5710 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5721 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5732 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6499 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6488 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5743 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5754 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5765 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5776 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5787 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5798 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9081 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9081/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9070 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9070/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9092 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9092/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8391 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8391/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8380 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8380/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7690 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_704 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_737 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_726 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_715 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5006 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5017 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5028 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_759 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_748 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4305 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4316 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5039 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3604 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3615 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4327 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4338 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4349 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2903 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3626 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3637 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3648 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2914 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2925 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2936 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3659 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2947 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2958 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2969 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6252 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6241 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6230 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6285 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6274 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6263 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5540 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6296 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5551 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5562 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5573 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5584 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4850 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4861 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4872 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5595 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4883 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4894 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1509 GRING VDD GND VREF ROW_SEL[15] NB1 VBIAS NB2 pixel_fill_1509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9839 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9839/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9828 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9828/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9817 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9817/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9806 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9806/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_512 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_501 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_545 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_534 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_523 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_589 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_578 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_567 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_556 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4102 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4113 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4124 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3401 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3412 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3423 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4135 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4146 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4157 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4168 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2700 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2711 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3434 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3445 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3456 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4179 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2722 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2733 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2744 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2755 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3467 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3478 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3489 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2766 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2777 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2788 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2799 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6060 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6071 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6082 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6093 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5370 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5381 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5392 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4680 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4691 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3990 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2007 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2018 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2029 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1339 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1328 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1317 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1306 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9603 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9603/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9647 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9647/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9636 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9636/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9625 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9625/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9614 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9614/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8902 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8902/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9669 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9669/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9658 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9658/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8935 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8935/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8924 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8924/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8913 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8913/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8968 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8968/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8957 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8957/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8946 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8946/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8979 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8979/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_320 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_331 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_342 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_353 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_397 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_386 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_364 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_375 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3220 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3231 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2530 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3242 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3253 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3264 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2541 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2552 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2563 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3275 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3286 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3297 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1840 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1851 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2574 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2585 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2596 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1862 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1873 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1884 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1895 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8209 GRING VDD GND VREF ROW_SEL[82] NB1 VBIAS NB2 pixel_fill_8209/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7519 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7508 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6818 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6807 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6829 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1114 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1103 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1147 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1136 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1125 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1169 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1158 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9422 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9422/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9411 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9411/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9400 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9400/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9455 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9455/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9444 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9444/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9433 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9433/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8710 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8710/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9488 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9488/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9477 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9477/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9466 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9466/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8743 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8743/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8732 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8732/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8721 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8721/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9499 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9499/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8787 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8787/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8776 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8776/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8765 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8765/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8754 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8754/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8798 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8798/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_150 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_161 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_172 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_183 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_194 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3050 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3061 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3072 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3083 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2360 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2371 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3094 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2382 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2393 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1670 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1681 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1692 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8006 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8006/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8039 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8039/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8028 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8028/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8017 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8017/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7338 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7338/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7327 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7327/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7316 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7316/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7305 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7305/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7349 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7349/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6626 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6615 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6604 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6659 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6648 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6637 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5903 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5914 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5925 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5936 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5947 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5958 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5969 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9230 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9230/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9263 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9263/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9252 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9252/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9241 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9241/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9296 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9296/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9285 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9285/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9274 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9274/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8562 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8562/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8551 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8551/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8540 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8540/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8595 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8595/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8584 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8584/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8573 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8573/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7850 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7850/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7883 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7883/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7872 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7872/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7861 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7861/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7894 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7894/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2190 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_919 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_908 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4509 GRING VDD GND VREF ROW_SEL[45] NB1 VBIAS NB2 pixel_fill_4509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3808 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3819 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7102 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7102/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7146 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7146/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7135 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7135/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7124 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7124/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7113 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7113/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6401 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7179 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7179/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7168 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7168/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7157 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7157/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6434 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6423 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6412 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_16 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_16/AMP_IN SF_IB
+ pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6467 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6456 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6445 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_49 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_49/AMP_IN SF_IB
+ pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_38 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_38/AMP_IN SF_IB
+ pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_27 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_27/AMP_IN SF_IB
+ pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5700 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5711 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5722 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5733 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6489 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6478 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5744 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5755 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5766 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5777 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5788 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5799 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9071 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9071/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9060 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9060/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9093 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9093/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9082 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9082/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8370 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8370/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8392 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8392/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8381 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8381/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7691 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7691/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7680 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7680/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6990 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_738 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_727 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_716 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_705 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5007 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5018 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_749 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4306 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4317 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5029 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3605 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4328 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4339 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2904 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3616 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3627 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3638 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2915 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2926 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2937 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3649 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2948 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2959 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6242 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6231 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6220 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6286 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6275 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6264 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6253 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5530 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5541 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6297 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5552 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5563 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5574 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4840 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4851 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4862 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4873 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5585 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5596 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4884 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4895 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9829 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9829/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9818 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9818/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9807 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9807/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_502 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_546 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_535 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_524 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_513 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_579 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_568 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_557 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4103 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4114 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4125 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3402 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3413 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4136 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4147 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4158 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2701 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2712 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3424 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3435 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3446 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3457 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4169 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2723 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2734 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2745 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3468 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3479 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2756 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2767 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2778 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2789 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6050 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6061 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6072 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6083 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6094 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5360 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5371 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5382 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4670 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4681 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5393 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4692 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3980 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3991 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2008 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2019 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1329 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1318 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1307 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9604 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9604/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9637 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9637/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9626 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9626/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9615 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9615/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9659 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9659/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9648 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9648/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8936 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8936/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8925 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8925/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8914 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8914/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8903 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8903/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8969 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8969/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8958 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8958/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8947 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8947/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_310 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_321 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_332 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_343 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_354 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_387 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_365 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_376 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_398 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3210 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3221 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3232 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2520 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3243 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3254 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3265 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2531 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2542 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2553 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3276 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3287 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3298 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1830 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1841 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1852 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2564 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2575 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2586 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2597 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1863 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1874 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1885 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1896 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5190 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7509 GRING VDD GND VREF ROW_SEL[75] NB1 VBIAS NB2 pixel_fill_7509/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6808 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6819 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1104 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1137 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1126 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1115 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1159 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1148 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9412 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9412/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9401 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9401/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9445 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9445/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9434 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9434/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9423 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9423/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8711 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8711/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8700 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8700/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9489 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9489/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9478 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9478/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9467 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9467/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9456 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9456/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8744 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8744/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8733 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8733/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8722 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8722/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8777 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8777/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8766 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8766/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8755 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8755/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8799 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8799/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8788 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8788/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_140 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_151 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_162 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_173 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_184 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_195 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3040 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3051 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3062 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3073 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2350 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2361 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2372 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3084 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3095 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1660 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2383 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2394 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1671 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1682 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1693 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9990 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9990/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8029 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8029/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8018 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8018/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8007 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8007/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7328 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7328/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7317 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7317/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7306 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7306/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7339 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7339/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6616 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6605 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6649 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6638 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6627 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5904 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5915 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5926 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5937 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5948 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5959 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9220 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9220/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9264 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9264/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9253 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9253/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9242 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9242/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9231 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9231/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9297 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9297/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9286 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9286/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9275 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9275/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8552 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8552/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8541 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8541/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8530 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8530/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8585 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8585/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8574 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8574/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8563 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8563/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7851 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7851/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7840 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7840/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8596 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8596/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7884 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7884/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7873 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7873/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7862 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7862/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7895 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7895/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2180 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2191 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1490 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_909 GRING VDD GND VREF ROW_SEL[9] NB1 VBIAS NB2 pixel_fill_909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3809 GRING VDD GND VREF ROW_SEL[38] NB1 VBIAS NB2 pixel_fill_3809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7103 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7103/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7136 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7136/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7125 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7125/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7114 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7114/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7169 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7169/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7158 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7158/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7147 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7147/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6435 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6424 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6413 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6402 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6468 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6457 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6446 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_39 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_39/AMP_IN SF_IB
+ pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_28 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_28/AMP_IN SF_IB
+ pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_17 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_17/AMP_IN SF_IB
+ pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5701 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5712 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5723 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6479 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5734 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5745 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5756 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5767 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5778 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5789 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9072 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9072/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9061 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9061/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9050 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9050/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9094 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9094/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9083 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9083/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8360 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8360/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8393 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8393/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8382 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8382/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8371 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8371/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7692 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7692/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7681 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7681/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7670 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7670/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6980 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6991 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_728 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_717 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_706 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5008 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5019 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_739 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4307 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3606 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4318 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4329 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3617 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3628 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3639 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2905 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2916 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2927 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2938 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2949 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6210 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6243 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6232 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6221 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6276 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6265 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6254 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5520 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5531 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6298 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6287 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4830 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5542 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5553 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5564 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5575 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4841 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4852 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4863 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5586 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5597 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4874 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4885 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4896 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8190 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8190/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9819 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9819/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9808 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9808/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_503 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_536 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_525 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_514 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_569 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_558 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_547 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4104 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4115 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3403 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3414 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4126 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4137 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4148 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4159 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2702 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3425 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3436 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3447 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2713 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2724 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2735 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2746 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3458 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3469 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2757 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2768 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2779 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6040 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6051 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5350 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6062 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6073 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6084 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5361 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5372 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5383 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6095 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4660 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4671 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5394 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3970 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4682 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4693 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3981 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3992 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2009 GRING VDD GND VREF ROW_SEL[20] NB1 VBIAS NB2 pixel_fill_2009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1319 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1308 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9638 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9638/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9627 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9627/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9616 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9616/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9605 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9605/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9649 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9649/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8926 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8926/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8915 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8915/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8904 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8904/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8959 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8959/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8948 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8948/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8937 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8937/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_300 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_311 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_322 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_333 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_344 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_388 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_355 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_366 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_377 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_399 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3200 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3211 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3222 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2510 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2521 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3233 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3244 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3255 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2532 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2543 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2554 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3266 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3277 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3288 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3299 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1820 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1831 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1842 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2565 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2576 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2587 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1853 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1864 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1875 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1886 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2598 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1897 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5180 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5191 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4490 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6809 GRING VDD GND VREF ROW_SEL[68] NB1 VBIAS NB2 pixel_fill_6809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1105 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1138 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1127 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1116 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1149 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9413 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9413/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9402 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9402/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9446 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9446/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9435 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9435/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9424 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9424/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8701 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8701/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9479 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9479/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9468 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9468/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9457 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9457/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8734 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8734/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8723 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8723/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8712 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8712/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8778 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8778/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8767 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8767/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8756 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8756/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8745 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8745/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8789 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8789/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_130 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_141 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_152 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_163 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_174 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_185 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_196 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3030 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3041 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3052 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3063 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3074 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2340 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2351 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2362 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3085 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3096 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1650 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2373 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2384 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2395 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1661 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1672 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1683 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1694 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9991 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9991/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9980 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9980/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8019 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8019/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8008 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8008/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7329 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7329/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7318 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7318/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7307 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7307/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6617 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6606 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6639 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6628 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5905 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5916 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5927 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5938 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5949 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9221 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9221/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9210 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9210/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9254 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9254/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9243 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9243/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9232 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9232/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9287 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9287/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9276 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9276/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9265 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9265/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8553 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8553/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8542 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8542/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8531 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8531/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8520 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8520/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9298 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9298/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8586 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8586/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8575 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8575/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8564 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8564/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7841 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7841/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7830 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7830/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8597 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8597/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7874 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7874/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7863 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7863/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7852 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7852/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7896 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7896/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7885 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7885/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2170 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2181 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2192 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1491 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1480 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7137 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7137/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7126 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7126/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7115 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7115/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7104 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7104/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7159 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7159/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7148 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7148/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6425 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6414 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6403 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6458 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6447 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6436 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_29 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_29/AMP_IN SF_IB
+ pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_18 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_18/AMP_IN SF_IB
+ pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5702 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5713 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5724 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6469 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5735 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5746 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5757 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5768 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5779 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9062 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9062/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9051 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9051/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9040 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9040/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9095 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9095/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9084 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9084/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9073 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9073/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8361 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8361/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8350 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8350/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8394 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8394/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8383 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8383/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8372 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8372/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7693 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7693/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7682 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7682/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7671 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7671/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7660 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7660/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6981 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6970 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6992 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_729 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_718 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_707 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5009 GRING VDD GND VREF ROW_SEL[50] NB1 VBIAS NB2 pixel_fill_5009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4308 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4319 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3607 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3618 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3629 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2906 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2917 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2928 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2939 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6200 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6233 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6222 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6211 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6277 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6266 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6255 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6244 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5510 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5521 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5532 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6299 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6288 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4820 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5543 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5554 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5565 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4831 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4842 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4853 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4864 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5576 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5587 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5598 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4875 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4886 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4897 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8191 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8191/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8180 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8180/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7490 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7490/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9809 GRING VDD GND VREF ROW_SEL[98] NB1 VBIAS NB2 pixel_fill_9809/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_537 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_537/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_526 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_526/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_515 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_515/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_504 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_504/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_559 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_559/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_548 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_548/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4105 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4116 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3404 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4127 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4138 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4149 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2703 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3415 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3426 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3437 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3448 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2714 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2725 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2736 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3459 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2747 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2758 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2769 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6030 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6041 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6052 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5340 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6063 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6074 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6085 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5351 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5362 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5373 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6096 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4650 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4661 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4672 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5384 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5395 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3960 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4683 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4694 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3971 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3982 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3993 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1309 GRING VDD GND VREF ROW_SEL[13] NB1 VBIAS NB2 pixel_fill_1309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9628 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9628/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9617 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9617/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9606 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9606/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9639 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9639/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8927 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8927/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8916 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8916/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8905 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8905/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8949 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8949/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8938 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8938/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_301 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_301/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_312 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_312/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_323 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_323/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_334 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_334/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_345 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_345/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_356 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_356/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_367 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_367/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_378 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_378/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_389 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_389/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3201 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3212 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3223 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2500 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2511 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3234 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3245 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3256 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2522 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2533 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2544 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3267 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3278 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3289 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1810 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1821 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1832 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1843 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2555 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2566 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2577 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2588 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1854 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1865 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1876 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2599 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1887 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1898 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_890 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_890/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5170 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5181 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5192 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4480 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4491 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3790 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1128 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1117 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1106 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1139 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9403 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9403/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9436 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9436/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9425 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9425/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9414 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9414/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8702 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8702/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9469 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9469/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9458 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9458/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9447 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9447/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8735 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8735/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8724 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8724/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8713 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8713/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8768 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8768/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8757 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8757/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8746 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8746/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8779 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8779/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_120 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_120/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_131 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_131/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_142 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_142/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_153 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_153/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_164 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_164/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_175 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_175/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_186 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_186/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_197 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_197/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3020 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3031 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3042 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3053 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3064 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2330 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2341 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2352 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2363 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3075 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3086 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3097 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1640 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1651 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2374 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2385 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2396 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1662 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1673 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1684 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1695 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9992 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9992/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9981 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9981/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9970 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9970/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8009 GRING VDD GND VREF ROW_SEL[80] NB1 VBIAS NB2 pixel_fill_8009/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7319 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7319/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7308 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7308/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6607 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6629 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6618 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5906 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5917 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5928 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5939 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9211 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9211/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9200 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9200/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9255 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9255/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9244 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9244/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9233 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9233/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9222 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9222/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8510 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8510/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9288 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9288/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9277 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9277/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9266 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9266/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8543 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8543/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8532 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8532/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8521 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8521/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9299 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9299/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8576 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8576/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8565 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8565/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8554 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8554/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7842 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7842/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7831 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7831/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7820 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7820/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8598 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8598/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8587 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8587/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7875 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7875/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7864 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7864/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7853 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7853/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7897 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7897/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7886 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7886/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2160 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2171 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2182 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2193 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1492 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1481 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1470 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7127 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7127/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7116 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7116/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7105 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7105/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7149 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7149/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7138 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7138/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6426 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6415 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6404 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6459 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6448 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6437 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_19 GRING VDD GND VREF ROW_SEL[0] NB1 VBIAS NB2 pixel_fill_19/AMP_IN SF_IB
+ pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5703 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5714 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5725 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5736 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5747 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5758 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5769 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9030 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9030/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9063 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9063/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9052 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9052/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9041 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9041/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9096 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9096/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9085 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9085/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9074 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9074/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8351 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8351/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8340 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8340/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8395 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8395/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8384 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8384/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8373 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8373/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8362 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8362/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7650 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7650/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7683 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7683/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7672 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7672/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7661 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7661/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7694 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7694/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6971 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6960 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6993 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6982 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_719 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_719/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_708 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_708/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4309 GRING VDD GND VREF ROW_SEL[43] NB1 VBIAS NB2 pixel_fill_4309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3608 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3619 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2907 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2918 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2929 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6201 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6234 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6223 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6212 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6267 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6256 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6245 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5500 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5511 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5522 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6289 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6278 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4810 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4821 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5533 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5544 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5555 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5566 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4832 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4843 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4854 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5577 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5588 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5599 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4865 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4876 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4887 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4898 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8192 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8192/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8181 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8181/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8170 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8170/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7491 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7491/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7480 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7480/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6790 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_527 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_527/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_516 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_516/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_505 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_505/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_549 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_549/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_538 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_538/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4106 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3405 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4117 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4128 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4139 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3416 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3427 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3438 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2704 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2715 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2726 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2737 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3449 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2748 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2759 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6020 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6031 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6042 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5330 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5341 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6053 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6064 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6075 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5352 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5363 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5374 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6086 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6097 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4640 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4651 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4662 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5385 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5396 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3950 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3961 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4673 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4684 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4695 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3972 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3983 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3994 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9629 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9629/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9618 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9618/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9607 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9607/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8917 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8917/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8906 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8906/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8939 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8939/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8928 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8928/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_302 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_302/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_313 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_313/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_324 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_324/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_335 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_335/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_346 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_346/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_357 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_357/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_368 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_368/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_379 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_379/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3202 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3213 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2501 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2512 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3224 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3235 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3246 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1800 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2523 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2534 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2545 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3257 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3268 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3279 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1811 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1822 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1833 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2556 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2567 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2578 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1844 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1855 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1866 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1877 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2589 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1888 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1899 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_891 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_891/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_880 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_880/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5160 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5171 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5182 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4470 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5193 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4481 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4492 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3780 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3791 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1129 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1118 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1107 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9404 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9404/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9437 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9437/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9426 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9426/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9415 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9415/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9459 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9459/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9448 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9448/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8725 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8725/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8714 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8714/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8703 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8703/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8769 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8769/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8758 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8758/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8747 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8747/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8736 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8736/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_110 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_110/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_121 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_121/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_132 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_132/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_143 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_143/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_154 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_154/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_165 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_165/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_176 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_176/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_187 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_187/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_198 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_198/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3010 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3021 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2320 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3032 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3043 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3054 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3065 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2331 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2342 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2353 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3076 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3087 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3098 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1630 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1641 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2364 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2375 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2386 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1652 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1663 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1674 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1685 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2397 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1696 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9993 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9993/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9982 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9982/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9971 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9971/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9960 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9960/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7309 GRING VDD GND VREF ROW_SEL[73] NB1 VBIAS NB2 pixel_fill_7309/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6608 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6619 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5907 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5918 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5929 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9212 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9212/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9201 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9201/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9245 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9245/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9234 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9234/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9223 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9223/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8500 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8500/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9278 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9278/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9267 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9267/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9256 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9256/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8544 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8544/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8533 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8533/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8522 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8522/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8511 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8511/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9289 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9289/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8577 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8577/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8566 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8566/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8555 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8555/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7832 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7832/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7821 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7821/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7810 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7810/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8599 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8599/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8588 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8588/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7865 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7865/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7854 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7854/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7843 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7843/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7898 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7898/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7887 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7887/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7876 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7876/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2150 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2161 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1460 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2172 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2183 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2194 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1493 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1482 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1471 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9790 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9790/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7128 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7128/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7117 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7117/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7106 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7106/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7139 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7139/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6416 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6405 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6449 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6438 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6427 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5704 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5715 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5726 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5737 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5748 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5759 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9020 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9020/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9053 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9053/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9042 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9042/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9031 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9031/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9097 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9097/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9086 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9086/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9075 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9075/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9064 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9064/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8352 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8352/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8341 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8341/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8330 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8330/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8385 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8385/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8374 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8374/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8363 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8363/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7640 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7640/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8396 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8396/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7684 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7684/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7673 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7673/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7662 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7662/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7651 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7651/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7695 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7695/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6972 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6961 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6950 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6994 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6983 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1290 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_709 GRING VDD GND VREF ROW_SEL[7] NB1 VBIAS NB2 pixel_fill_709/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3609 GRING VDD GND VREF ROW_SEL[36] NB1 VBIAS NB2 pixel_fill_3609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2908 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2919 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6224 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6213 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6202 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6268 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6257 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6246 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6235 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5501 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5512 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5523 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6279 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4800 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4811 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5534 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5545 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5556 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4822 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4833 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4844 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4855 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5567 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5578 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5589 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4866 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4877 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4888 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4899 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8160 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8160/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8193 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8193/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8182 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8182/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8171 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8171/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7492 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7492/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7481 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7481/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7470 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7470/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6780 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6791 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_528 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_528/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_517 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_517/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_506 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_506/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_539 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_539/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4107 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4118 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4129 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3406 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3417 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3428 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3439 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2705 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2716 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2727 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2738 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2749 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6010 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6021 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6032 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6043 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5320 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5331 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6054 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6065 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6076 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5342 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5353 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5364 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6087 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6098 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4630 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4641 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4652 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4663 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5375 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5386 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5397 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3940 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3951 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4674 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4685 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4696 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3962 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3973 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3984 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3995 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9619 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9619/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9608 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9608/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8918 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8918/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8907 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8907/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8929 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8929/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_303 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_303/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_314 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_314/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_325 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_325/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_336 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_336/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_347 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_347/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_358 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_358/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_369 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_369/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3203 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3214 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2502 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3225 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3236 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3247 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2513 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2524 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2535 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3258 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3269 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1801 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1812 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1823 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1834 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2546 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2557 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2568 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2579 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1845 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1856 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1867 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1878 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1889 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_892 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_892/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_881 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_881/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_870 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_870/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5150 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5161 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5172 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5183 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4460 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4471 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5194 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4482 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4493 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3770 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3781 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3792 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1119 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1108 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9427 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9427/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9416 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9416/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9405 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9405/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9449 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9449/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9438 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9438/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8726 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8726/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8715 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8715/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8704 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8704/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8759 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8759/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8748 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8748/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8737 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8737/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_100 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_100/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_111 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_111/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_122 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_122/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_133 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_133/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_144 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_144/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_155 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_155/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_166 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_166/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_177 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_177/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_188 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_188/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_199 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_199/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3000 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3011 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3022 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2310 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3033 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3044 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3055 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2321 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2332 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2343 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2354 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3066 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3077 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3088 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1620 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1631 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1642 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2365 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2376 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2387 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3099 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1653 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1664 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1675 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2398 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1686 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1697 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9950 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9950/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9983 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9983/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9972 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9972/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9961 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9961/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9994 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9994/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4290 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6609 GRING VDD GND VREF ROW_SEL[66] NB1 VBIAS NB2 pixel_fill_6609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5908 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5919 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9202 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9202/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9246 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9246/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9235 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9235/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9224 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9224/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9213 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9213/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8501 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8501/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9279 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9279/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9268 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9268/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9257 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9257/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8534 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8534/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8523 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8523/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8512 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8512/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8567 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8567/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8556 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8556/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8545 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8545/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7833 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7833/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7822 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7822/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7811 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7811/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7800 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7800/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8589 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8589/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8578 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8578/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7866 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7866/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7855 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7855/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7844 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7844/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7899 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7899/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7888 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7888/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7877 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7877/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2140 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2151 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2162 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1450 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2173 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2184 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2195 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1483 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1472 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1461 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1494 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9791 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9791/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9780 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9780/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7118 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7118/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7107 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7107/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7129 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7129/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6417 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6406 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6439 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6428 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5705 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5716 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5727 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5738 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5749 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9021 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9021/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9010 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9010/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9054 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9054/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9043 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9043/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9032 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9032/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9087 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9087/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9076 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9076/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9065 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9065/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8342 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8342/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8331 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8331/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8320 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8320/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9098 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9098/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8386 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8386/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8375 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8375/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8364 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8364/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8353 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8353/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7641 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7641/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7630 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7630/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8397 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8397/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7674 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7674/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7663 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7663/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7652 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7652/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7696 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7696/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7685 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7685/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6962 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6951 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6940 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6995 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6984 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6973 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1291 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1280 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2909 GRING VDD GND VREF ROW_SEL[29] NB1 VBIAS NB2 pixel_fill_2909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6225 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6214 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6203 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6258 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6247 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6236 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5502 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5513 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6269 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4801 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4812 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5524 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5535 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5546 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5557 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4823 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4834 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4845 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5568 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5579 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4856 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4867 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4878 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4889 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8150 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8150/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8194 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8194/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8183 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8183/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8172 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8172/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8161 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8161/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7482 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7482/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7471 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7471/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7460 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7460/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7493 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7493/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6781 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6770 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6792 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_518 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_518/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_507 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_507/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_529 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_529/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4108 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4119 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3407 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3418 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3429 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2706 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2717 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2728 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2739 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6000 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6011 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6022 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6033 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5310 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5321 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6044 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6055 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6066 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4620 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5332 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5343 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5354 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5365 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6077 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6088 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6099 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4631 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4642 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4653 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5376 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5387 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5398 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3930 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3941 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3952 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4664 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4675 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4686 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4697 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3963 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3974 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3985 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3996 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7290 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7290/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9609 GRING VDD GND VREF ROW_SEL[96] NB1 VBIAS NB2 pixel_fill_9609/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8908 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8908/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8919 GRING VDD GND VREF ROW_SEL[89] NB1 VBIAS NB2 pixel_fill_8919/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_304 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_304/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_315 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_315/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_326 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_326/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_337 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_337/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_348 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_348/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_359 GRING VDD GND VREF ROW_SEL[3] NB1 VBIAS NB2 pixel_fill_359/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3204 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2503 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3215 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3226 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3237 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2514 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2525 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2536 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3248 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3259 GRING VDD GND VREF ROW_SEL[32] NB1 VBIAS NB2 pixel_fill_3259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1802 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1813 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1824 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2547 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2558 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2569 GRING VDD GND VREF ROW_SEL[25] NB1 VBIAS NB2 pixel_fill_2569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1835 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1846 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1857 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1868 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1879 GRING VDD GND VREF ROW_SEL[18] NB1 VBIAS NB2 pixel_fill_1879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5140 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_882 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_882/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_871 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_871/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_860 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_860/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5151 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5162 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5173 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_893 GRING VDD GND VREF ROW_SEL[8] NB1 VBIAS NB2 pixel_fill_893/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4450 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4461 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5184 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5195 GRING VDD GND VREF ROW_SEL[51] NB1 VBIAS NB2 pixel_fill_5195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3760 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4472 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4483 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4494 GRING VDD GND VREF ROW_SEL[44] NB1 VBIAS NB2 pixel_fill_4494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3771 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3782 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3793 GRING VDD GND VREF ROW_SEL[37] NB1 VBIAS NB2 pixel_fill_3793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1109 GRING VDD GND VREF ROW_SEL[11] NB1 VBIAS NB2 pixel_fill_1109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9428 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9428/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9417 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9417/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9406 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9406/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9439 GRING VDD GND VREF ROW_SEL[94] NB1 VBIAS NB2 pixel_fill_9439/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8716 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8716/AMP_IN
+ SF_IB pixel_fill_16/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8705 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8705/AMP_IN
+ SF_IB pixel_fill_5/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8749 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8749/AMP_IN
+ SF_IB pixel_fill_49/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8738 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8738/AMP_IN
+ SF_IB pixel_fill_38/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8727 GRING VDD GND VREF ROW_SEL[87] NB1 VBIAS NB2 pixel_fill_8727/AMP_IN
+ SF_IB pixel_fill_27/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_101 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_101/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_112 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_112/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_123 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_123/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_134 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_134/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_145 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_145/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_156 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_156/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_167 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_167/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_178 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_178/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_189 GRING VDD GND VREF ROW_SEL[1] NB1 VBIAS NB2 pixel_fill_189/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3001 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3012 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2300 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2311 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3023 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3034 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3045 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3056 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2322 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2333 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2344 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3067 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3078 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3089 GRING VDD GND VREF ROW_SEL[30] NB1 VBIAS NB2 pixel_fill_3089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1610 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1621 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1632 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2355 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2366 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2377 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1643 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1654 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1665 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1676 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2388 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2399 GRING VDD GND VREF ROW_SEL[23] NB1 VBIAS NB2 pixel_fill_2399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1687 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1698 GRING VDD GND VREF ROW_SEL[16] NB1 VBIAS NB2 pixel_fill_1698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9940 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9940/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9984 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9984/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9973 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9973/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9962 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9962/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9951 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9951/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9995 GRING VDD GND VREF ROW_SEL[99] NB1 VBIAS NB2 pixel_fill_9995/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_690 GRING VDD GND VREF ROW_SEL[6] NB1 VBIAS NB2 pixel_fill_690/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4280 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4291 GRING VDD GND VREF ROW_SEL[42] NB1 VBIAS NB2 pixel_fill_4291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3590 GRING VDD GND VREF ROW_SEL[35] NB1 VBIAS NB2 pixel_fill_3590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5909 GRING VDD GND VREF ROW_SEL[59] NB1 VBIAS NB2 pixel_fill_5909/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9203 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9203/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9236 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9236/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9225 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9225/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9214 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9214/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9269 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9269/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9258 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9258/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9247 GRING VDD GND VREF ROW_SEL[92] NB1 VBIAS NB2 pixel_fill_9247/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8535 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8535/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8524 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8524/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8513 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8513/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8502 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8502/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8568 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8568/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8557 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8557/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8546 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8546/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7823 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7823/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7812 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7812/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7801 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7801/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8579 GRING VDD GND VREF ROW_SEL[85] NB1 VBIAS NB2 pixel_fill_8579/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7856 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7856/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7845 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7845/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7834 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7834/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7889 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7889/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7878 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7878/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7867 GRING VDD GND VREF ROW_SEL[78] NB1 VBIAS NB2 pixel_fill_7867/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2130 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2130/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2141 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2141/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2152 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2152/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1451 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1451/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1440 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1440/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2163 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2163/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2174 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2174/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2185 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2185/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2196 GRING VDD GND VREF ROW_SEL[21] NB1 VBIAS NB2 pixel_fill_2196/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1484 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1484/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1473 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1473/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1462 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1462/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1495 GRING VDD GND VREF ROW_SEL[14] NB1 VBIAS NB2 pixel_fill_1495/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9792 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9792/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9781 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9781/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9770 GRING VDD GND VREF ROW_SEL[97] NB1 VBIAS NB2 pixel_fill_9770/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7119 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7119/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7108 GRING VDD GND VREF ROW_SEL[71] NB1 VBIAS NB2 pixel_fill_7108/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6407 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6407/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6429 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6429/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6418 GRING VDD GND VREF ROW_SEL[64] NB1 VBIAS NB2 pixel_fill_6418/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5706 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5706/AMP_IN
+ SF_IB pixel_fill_6/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5717 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5717/AMP_IN
+ SF_IB pixel_fill_17/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5728 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5728/AMP_IN
+ SF_IB pixel_fill_28/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5739 GRING VDD GND VREF ROW_SEL[57] NB1 VBIAS NB2 pixel_fill_5739/AMP_IN
+ SF_IB pixel_fill_39/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9011 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9011/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9000 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9000/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9044 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9044/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9033 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9033/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9022 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9022/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9088 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9088/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9077 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9077/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9066 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9066/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9055 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9055/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8343 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8343/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8332 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8332/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8321 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8321/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8310 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8310/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_9099 GRING VDD GND VREF ROW_SEL[90] NB1 VBIAS NB2 pixel_fill_9099/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8376 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8376/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8365 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8365/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8354 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8354/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7631 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7631/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7620 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7620/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8398 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8398/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8387 GRING VDD GND VREF ROW_SEL[83] NB1 VBIAS NB2 pixel_fill_8387/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7675 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7675/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7664 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7664/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7653 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7653/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7642 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7642/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6930 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6930/AMP_IN
+ SF_IB pixel_fill_30/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7697 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7697/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7686 GRING VDD GND VREF ROW_SEL[76] NB1 VBIAS NB2 pixel_fill_7686/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6963 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6963/AMP_IN
+ SF_IB pixel_fill_63/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6952 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6952/AMP_IN
+ SF_IB pixel_fill_52/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6941 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6941/AMP_IN
+ SF_IB pixel_fill_41/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6996 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6996/AMP_IN
+ SF_IB pixel_fill_96/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6985 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6985/AMP_IN
+ SF_IB pixel_fill_85/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6974 GRING VDD GND VREF ROW_SEL[69] NB1 VBIAS NB2 pixel_fill_6974/AMP_IN
+ SF_IB pixel_fill_74/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1292 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1292/AMP_IN
+ SF_IB pixel_fill_92/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1281 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1281/AMP_IN
+ SF_IB pixel_fill_81/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_1270 GRING VDD GND VREF ROW_SEL[12] NB1 VBIAS NB2 pixel_fill_1270/AMP_IN
+ SF_IB pixel_fill_70/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6215 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6215/AMP_IN
+ SF_IB pixel_fill_15/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6204 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6204/AMP_IN
+ SF_IB pixel_fill_4/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6259 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6259/AMP_IN
+ SF_IB pixel_fill_59/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6248 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6248/AMP_IN
+ SF_IB pixel_fill_48/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6237 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6237/AMP_IN
+ SF_IB pixel_fill_37/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6226 GRING VDD GND VREF ROW_SEL[62] NB1 VBIAS NB2 pixel_fill_6226/AMP_IN
+ SF_IB pixel_fill_26/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5503 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5503/AMP_IN
+ SF_IB pixel_fill_3/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5514 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5514/AMP_IN
+ SF_IB pixel_fill_14/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4802 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4802/AMP_IN
+ SF_IB pixel_fill_2/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5525 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5525/AMP_IN
+ SF_IB pixel_fill_25/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5536 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5536/AMP_IN
+ SF_IB pixel_fill_36/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5547 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5547/AMP_IN
+ SF_IB pixel_fill_47/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4813 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4813/AMP_IN
+ SF_IB pixel_fill_13/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4824 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4824/AMP_IN
+ SF_IB pixel_fill_24/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4835 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4835/AMP_IN
+ SF_IB pixel_fill_35/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4846 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4846/AMP_IN
+ SF_IB pixel_fill_46/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5558 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5558/AMP_IN
+ SF_IB pixel_fill_58/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5569 GRING VDD GND VREF ROW_SEL[55] NB1 VBIAS NB2 pixel_fill_5569/AMP_IN
+ SF_IB pixel_fill_69/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4857 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4857/AMP_IN
+ SF_IB pixel_fill_57/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4868 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4868/AMP_IN
+ SF_IB pixel_fill_68/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4879 GRING VDD GND VREF ROW_SEL[48] NB1 VBIAS NB2 pixel_fill_4879/AMP_IN
+ SF_IB pixel_fill_79/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8151 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8151/AMP_IN
+ SF_IB pixel_fill_51/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8140 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8140/AMP_IN
+ SF_IB pixel_fill_40/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8184 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8184/AMP_IN
+ SF_IB pixel_fill_84/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8173 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8173/AMP_IN
+ SF_IB pixel_fill_73/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8162 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8162/AMP_IN
+ SF_IB pixel_fill_62/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_8195 GRING VDD GND VREF ROW_SEL[81] NB1 VBIAS NB2 pixel_fill_8195/AMP_IN
+ SF_IB pixel_fill_95/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7483 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7483/AMP_IN
+ SF_IB pixel_fill_83/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7472 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7472/AMP_IN
+ SF_IB pixel_fill_72/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7461 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7461/AMP_IN
+ SF_IB pixel_fill_61/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7450 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7450/AMP_IN
+ SF_IB pixel_fill_50/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7494 GRING VDD GND VREF ROW_SEL[74] NB1 VBIAS NB2 pixel_fill_7494/AMP_IN
+ SF_IB pixel_fill_94/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6771 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6771/AMP_IN
+ SF_IB pixel_fill_71/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6760 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6760/AMP_IN
+ SF_IB pixel_fill_60/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6793 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6793/AMP_IN
+ SF_IB pixel_fill_93/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6782 GRING VDD GND VREF ROW_SEL[67] NB1 VBIAS NB2 pixel_fill_6782/AMP_IN
+ SF_IB pixel_fill_82/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_519 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_519/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_508 GRING VDD GND VREF ROW_SEL[5] NB1 VBIAS NB2 pixel_fill_508/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4109 GRING VDD GND VREF ROW_SEL[41] NB1 VBIAS NB2 pixel_fill_4109/AMP_IN
+ SF_IB pixel_fill_9/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3408 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3408/AMP_IN
+ SF_IB pixel_fill_8/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3419 GRING VDD GND VREF ROW_SEL[34] NB1 VBIAS NB2 pixel_fill_3419/AMP_IN
+ SF_IB pixel_fill_19/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2707 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2707/AMP_IN
+ SF_IB pixel_fill_7/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2718 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2718/AMP_IN
+ SF_IB pixel_fill_18/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_2729 GRING VDD GND VREF ROW_SEL[27] NB1 VBIAS NB2 pixel_fill_2729/AMP_IN
+ SF_IB pixel_fill_29/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6001 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6001/AMP_IN
+ SF_IB pixel_fill_901/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6012 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6012/AMP_IN
+ SF_IB pixel_fill_12/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6023 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6023/AMP_IN
+ SF_IB pixel_fill_23/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6034 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6034/AMP_IN
+ SF_IB pixel_fill_34/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5300 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5300/AMP_IN
+ SF_IB pixel_fill_900/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5311 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5311/AMP_IN
+ SF_IB pixel_fill_11/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5322 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5322/AMP_IN
+ SF_IB pixel_fill_22/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6045 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6045/AMP_IN
+ SF_IB pixel_fill_45/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6056 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6056/AMP_IN
+ SF_IB pixel_fill_56/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6067 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6067/AMP_IN
+ SF_IB pixel_fill_67/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4610 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4610/AMP_IN
+ SF_IB pixel_fill_10/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5333 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5333/AMP_IN
+ SF_IB pixel_fill_33/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5344 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5344/AMP_IN
+ SF_IB pixel_fill_44/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5355 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5355/AMP_IN
+ SF_IB pixel_fill_55/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6078 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6078/AMP_IN
+ SF_IB pixel_fill_78/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6089 GRING VDD GND VREF ROW_SEL[60] NB1 VBIAS NB2 pixel_fill_6089/AMP_IN
+ SF_IB pixel_fill_89/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4621 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4621/AMP_IN
+ SF_IB pixel_fill_21/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4632 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4632/AMP_IN
+ SF_IB pixel_fill_32/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4643 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4643/AMP_IN
+ SF_IB pixel_fill_43/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4654 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4654/AMP_IN
+ SF_IB pixel_fill_54/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5366 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5366/AMP_IN
+ SF_IB pixel_fill_66/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5377 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5377/AMP_IN
+ SF_IB pixel_fill_77/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5388 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5388/AMP_IN
+ SF_IB pixel_fill_88/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_5399 GRING VDD GND VREF ROW_SEL[53] NB1 VBIAS NB2 pixel_fill_5399/AMP_IN
+ SF_IB pixel_fill_99/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3920 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3920/AMP_IN
+ SF_IB pixel_fill_20/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3931 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3931/AMP_IN
+ SF_IB pixel_fill_31/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3942 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3942/AMP_IN
+ SF_IB pixel_fill_42/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4665 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4665/AMP_IN
+ SF_IB pixel_fill_65/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4676 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4676/AMP_IN
+ SF_IB pixel_fill_76/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4687 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4687/AMP_IN
+ SF_IB pixel_fill_87/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3953 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3953/AMP_IN
+ SF_IB pixel_fill_53/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3964 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3964/AMP_IN
+ SF_IB pixel_fill_64/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3975 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3975/AMP_IN
+ SF_IB pixel_fill_75/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_4698 GRING VDD GND VREF ROW_SEL[46] NB1 VBIAS NB2 pixel_fill_4698/AMP_IN
+ SF_IB pixel_fill_98/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3986 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3986/AMP_IN
+ SF_IB pixel_fill_86/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_3997 GRING VDD GND VREF ROW_SEL[39] NB1 VBIAS NB2 pixel_fill_3997/AMP_IN
+ SF_IB pixel_fill_97/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7291 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7291/AMP_IN
+ SF_IB pixel_fill_91/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_7280 GRING VDD GND VREF ROW_SEL[72] NB1 VBIAS NB2 pixel_fill_7280/AMP_IN
+ SF_IB pixel_fill_80/PIX_OUT CSA_VREF pixel_fill
Xpixel_fill_6590 GRING VDD GND VREF ROW_SEL[65] NB1 VBIAS NB2 pixel_fill_6590/AMP_IN
+ SF_IB pixel_fill_90/PIX_OUT CSA_VREF pixel_fill
X0 pixel_fill_83/PIX_OUT COL_SEL[83] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X1 pixel_fill_79/PIX_OUT COL_SEL[79] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X2 pixel_fill_75/PIX_OUT COL_SEL[75] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X3 pixel_fill_71/PIX_OUT COL_SEL[71] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X4 pixel_fill_67/PIX_OUT COL_SEL[67] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X5 pixel_fill_26/PIX_OUT COL_SEL[26] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X6 pixel_fill_64/PIX_OUT COL_SEL[64] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X7 pixel_fill_22/PIX_OUT COL_SEL[22] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X8 pixel_fill_18/PIX_OUT COL_SEL[18] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X9 pixel_fill_60/PIX_OUT COL_SEL[60] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X10 pixel_fill_14/PIX_OUT COL_SEL[14] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X11 pixel_fill_10/PIX_OUT COL_SEL[10] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X12 pixel_fill_86/PIX_OUT COL_SEL[86] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X13 pixel_fill_82/PIX_OUT COL_SEL[82] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X14 pixel_fill_78/PIX_OUT COL_SEL[78] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X15 pixel_fill_74/PIX_OUT COL_SEL[74] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X16 pixel_fill_70/PIX_OUT COL_SEL[70] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X17 pixel_fill_33/PIX_OUT COL_SEL[33] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X18 pixel_fill_29/PIX_OUT COL_SEL[29] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X19 pixel_fill_25/PIX_OUT COL_SEL[25] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X20 pixel_fill_21/PIX_OUT COL_SEL[21] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X21 pixel_fill_17/PIX_OUT COL_SEL[17] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X22 pixel_fill_93/PIX_OUT COL_SEL[93] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X23 pixel_fill_89/PIX_OUT COL_SEL[89] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X24 pixel_fill_85/PIX_OUT COL_SEL[85] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X25 pixel_fill_81/PIX_OUT COL_SEL[81] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X26 pixel_fill_77/PIX_OUT COL_SEL[77] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X27 pixel_fill_36/PIX_OUT COL_SEL[36] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X28 pixel_fill_32/PIX_OUT COL_SEL[32] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X29 pixel_fill_28/PIX_OUT COL_SEL[28] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X30 pixel_fill_24/PIX_OUT COL_SEL[24] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X31 pixel_fill_20/PIX_OUT COL_SEL[20] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X32 pixel_fill_3/PIX_OUT COL_SEL[3] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X33 pixel_fill_96/PIX_OUT COL_SEL[96] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X34 pixel_fill_92/PIX_OUT COL_SEL[92] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X35 pixel_fill_88/PIX_OUT COL_SEL[88] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X36 pixel_fill_84/PIX_OUT COL_SEL[84] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X37 pixel_fill_80/PIX_OUT COL_SEL[80] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X38 pixel_fill_43/PIX_OUT COL_SEL[43] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X39 pixel_fill_900/PIX_OUT COL_SEL[0] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X40 pixel_fill_39/PIX_OUT COL_SEL[39] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X41 pixel_fill_35/PIX_OUT COL_SEL[35] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X42 pixel_fill_31/PIX_OUT COL_SEL[31] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X43 pixel_fill_27/PIX_OUT COL_SEL[27] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X44 pixel_fill_2/PIX_OUT COL_SEL[2] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X45 pixel_fill_99/PIX_OUT COL_SEL[99] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X46 pixel_fill_95/PIX_OUT COL_SEL[95] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X47 pixel_fill_91/PIX_OUT COL_SEL[91] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X48 pixel_fill_87/PIX_OUT COL_SEL[87] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X49 pixel_fill_46/PIX_OUT COL_SEL[46] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X50 pixel_fill_42/PIX_OUT COL_SEL[42] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X51 pixel_fill_38/PIX_OUT COL_SEL[38] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X52 pixel_fill_34/PIX_OUT COL_SEL[34] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X53 pixel_fill_30/PIX_OUT COL_SEL[30] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X54 pixel_fill_901/PIX_OUT COL_SEL[1] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X55 pixel_fill_98/PIX_OUT COL_SEL[98] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X56 pixel_fill_94/PIX_OUT COL_SEL[94] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X57 pixel_fill_90/PIX_OUT COL_SEL[90] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X58 pixel_fill_53/PIX_OUT COL_SEL[53] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X59 pixel_fill_49/PIX_OUT COL_SEL[49] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X60 pixel_fill_45/PIX_OUT COL_SEL[45] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X61 pixel_fill_41/PIX_OUT COL_SEL[41] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X62 pixel_fill_37/PIX_OUT COL_SEL[37] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X63 pixel_fill_97/PIX_OUT COL_SEL[97] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X64 pixel_fill_56/PIX_OUT COL_SEL[56] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X65 pixel_fill_52/PIX_OUT COL_SEL[52] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X66 pixel_fill_6/PIX_OUT COL_SEL[6] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X67 pixel_fill_48/PIX_OUT COL_SEL[48] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X68 pixel_fill_44/PIX_OUT COL_SEL[44] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X69 pixel_fill_40/PIX_OUT COL_SEL[40] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X70 pixel_fill_63/PIX_OUT COL_SEL[63] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X71 pixel_fill_59/PIX_OUT COL_SEL[59] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X72 pixel_fill_55/PIX_OUT COL_SEL[55] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X73 pixel_fill_13/PIX_OUT COL_SEL[13] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X74 pixel_fill_9/PIX_OUT COL_SEL[9] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X75 pixel_fill_51/PIX_OUT COL_SEL[51] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X76 pixel_fill_5/PIX_OUT COL_SEL[5] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X77 pixel_fill_47/PIX_OUT COL_SEL[47] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X78 pixel_fill_73/PIX_OUT COL_SEL[73] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X79 pixel_fill_69/PIX_OUT COL_SEL[69] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X80 pixel_fill_66/PIX_OUT COL_SEL[66] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X81 pixel_fill_62/PIX_OUT COL_SEL[62] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X82 pixel_fill_16/PIX_OUT COL_SEL[16] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X83 pixel_fill_12/PIX_OUT COL_SEL[12] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X84 pixel_fill_58/PIX_OUT COL_SEL[58] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X85 pixel_fill_54/PIX_OUT COL_SEL[54] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X86 pixel_fill_8/PIX_OUT COL_SEL[8] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X87 pixel_fill_50/PIX_OUT COL_SEL[50] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X88 pixel_fill_4/PIX_OUT COL_SEL[4] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X89 pixel_fill_76/PIX_OUT COL_SEL[76] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X90 pixel_fill_72/PIX_OUT COL_SEL[72] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X91 pixel_fill_68/PIX_OUT COL_SEL[68] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X92 pixel_fill_23/PIX_OUT COL_SEL[23] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X93 pixel_fill_19/PIX_OUT COL_SEL[19] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X94 pixel_fill_65/PIX_OUT COL_SEL[65] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X95 pixel_fill_61/PIX_OUT COL_SEL[61] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X96 pixel_fill_15/PIX_OUT COL_SEL[15] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X97 pixel_fill_11/PIX_OUT COL_SEL[11] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X98 pixel_fill_57/PIX_OUT COL_SEL[57] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
X99 pixel_fill_7/PIX_OUT COL_SEL[7] ARRAY_OUT GND sky130_fd_pr__nfet_01v8_lvt ad=4 pd=17 as=3.2 ps=16.8 w=8 l=2
.ends

.subckt array_SR VDD COL_ENA COL_RST COL_DIN COL_CLK CSA_VREF ARRAY_OUT NB1 NB2 VBIAS
+ VREF SF_IB ROW_DIN gring ROW_CLK ROW_RST ROW_ENA GND
Xshift_registerC_0 shift_registerC_0/COL_SEL[0] shift_registerC_0/COL_SEL[10] shift_registerC_0/COL_SEL[11]
+ shift_registerC_0/COL_SEL[12] shift_registerC_0/COL_SEL[13] shift_registerC_0/COL_SEL[14]
+ shift_registerC_0/COL_SEL[15] shift_registerC_0/COL_SEL[16] shift_registerC_0/COL_SEL[17]
+ shift_registerC_0/COL_SEL[18] shift_registerC_0/COL_SEL[19] shift_registerC_0/COL_SEL[1]
+ shift_registerC_0/COL_SEL[20] shift_registerC_0/COL_SEL[21] shift_registerC_0/COL_SEL[22]
+ shift_registerC_0/COL_SEL[23] shift_registerC_0/COL_SEL[24] shift_registerC_0/COL_SEL[25]
+ shift_registerC_0/COL_SEL[26] shift_registerC_0/COL_SEL[27] shift_registerC_0/COL_SEL[28]
+ shift_registerC_0/COL_SEL[29] shift_registerC_0/COL_SEL[2] shift_registerC_0/COL_SEL[30]
+ shift_registerC_0/COL_SEL[31] shift_registerC_0/COL_SEL[32] shift_registerC_0/COL_SEL[33]
+ shift_registerC_0/COL_SEL[34] shift_registerC_0/COL_SEL[35] shift_registerC_0/COL_SEL[36]
+ shift_registerC_0/COL_SEL[37] shift_registerC_0/COL_SEL[38] shift_registerC_0/COL_SEL[39]
+ shift_registerC_0/COL_SEL[3] shift_registerC_0/COL_SEL[40] shift_registerC_0/COL_SEL[41]
+ shift_registerC_0/COL_SEL[42] shift_registerC_0/COL_SEL[43] shift_registerC_0/COL_SEL[44]
+ shift_registerC_0/COL_SEL[45] shift_registerC_0/COL_SEL[46] shift_registerC_0/COL_SEL[47]
+ shift_registerC_0/COL_SEL[48] shift_registerC_0/COL_SEL[49] shift_registerC_0/COL_SEL[4]
+ shift_registerC_0/COL_SEL[50] shift_registerC_0/COL_SEL[51] shift_registerC_0/COL_SEL[52]
+ shift_registerC_0/COL_SEL[53] shift_registerC_0/COL_SEL[54] shift_registerC_0/COL_SEL[55]
+ shift_registerC_0/COL_SEL[56] shift_registerC_0/COL_SEL[57] shift_registerC_0/COL_SEL[58]
+ shift_registerC_0/COL_SEL[59] shift_registerC_0/COL_SEL[5] shift_registerC_0/COL_SEL[60]
+ shift_registerC_0/COL_SEL[61] shift_registerC_0/COL_SEL[62] shift_registerC_0/COL_SEL[63]
+ shift_registerC_0/COL_SEL[64] shift_registerC_0/COL_SEL[65] shift_registerC_0/COL_SEL[66]
+ shift_registerC_0/COL_SEL[67] shift_registerC_0/COL_SEL[68] shift_registerC_0/COL_SEL[69]
+ shift_registerC_0/COL_SEL[6] shift_registerC_0/COL_SEL[70] shift_registerC_0/COL_SEL[71]
+ shift_registerC_0/COL_SEL[72] shift_registerC_0/COL_SEL[73] shift_registerC_0/COL_SEL[74]
+ shift_registerC_0/COL_SEL[75] shift_registerC_0/COL_SEL[76] shift_registerC_0/COL_SEL[77]
+ shift_registerC_0/COL_SEL[78] shift_registerC_0/COL_SEL[79] shift_registerC_0/COL_SEL[7]
+ shift_registerC_0/COL_SEL[80] shift_registerC_0/COL_SEL[81] shift_registerC_0/COL_SEL[82]
+ shift_registerC_0/COL_SEL[83] shift_registerC_0/COL_SEL[84] shift_registerC_0/COL_SEL[85]
+ shift_registerC_0/COL_SEL[86] shift_registerC_0/COL_SEL[87] shift_registerC_0/COL_SEL[88]
+ shift_registerC_0/COL_SEL[89] shift_registerC_0/COL_SEL[8] shift_registerC_0/COL_SEL[90]
+ shift_registerC_0/COL_SEL[91] shift_registerC_0/COL_SEL[92] shift_registerC_0/COL_SEL[93]
+ shift_registerC_0/COL_SEL[94] shift_registerC_0/COL_SEL[95] shift_registerC_0/COL_SEL[96]
+ shift_registerC_0/COL_SEL[97] shift_registerC_0/COL_SEL[98] shift_registerC_0/COL_SEL[99]
+ shift_registerC_0/COL_SEL[9] COL_CLK COL_DIN shift_registerC_0/data_out COL_ENA
+ COL_RST VDD GND shift_registerC
Xshift_registerC_1 shift_registerC_1/COL_SEL[0] shift_registerC_1/COL_SEL[10] shift_registerC_1/COL_SEL[11]
+ shift_registerC_1/COL_SEL[12] shift_registerC_1/COL_SEL[13] shift_registerC_1/COL_SEL[14]
+ shift_registerC_1/COL_SEL[15] shift_registerC_1/COL_SEL[16] shift_registerC_1/COL_SEL[17]
+ shift_registerC_1/COL_SEL[18] shift_registerC_1/COL_SEL[19] shift_registerC_1/COL_SEL[1]
+ shift_registerC_1/COL_SEL[20] shift_registerC_1/COL_SEL[21] shift_registerC_1/COL_SEL[22]
+ shift_registerC_1/COL_SEL[23] shift_registerC_1/COL_SEL[24] shift_registerC_1/COL_SEL[25]
+ shift_registerC_1/COL_SEL[26] shift_registerC_1/COL_SEL[27] shift_registerC_1/COL_SEL[28]
+ shift_registerC_1/COL_SEL[29] shift_registerC_1/COL_SEL[2] shift_registerC_1/COL_SEL[30]
+ shift_registerC_1/COL_SEL[31] shift_registerC_1/COL_SEL[32] shift_registerC_1/COL_SEL[33]
+ shift_registerC_1/COL_SEL[34] shift_registerC_1/COL_SEL[35] shift_registerC_1/COL_SEL[36]
+ shift_registerC_1/COL_SEL[37] shift_registerC_1/COL_SEL[38] shift_registerC_1/COL_SEL[39]
+ shift_registerC_1/COL_SEL[3] shift_registerC_1/COL_SEL[40] shift_registerC_1/COL_SEL[41]
+ shift_registerC_1/COL_SEL[42] shift_registerC_1/COL_SEL[43] shift_registerC_1/COL_SEL[44]
+ shift_registerC_1/COL_SEL[45] shift_registerC_1/COL_SEL[46] shift_registerC_1/COL_SEL[47]
+ shift_registerC_1/COL_SEL[48] shift_registerC_1/COL_SEL[49] shift_registerC_1/COL_SEL[4]
+ shift_registerC_1/COL_SEL[50] shift_registerC_1/COL_SEL[51] shift_registerC_1/COL_SEL[52]
+ shift_registerC_1/COL_SEL[53] shift_registerC_1/COL_SEL[54] shift_registerC_1/COL_SEL[55]
+ shift_registerC_1/COL_SEL[56] shift_registerC_1/COL_SEL[57] shift_registerC_1/COL_SEL[58]
+ shift_registerC_1/COL_SEL[59] shift_registerC_1/COL_SEL[5] shift_registerC_1/COL_SEL[60]
+ shift_registerC_1/COL_SEL[61] shift_registerC_1/COL_SEL[62] shift_registerC_1/COL_SEL[63]
+ shift_registerC_1/COL_SEL[64] shift_registerC_1/COL_SEL[65] shift_registerC_1/COL_SEL[66]
+ shift_registerC_1/COL_SEL[67] shift_registerC_1/COL_SEL[68] shift_registerC_1/COL_SEL[69]
+ shift_registerC_1/COL_SEL[6] shift_registerC_1/COL_SEL[70] shift_registerC_1/COL_SEL[71]
+ shift_registerC_1/COL_SEL[72] shift_registerC_1/COL_SEL[73] shift_registerC_1/COL_SEL[74]
+ shift_registerC_1/COL_SEL[75] shift_registerC_1/COL_SEL[76] shift_registerC_1/COL_SEL[77]
+ shift_registerC_1/COL_SEL[78] shift_registerC_1/COL_SEL[79] shift_registerC_1/COL_SEL[7]
+ shift_registerC_1/COL_SEL[80] shift_registerC_1/COL_SEL[81] shift_registerC_1/COL_SEL[82]
+ shift_registerC_1/COL_SEL[83] shift_registerC_1/COL_SEL[84] shift_registerC_1/COL_SEL[85]
+ shift_registerC_1/COL_SEL[86] shift_registerC_1/COL_SEL[87] shift_registerC_1/COL_SEL[88]
+ shift_registerC_1/COL_SEL[89] shift_registerC_1/COL_SEL[8] shift_registerC_1/COL_SEL[90]
+ shift_registerC_1/COL_SEL[91] shift_registerC_1/COL_SEL[92] shift_registerC_1/COL_SEL[93]
+ shift_registerC_1/COL_SEL[94] shift_registerC_1/COL_SEL[95] shift_registerC_1/COL_SEL[96]
+ shift_registerC_1/COL_SEL[97] shift_registerC_1/COL_SEL[98] shift_registerC_1/COL_SEL[99]
+ shift_registerC_1/COL_SEL[9] ROW_CLK ROW_DIN shift_registerC_1/data_out ROW_ENA
+ ROW_RST VDD GND shift_registerC
Xpixel_array100x100_fill_0 VBIAS VREF NB2 VDD NB1 shift_registerC_1/COL_SEL[0] gring
+ shift_registerC_1/COL_SEL[1] shift_registerC_1/COL_SEL[2] shift_registerC_1/COL_SEL[3]
+ shift_registerC_1/COL_SEL[4] shift_registerC_1/COL_SEL[5] shift_registerC_1/COL_SEL[6]
+ shift_registerC_1/COL_SEL[7] shift_registerC_1/COL_SEL[8] shift_registerC_1/COL_SEL[9]
+ shift_registerC_1/COL_SEL[10] shift_registerC_1/COL_SEL[11] shift_registerC_1/COL_SEL[12]
+ shift_registerC_1/COL_SEL[13] shift_registerC_1/COL_SEL[14] shift_registerC_1/COL_SEL[15]
+ shift_registerC_1/COL_SEL[16] shift_registerC_1/COL_SEL[17] shift_registerC_1/COL_SEL[18]
+ shift_registerC_1/COL_SEL[19] shift_registerC_1/COL_SEL[20] shift_registerC_1/COL_SEL[21]
+ shift_registerC_1/COL_SEL[22] shift_registerC_1/COL_SEL[23] shift_registerC_1/COL_SEL[24]
+ shift_registerC_1/COL_SEL[25] shift_registerC_1/COL_SEL[26] shift_registerC_1/COL_SEL[27]
+ shift_registerC_1/COL_SEL[28] shift_registerC_1/COL_SEL[29] shift_registerC_1/COL_SEL[30]
+ shift_registerC_1/COL_SEL[31] shift_registerC_1/COL_SEL[32] shift_registerC_1/COL_SEL[33]
+ shift_registerC_1/COL_SEL[34] shift_registerC_1/COL_SEL[35] shift_registerC_1/COL_SEL[36]
+ shift_registerC_1/COL_SEL[37] shift_registerC_1/COL_SEL[38] shift_registerC_1/COL_SEL[39]
+ shift_registerC_1/COL_SEL[40] shift_registerC_1/COL_SEL[41] shift_registerC_1/COL_SEL[42]
+ shift_registerC_1/COL_SEL[43] shift_registerC_1/COL_SEL[44] shift_registerC_1/COL_SEL[45]
+ shift_registerC_1/COL_SEL[46] shift_registerC_1/COL_SEL[47] shift_registerC_1/COL_SEL[48]
+ shift_registerC_1/COL_SEL[49] shift_registerC_1/COL_SEL[50] shift_registerC_1/COL_SEL[51]
+ shift_registerC_1/COL_SEL[52] shift_registerC_1/COL_SEL[53] shift_registerC_1/COL_SEL[54]
+ shift_registerC_1/COL_SEL[55] shift_registerC_1/COL_SEL[56] shift_registerC_1/COL_SEL[57]
+ shift_registerC_1/COL_SEL[58] shift_registerC_1/COL_SEL[59] shift_registerC_1/COL_SEL[60]
+ shift_registerC_1/COL_SEL[61] shift_registerC_1/COL_SEL[62] shift_registerC_1/COL_SEL[63]
+ shift_registerC_1/COL_SEL[64] shift_registerC_1/COL_SEL[65] shift_registerC_1/COL_SEL[66]
+ shift_registerC_1/COL_SEL[67] shift_registerC_1/COL_SEL[68] shift_registerC_1/COL_SEL[69]
+ shift_registerC_1/COL_SEL[70] shift_registerC_1/COL_SEL[71] shift_registerC_1/COL_SEL[72]
+ shift_registerC_1/COL_SEL[73] shift_registerC_1/COL_SEL[74] shift_registerC_1/COL_SEL[75]
+ shift_registerC_1/COL_SEL[76] shift_registerC_1/COL_SEL[77] shift_registerC_1/COL_SEL[78]
+ shift_registerC_1/COL_SEL[79] shift_registerC_1/COL_SEL[80] shift_registerC_1/COL_SEL[81]
+ shift_registerC_1/COL_SEL[82] shift_registerC_1/COL_SEL[83] shift_registerC_1/COL_SEL[84]
+ shift_registerC_1/COL_SEL[85] shift_registerC_1/COL_SEL[86] shift_registerC_1/COL_SEL[87]
+ shift_registerC_1/COL_SEL[88] shift_registerC_1/COL_SEL[89] shift_registerC_1/COL_SEL[90]
+ shift_registerC_1/COL_SEL[91] shift_registerC_1/COL_SEL[92] shift_registerC_1/COL_SEL[93]
+ shift_registerC_1/COL_SEL[94] shift_registerC_1/COL_SEL[95] shift_registerC_1/COL_SEL[96]
+ shift_registerC_1/COL_SEL[97] shift_registerC_1/COL_SEL[98] shift_registerC_0/COL_SEL[0]
+ CSA_VREF shift_registerC_1/COL_SEL[99] shift_registerC_0/COL_SEL[1] shift_registerC_0/COL_SEL[2]
+ shift_registerC_0/COL_SEL[3] shift_registerC_0/COL_SEL[4] shift_registerC_0/COL_SEL[5]
+ shift_registerC_0/COL_SEL[6] shift_registerC_0/COL_SEL[7] shift_registerC_0/COL_SEL[8]
+ shift_registerC_0/COL_SEL[9] shift_registerC_0/COL_SEL[10] shift_registerC_0/COL_SEL[11]
+ shift_registerC_0/COL_SEL[12] shift_registerC_0/COL_SEL[13] shift_registerC_0/COL_SEL[14]
+ shift_registerC_0/COL_SEL[15] shift_registerC_0/COL_SEL[16] shift_registerC_0/COL_SEL[17]
+ shift_registerC_0/COL_SEL[18] shift_registerC_0/COL_SEL[19] shift_registerC_0/COL_SEL[20]
+ shift_registerC_0/COL_SEL[21] shift_registerC_0/COL_SEL[22] shift_registerC_0/COL_SEL[23]
+ shift_registerC_0/COL_SEL[24] shift_registerC_0/COL_SEL[25] shift_registerC_0/COL_SEL[26]
+ shift_registerC_0/COL_SEL[27] shift_registerC_0/COL_SEL[28] shift_registerC_0/COL_SEL[29]
+ shift_registerC_0/COL_SEL[30] shift_registerC_0/COL_SEL[31] shift_registerC_0/COL_SEL[32]
+ shift_registerC_0/COL_SEL[33] shift_registerC_0/COL_SEL[34] shift_registerC_0/COL_SEL[35]
+ shift_registerC_0/COL_SEL[36] shift_registerC_0/COL_SEL[37] shift_registerC_0/COL_SEL[38]
+ shift_registerC_0/COL_SEL[39] shift_registerC_0/COL_SEL[40] shift_registerC_0/COL_SEL[41]
+ shift_registerC_0/COL_SEL[42] shift_registerC_0/COL_SEL[43] shift_registerC_0/COL_SEL[44]
+ shift_registerC_0/COL_SEL[45] shift_registerC_0/COL_SEL[46] shift_registerC_0/COL_SEL[47]
+ shift_registerC_0/COL_SEL[48] shift_registerC_0/COL_SEL[49] shift_registerC_0/COL_SEL[50]
+ shift_registerC_0/COL_SEL[51] shift_registerC_0/COL_SEL[52] shift_registerC_0/COL_SEL[53]
+ shift_registerC_0/COL_SEL[54] shift_registerC_0/COL_SEL[55] shift_registerC_0/COL_SEL[56]
+ shift_registerC_0/COL_SEL[57] shift_registerC_0/COL_SEL[58] shift_registerC_0/COL_SEL[59]
+ shift_registerC_0/COL_SEL[60] shift_registerC_0/COL_SEL[61] shift_registerC_0/COL_SEL[62]
+ shift_registerC_0/COL_SEL[63] shift_registerC_0/COL_SEL[64] shift_registerC_0/COL_SEL[65]
+ shift_registerC_0/COL_SEL[66] shift_registerC_0/COL_SEL[67] shift_registerC_0/COL_SEL[68]
+ shift_registerC_0/COL_SEL[69] shift_registerC_0/COL_SEL[70] shift_registerC_0/COL_SEL[71]
+ shift_registerC_0/COL_SEL[72] shift_registerC_0/COL_SEL[73] shift_registerC_0/COL_SEL[74]
+ shift_registerC_0/COL_SEL[75] shift_registerC_0/COL_SEL[76] shift_registerC_0/COL_SEL[77]
+ shift_registerC_0/COL_SEL[78] shift_registerC_0/COL_SEL[79] shift_registerC_0/COL_SEL[80]
+ shift_registerC_0/COL_SEL[81] shift_registerC_0/COL_SEL[82] shift_registerC_0/COL_SEL[83]
+ shift_registerC_0/COL_SEL[84] shift_registerC_0/COL_SEL[85] shift_registerC_0/COL_SEL[86]
+ shift_registerC_0/COL_SEL[87] shift_registerC_0/COL_SEL[88] shift_registerC_0/COL_SEL[89]
+ shift_registerC_0/COL_SEL[90] shift_registerC_0/COL_SEL[91] shift_registerC_0/COL_SEL[92]
+ shift_registerC_0/COL_SEL[93] shift_registerC_0/COL_SEL[94] shift_registerC_0/COL_SEL[95]
+ shift_registerC_0/COL_SEL[96] shift_registerC_0/COL_SEL[97] shift_registerC_0/COL_SEL[98]
+ ARRAY_OUT shift_registerC_0/COL_SEL[99] SF_IB GND pixel_array100x100_fill
.ends

.subckt sky130_fd_pr__pfet_01v8_YT7TV5 a_n505_21# a_n387_21# a_384_118# w_n1642_n937#
+ a_n623_21# a_620_118# a_n387_n815# a_n1150_118# a_n33_n815# a_n741_21# a_321_n815#
+ a_n560_n718# a_675_n815# a_1092_n718# a_n1331_n815# a_n1449_21# a_n914_n718# a_1446_n718#
+ a_1029_n815# a_n151_21# a_n560_118# a_1092_118# a_n269_n815# a_620_n718# a_1328_118#
+ a_30_118# a_203_n815# a_974_n718# a_n442_n718# a_557_n815# a_n796_n718# a_439_21#
+ a_n1213_n815# a_n1213_21# a_n1095_21# a_557_21# a_1328_n718# a_n1331_21# a_n206_118#
+ a_675_21# a_738_118# a_911_21# a_n1268_118# a_793_21# a_n1504_118# a_502_n718# a_n1095_n815#
+ a_856_n718# a_85_n815# a_n324_n718# a_439_n815# a_203_21# a_n678_n718# a_148_118#
+ a_n1449_n815# a_321_21# a_n678_118# a_n33_21# a_n914_118# a_1446_118# a_384_n718#
+ a_1029_21# a_n741_n815# a_30_n718# a_1147_21# a_738_n718# a_n206_n718# a_n324_118#
+ a_1265_21# a_n1150_n718# a_856_118# a_1383_n815# a_1383_21# a_n1386_118# a_n1504_n718#
+ a_266_n718# a_n88_118# a_266_118# a_n623_n815# a_n977_n815# a_502_118# a_n796_118#
+ a_n88_n718# a_n1032_118# a_911_n815# a_n1032_n718# a_1265_n815# a_n1386_n718# a_n151_n815#
+ a_n859_21# a_148_n718# a_n442_118# a_974_118# a_n505_n815# a_n977_21# a_1210_118#
+ a_793_n815# a_n859_n815# a_85_21# a_1210_n718# a_n269_21# a_1147_n815# a_n1268_n718#
X0 a_1446_118# a_1383_21# a_1328_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X1 a_n1032_n718# a_n1095_n815# a_n1150_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_n796_118# a_n859_21# a_n914_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_384_118# a_321_21# a_266_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_384_n718# a_321_n815# a_266_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n88_n718# a_n151_n815# a_n206_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_1328_118# a_1265_21# a_1210_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_n1150_n718# a_n1213_n815# a_n1268_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_n678_118# a_n741_21# a_n796_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_1210_n718# a_1147_n815# a_1092_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_266_118# a_203_21# a_148_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_30_n718# a_n33_n815# a_n88_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_1210_118# a_1147_21# a_1092_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n914_n718# a_n977_n815# a_n1032_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_n560_n718# a_n623_n815# a_n678_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_1446_n718# a_1383_n815# a_1328_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X16 a_n560_118# a_n623_21# a_n678_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_266_n718# a_203_n815# a_148_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_620_n718# a_557_n815# a_502_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_n1386_118# a_n1449_21# a_n1504_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X20 a_n324_118# a_n387_21# a_n442_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_856_118# a_793_21# a_738_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_1092_118# a_1029_21# a_974_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_n324_n718# a_n387_n815# a_n442_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_n442_118# a_n505_21# a_n560_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_148_118# a_85_21# a_30_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_n1386_n718# a_n1449_n815# a_n1504_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X27 a_856_n718# a_793_n815# a_738_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_974_118# a_911_21# a_856_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_1092_n718# a_1029_n815# a_974_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X30 a_n1268_118# a_n1331_21# a_n1386_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X31 a_n206_118# a_n269_21# a_n324_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X32 a_738_118# a_675_21# a_620_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X33 a_n796_n718# a_n859_n815# a_n914_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X34 a_n1032_118# a_n1095_21# a_n1150_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X35 a_148_n718# a_85_n815# a_30_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X36 a_1328_n718# a_1265_n815# a_1210_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X37 a_n88_118# a_n151_21# a_n206_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X38 a_30_118# a_n33_21# a_n88_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X39 a_620_118# a_557_21# a_502_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X40 a_502_n718# a_439_n815# a_384_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X41 a_n1150_118# a_n1213_21# a_n1268_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X42 a_n206_n718# a_n269_n815# a_n324_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X43 a_738_n718# a_675_n815# a_620_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X44 a_n1268_n718# a_n1331_n815# a_n1386_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X45 a_n914_118# a_n977_21# a_n1032_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X46 a_n442_n718# a_n505_n815# a_n560_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X47 a_502_118# a_439_21# a_384_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X48 a_974_n718# a_911_n815# a_856_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X49 a_n678_n718# a_n741_n815# a_n796_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_8HUREQ a_384_n709# a_557_n797# a_203_n797# a_n387_21#
+ a_n505_21# a_30_n709# a_n623_21# a_738_n709# a_n206_n709# a_n741_21# a_n324_109#
+ a_856_109# a_85_n797# a_n151_21# a_266_n709# a_439_n797# a_n88_109# a_266_109# a_n88_n709#
+ a_502_109# a_n796_109# a_439_21# a_n741_n797# a_557_21# a_148_n709# a_675_21# a_n442_109#
+ a_793_21# a_203_21# a_n623_n797# a_321_21# a_620_109# a_384_109# a_n33_21# a_n560_n709#
+ a_n151_n797# a_n914_n709# a_n1016_n883# a_793_n797# a_n505_n797# a_n859_n797# a_n560_109#
+ a_620_n709# a_n442_n709# a_30_109# a_n796_n709# a_n387_n797# a_321_n797# a_n33_n797#
+ a_n206_109# a_675_n797# a_738_109# a_502_n709# a_n859_21# a_856_n709# a_n324_n709#
+ a_n678_n709# a_148_109# a_85_21# a_n269_n797# a_n678_109# a_n914_109# a_n269_21#
X0 a_n678_109# a_n741_21# a_n796_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_266_109# a_203_21# a_148_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_30_n709# a_n33_n797# a_n88_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_n560_n709# a_n623_n797# a_n678_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_n560_109# a_n623_21# a_n678_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n324_109# a_n387_21# a_n442_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_266_n709# a_203_n797# a_148_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_620_n709# a_557_n797# a_502_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_856_109# a_793_21# a_738_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X9 a_n324_n709# a_n387_n797# a_n442_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_n442_109# a_n505_21# a_n560_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_148_109# a_85_21# a_30_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_856_n709# a_793_n797# a_738_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n206_109# a_n269_21# a_n324_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_738_109# a_675_21# a_620_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_n796_n709# a_n859_n797# a_n914_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X16 a_148_n709# a_85_n797# a_30_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_620_109# a_557_21# a_502_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_n88_109# a_n151_21# a_n206_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_30_109# a_n33_21# a_n88_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X20 a_502_n709# a_439_n797# a_384_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_n206_n709# a_n269_n797# a_n324_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_738_n709# a_675_n797# a_620_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_n442_n709# a_n505_n797# a_n560_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_502_109# a_439_21# a_384_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_n678_n709# a_n741_n797# a_n796_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_n796_109# a_n859_21# a_n914_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X27 a_384_109# a_321_21# a_266_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_384_n709# a_321_n797# a_266_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_n88_n709# a_n151_n797# a_n206_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_BLS9H9 m3_n1941_n1600# c1_n1841_n1500#
X0 c1_n1841_n1500# m3_n1941_n1600# sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
.ends

.subckt sky130_fd_pr__pfet_01v8_YC9MKB a_856_n300# a_n324_n300# a_n505_n397# a_n678_n300#
+ a_793_n397# a_n859_n397# a_384_n300# a_n387_n397# a_30_n300# a_321_n397# a_n33_n397#
+ a_738_n300# a_n206_n300# a_675_n397# a_266_n300# a_n269_n397# a_n88_n300# a_203_n397#
+ a_557_n397# a_148_n300# a_439_n397# a_85_n397# w_n1052_n519# a_n560_n300# a_n741_n397#
+ a_n914_n300# a_620_n300# a_n442_n300# a_n796_n300# a_n623_n397# a_n151_n397# a_502_n300#
X0 a_n560_n300# a_n623_n397# a_n678_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_30_n300# a_n33_n397# a_n88_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_266_n300# a_203_n397# a_148_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_620_n300# a_557_n397# a_502_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_n324_n300# a_n387_n397# a_n442_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_856_n300# a_793_n397# a_738_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X6 a_n796_n300# a_n859_n397# a_n914_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X7 a_148_n300# a_85_n397# a_30_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_502_n300# a_439_n397# a_384_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_n206_n300# a_n269_n397# a_n324_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_738_n300# a_675_n397# a_620_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_n442_n300# a_n505_n397# a_n560_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_n678_n300# a_n741_n397# a_n796_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_384_n300# a_321_n397# a_266_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_n88_n300# a_n151_n397# a_n206_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_GQFJAV a_15_n75# a_n69_97# a_n175_n249# a_n73_n75#
X0 a_15_n75# a_n69_97# a_n73_n75# a_n175_n249# sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_YCMRKB a_n1390_n815# a_89_n718# a_1678_21# a_915_118#
+ a_1151_n718# a_1914_21# a_n2216_21# a_734_n815# a_n2153_n718# a_380_21# a_n2098_21#
+ a_2032_n815# a_n973_n718# a_n1445_118# a_1796_21# a_1977_118# a_n92_21# a_2386_n815#
+ a_n1744_n815# a_1088_n815# a_n2334_21# w_n3117_n937# a_2803_n718# a_1206_21# a_1505_n718#
+ a_n2507_n718# a_n1209_n718# a_1088_21# a_1859_n718# a_2213_118# a_n2452_21# a_325_118#
+ a_1324_21# a_262_n815# a_n855_118# a_n2743_118# a_n2570_21# a_n328_n815# a_1387_118#
+ a_1442_21# a_1623_118# a_n2570_n815# a_n1272_n815# a_n501_n718# a_1033_n718# a_2331_n718#
+ a_1560_21# a_616_n815# a_n2035_n718# a_89_118# a_n855_n718# a_2685_n718# a_1387_n718#
+ a_2268_n815# a_n2389_n718# a_n2924_n815# a_n1626_n815# a_2685_118# a_n265_118# a_n2153_118#
+ a_797_118# a_n501_118# a_2921_118# a_1033_118# a_2858_21# a_561_n718# a_144_n815#
+ a_n1563_118# a_n383_n718# a_498_n815# a_n2452_n815# a_n1154_n815# a_915_n718# a_2095_118#
+ a_2213_n718# a_2268_21# a_n918_21# a_2331_118# a_n737_n718# a_2567_n718# a_1269_n718#
+ a_443_118# a_n2806_n815# a_2504_21# a_n1508_n815# a_n1681_n718# a_2386_21# a_26_21#
+ a_1560_n815# a_n973_118# a_n2861_118# a_2622_21# a_1741_118# a_1914_n815# a_443_n718#
+ a_n328_21# a_2740_21# a_797_n718# a_n1209_118# a_n800_n815# a_n265_n718# a_2095_n718#
+ a_n446_21# a_n2334_n815# a_n1036_n815# a_n383_118# a_n2271_118# a_n2688_n815# a_2032_21#
+ a_26_n815# a_1151_118# a_n564_21# a_n619_n718# a_2449_n718# a_2150_21# a_n800_21#
+ a_2740_n815# a_n2861_n718# a_n1563_n718# a_1442_n815# a_n619_118# a_n1681_118# a_n682_21#
+ a_n2507_118# a_1796_n815# a_n1508_21# a_n682_n815# a_n1917_n718# a_325_n718# a_n1626_21#
+ a_679_n718# a_n1917_118# a_n210_21# a_n147_n718# a_561_118# a_n2216_n815# a_970_n815#
+ a_n1744_21# a_n1091_n718# a_n1091_118# a_2449_118# a_n1980_n815# a_n1862_21# a_1741_n718#
+ a_n2979_118# a_n1036_21# a_2622_n815# a_n2743_n718# a_n1445_n718# a_1324_n815# a_1859_118#
+ a_n1327_118# a_n1980_21# a_1678_n815# a_n1799_n718# a_n1154_21# a_n210_n815# a_n564_n815#
+ a_207_n718# a_616_21# a_n2098_n815# a_n1272_21# a_n29_118# a_498_21# a_207_118#
+ a_n2389_118# a_734_21# a_852_n815# a_n2271_n718# a_n1390_21# a_n918_n815# a_2150_n815#
+ a_n737_118# a_n2625_118# a_n29_n718# a_1269_118# a_n1862_n815# a_1505_118# a_852_21#
+ a_2921_n718# a_1623_n718# a_n1799_118# a_2504_n815# a_n2625_n718# a_n1327_n718#
+ a_1206_n815# a_1977_n718# a_970_21# a_n2806_21# a_n2979_n718# a_n2688_21# a_2858_n815#
+ a_144_21# a_n92_n815# a_380_n815# a_n147_118# a_n2035_118# a_n2924_21# a_n446_n815#
+ a_2567_118# a_2803_118# a_679_118# a_262_21#
X0 a_561_n718# a_498_n815# a_443_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_n383_118# a_n446_21# a_n501_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_n265_n718# a_n328_n815# a_n383_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_n1445_118# a_n1508_21# a_n1563_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_915_118# a_852_21# a_797_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n2625_n718# a_n2688_n815# a_n2743_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_1151_n718# a_1088_n815# a_1033_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_n2153_118# a_n2216_21# a_n2271_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_797_n718# a_734_n815# a_679_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_2803_118# a_2740_21# a_2685_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_2331_n718# a_2268_n815# a_2213_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_n29_118# a_n92_21# a_n147_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_n1681_n718# a_n1744_n815# a_n1799_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n1209_118# a_n1272_21# a_n1327_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_1859_118# a_1796_21# a_1741_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_n2861_n718# a_n2924_n815# a_n2979_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X16 a_n265_118# a_n328_21# a_n383_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_n1917_n718# a_n1980_n815# a_n2035_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_n2035_n718# a_n2098_n815# a_n2153_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_797_118# a_734_21# a_679_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X20 a_1977_118# a_1914_21# a_1859_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_1269_n718# a_1206_n815# a_1151_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_1623_n718# a_1560_n815# a_1505_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_207_n718# a_144_n815# a_89_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_89_n718# a_26_n815# a_n29_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_n1091_118# a_n1154_21# a_n1209_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_2685_118# a_2622_21# a_2567_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X27 a_1741_118# a_1678_21# a_1623_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_2803_n718# a_2740_n815# a_2685_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_n1091_n718# a_n1154_n815# a_n1209_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X30 a_89_118# a_26_21# a_n29_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X31 a_n2271_n718# a_n2334_n815# a_n2389_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X32 a_1859_n718# a_1796_n815# a_1741_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X33 a_2449_118# a_2386_21# a_2331_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X34 a_n1327_n718# a_n1390_n815# a_n1445_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X35 a_n147_118# a_n210_21# a_n265_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X36 a_n147_n718# a_n210_n815# a_n265_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X37 a_n2861_118# a_n2924_21# a_n2979_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X38 a_n501_n718# a_n564_n815# a_n619_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X39 a_n2507_n718# a_n2570_n815# a_n2625_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X40 a_679_118# a_616_21# a_561_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X41 a_443_118# a_380_21# a_325_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X42 a_n973_118# a_n1036_21# a_n1091_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X43 a_n1917_118# a_n1980_21# a_n2035_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X44 a_679_n718# a_616_n815# a_561_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X45 a_1623_118# a_1560_21# a_1505_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X46 a_2213_n718# a_2150_n815# a_2095_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X47 a_2567_118# a_2504_21# a_2449_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X48 a_1033_n718# a_970_n815# a_915_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X49 a_n2625_118# a_n2688_21# a_n2743_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X50 a_n1563_n718# a_n1626_n815# a_n1681_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X51 a_n737_n718# a_n800_n815# a_n855_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X52 a_2331_118# a_2268_21# a_2213_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X53 a_n2743_n718# a_n2806_n815# a_n2861_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X54 a_2449_n718# a_2386_n815# a_2331_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X55 a_561_118# a_498_21# a_443_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X56 a_n1799_n718# a_n1862_n815# a_n1917_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X57 a_n2743_118# a_n2806_21# a_n2861_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X58 a_n737_118# a_n800_21# a_n855_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X59 a_1505_n718# a_1442_n815# a_1387_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X60 a_n1799_118# a_n1862_21# a_n1917_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X61 a_325_118# a_262_21# a_207_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X62 a_443_n718# a_380_n815# a_325_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X63 a_1505_118# a_1442_21# a_1387_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X64 a_2685_n718# a_2622_n815# a_2567_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X65 a_n973_n718# a_n1036_n815# a_n1091_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X66 a_n2507_118# a_n2570_21# a_n2625_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X67 a_n2153_n718# a_n2216_n815# a_n2271_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X68 a_2213_118# a_2150_21# a_2095_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X69 a_n855_118# a_n918_21# a_n973_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X70 a_n1209_n718# a_n1272_n815# a_n1327_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X71 a_n383_n718# a_n446_n815# a_n501_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X72 a_n2389_n718# a_n2452_n815# a_n2507_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X73 a_n1681_118# a_n1744_21# a_n1799_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X74 a_n619_118# a_n682_21# a_n737_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X75 a_1977_n718# a_1914_n815# a_1859_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X76 a_207_118# a_144_21# a_89_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X77 a_2095_n718# a_2032_n815# a_1977_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X78 a_1387_118# a_1324_21# a_1269_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X79 a_915_n718# a_852_n815# a_797_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X80 a_n29_n718# a_n92_n815# a_n147_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X81 a_n1445_n718# a_n1508_n815# a_n1563_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X82 a_n619_n718# a_n682_n815# a_n737_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X83 a_n2389_118# a_n2452_21# a_n2507_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X84 a_2095_118# a_2032_21# a_1977_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X85 a_1151_118# a_1088_21# a_1033_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X86 a_n501_118# a_n564_21# a_n619_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X87 a_1033_118# a_970_21# a_915_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X88 a_n1563_118# a_n1626_21# a_n1681_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X89 a_n855_n718# a_n918_n815# a_n973_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X90 a_1387_n718# a_1324_n815# a_1269_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X91 a_n2271_118# a_n2334_21# a_n2389_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X92 a_1741_n718# a_1678_n815# a_1623_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X93 a_325_n718# a_262_n815# a_207_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X94 a_2921_118# a_2858_21# a_2803_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X95 a_1269_118# a_1206_21# a_1151_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X96 a_2567_n718# a_2504_n815# a_2449_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X97 a_2921_n718# a_2858_n815# a_2803_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X98 a_n1327_118# a_n1390_21# a_n1445_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X99 a_n2035_118# a_n2098_21# a_n2153_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_8JUMX6 a_2117_109# a_n399_n1009# a_1879_n1097# a_5225_109#
+ a_3301_109# a_3803_21# a_547_21# a_785_n1009# a_1377_n1009# a_n193_21# a_n2027_109#
+ a_n3301_21# a_n3597_n1097# a_n3211_109# a_n5135_109# a_2767_n1097# a_4189_n1009#
+ a_3893_109# a_4395_21# a_n1673_n1097# a_2265_n1009# a_4691_n1097# a_n103_109# a_637_n1009#
+ a_n4485_n1097# a_4247_21# a_1229_n1009# a_3655_n1097# a_5077_n1009# a_n2561_n1097#
+ a_785_109# a_3655_21# a_399_21# a_n251_n1009# a_1731_n1097# a_n3449_n1097# a_1969_109#
+ a_2619_n1097# a_3153_n1009# a_n1525_n1097# a_n695_109# a_n3153_21# a_2117_n1009#
+ a_n5373_n1097# a_4543_n1097# a_3507_21# a_n2561_21# a_n4929_21# a_n1879_109# a_n4337_n1097#
+ a_5077_109# a_n4987_109# a_2915_21# a_n3005_21# a_3507_n1097# a_4041_n1009# a_3153_109#
+ a_n1583_n1009# a_n103_n1009# a_n2413_n1097# a_4099_21# a_n2413_21# a_3005_n1009#
+ a_n933_n1097# a_5431_n1097# a_n1821_21# a_n5225_n1097# a_n4395_n1009# a_n3063_109#
+ a_1969_n1009# a_399_n1097# a_n3301_n1097# a_n2471_n1009# a_1229_109# a_n3359_n1009#
+ a_n991_n1009# a_4337_109# a_2413_109# a_3359_21# a_3893_n1009# a_5521_109# a_n1435_n1009#
+ a_2767_21# a_n5283_n1009# a_2857_n1009# a_n1139_109# a_n2265_21# a_n4247_n1009#
+ a_n2323_109# a_n4247_109# a_n5431_109# a_2619_21# a_n1673_21# a_n2323_n1009# a_4781_n1009#
+ a_n843_n1009# a_n2117_21# a_3745_n1009# a_n45_n1097# a_n1525_21# a_n5135_n1009#
+ a_1821_n1009# a_251_n1097# a_45_109# a_2709_n1009# a_n193_n1097# a_1081_109# a_n3211_n1009#
+ a_n3507_109# a_n4929_n1097# a_4633_n1009# a_n991_109# a_n5521_21# a_103_n1097# a_4189_109#
+ a_1879_21# a_251_21# a_n4987_n1009# a_2265_109# a_5521_n1009# a_5373_109# a_n1377_21#
+ a_489_n1009# a_103_21# a_n4099_109# a_n2175_109# a_991_n1097# a_n5283_109# a_n45_21#
+ a_n1229_21# a_1583_n1097# a_341_109# a_n3951_n1009# a_n1377_n1097# a_3449_109# a_1525_109#
+ a_n4839_n1009# a_1081_n1009# a_4633_109# a_n933_21# a_n5373_21# a_n251_109# a_4395_n1097#
+ a_n2915_n1009# a_n4781_21# a_n4189_n1097# a_3359_n1097# a_2471_n1097# a_n1435_109#
+ a_n3359_109# a_n5225_21# a_843_n1097# a_n2265_n1097# a_n4543_109# a_1435_n1097#
+ a_n785_n1097# a_3211_21# a_n4633_21# a_5283_n1097# a_n3803_n1009# a_2709_109# a_341_n1009#
+ a_n1229_n1097# a_n5077_n1097# a_4247_n1097# a_n3153_n1097# a_n785_21# a_2323_n1097#
+ a_n2619_109# a_n2117_n1097# a_n1287_n1009# a_n637_n1097# a_n3803_109# a_4987_21#
+ a_n5077_21# a_5135_n1097# a_n637_21# a_n4041_n1097# a_193_109# a_3063_21# a_n4485_21#
+ a_3211_n1097# a_n4099_n1009# a_n3005_n1097# a_1377_109# a_2471_21# a_n3893_21# a_n2175_n1009#
+ a_4485_109# a_2561_109# a_4839_21# a_n695_n1009# a_n1139_n1009# a_45_n1009# a_3597_n1009#
+ a_n4337_21# a_n1969_n1097# a_2323_21# a_1673_n1009# a_n1287_109# a_n3745_21# a_4987_n1097#
+ a_n2471_109# a_n4395_109# a_1731_21# a_n5681_n1183# a_n3063_n1009# a_n3893_n1097#
+ a_n489_21# a_4485_n1009# a_n2027_n1009# a_3745_109# a_n547_n1009# a_2561_n1009#
+ a_n2857_n1097# a_1821_109# a_3449_n1009# a_933_n1009# a_1525_n1009# a_n4781_n1097#
+ a_3951_n1097# a_4839_n1097# a_5373_n1009# a_n3655_109# a_n5579_109# a_n4189_21#
+ a_n3745_n1097# a_637_109# a_n1731_109# a_2175_21# a_2915_n1097# a_n3597_21# a_4337_n1009#
+ a_n1821_n1097# a_4929_109# a_1583_21# a_n1879_n1009# a_n2709_n1097# a_n547_109#
+ a_2413_n1009# a_2027_21# a_n1081_21# a_n3449_21# a_n4633_n1097# a_3803_n1097# a_5225_n1009#
+ a_n4839_109# a_1435_21# a_n2857_21# a_3005_109# a_n2915_109# a_n2767_n1009# a_3301_n1009#
+ a_n4691_n1009# a_n5521_n1097# a_n2709_21# a_n5579_n1009# a_695_n1097# a_1287_n1097#
+ a_3597_109# a_1673_109# a_5431_21# a_n3655_n1009# a_193_n1009# a_4781_109# a_4099_n1097#
+ a_n2619_n1009# a_n1731_n1009# a_1287_21# a_991_21# a_2175_n1097# a_489_109# a_n1583_109#
+ a_n1081_n1097# a_n4691_109# a_n4543_n1009# a_547_n1097# a_1139_n1097# a_n489_n1097#
+ a_2857_109# a_n399_109# a_1139_21# a_843_21# a_n3507_n1009# a_3063_n1097# a_4929_n1009#
+ a_5283_21# a_n1969_21# a_n5431_n1009# a_n2767_109# a_4691_21# a_2027_n1097# a_n341_21#
+ a_4041_109# a_933_109# a_n3951_109# a_5135_21# a_n843_109# a_4543_21# a_695_21#
+ a_3951_21# a_n4041_21# a_n341_n1097#
X0 a_n4099_109# a_n4189_21# a_n4247_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X1 a_489_n1009# a_399_n1097# a_341_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X2 a_n843_n1009# a_n933_n1097# a_n991_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X3 a_n1731_n1009# a_n1821_n1097# a_n1879_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X4 a_3597_109# a_3507_21# a_3449_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X5 a_n1287_109# a_n1377_21# a_n1435_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X6 a_4633_109# a_4543_21# a_4485_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X7 a_4485_n1009# a_4395_n1097# a_4337_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X8 a_489_109# a_399_21# a_341_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X9 a_2709_109# a_2619_21# a_2561_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X10 a_1821_109# a_1731_21# a_1673_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X11 a_n2027_n1009# a_n2117_n1097# a_n2175_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X12 a_n547_n1009# a_n637_n1097# a_n695_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X13 a_n1435_n1009# a_n1525_n1097# a_n1583_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X14 a_3745_109# a_3655_21# a_3597_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X15 a_4781_109# a_4691_21# a_4633_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X16 a_4189_n1009# a_4099_n1097# a_4041_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X17 a_2857_109# a_2767_21# a_2709_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X18 a_n4839_109# a_n4929_21# a_n4987_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X19 a_5077_n1009# a_4987_n1097# a_4929_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X20 a_n1139_n1009# a_n1229_n1097# a_n1287_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X21 a_1969_109# a_1879_21# a_1821_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X22 a_n2619_n1009# a_n2709_n1097# a_n2767_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X23 a_193_n1009# a_103_n1097# a_45_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X24 a_n3951_n1009# a_n4041_n1097# a_n4099_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X25 a_n5431_n1009# a_n5521_n1097# a_n5579_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.45
X26 a_n547_109# a_n637_21# a_n695_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X27 a_45_109# a_n45_21# a_n103_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X28 a_2117_109# a_2027_21# a_1969_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X29 a_3153_109# a_3063_21# a_3005_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X30 a_n3211_109# a_n3301_21# a_n3359_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X31 a_45_n1009# a_n45_n1097# a_n103_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X32 a_n5135_n1009# a_n5225_n1097# a_n5283_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X33 a_n103_n1009# a_n193_n1097# a_n251_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X34 a_n991_n1009# a_n1081_n1097# a_n1139_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X35 a_n3063_n1009# a_n3153_n1097# a_n3211_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X36 a_n5135_109# a_n5225_21# a_n5283_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X37 a_1229_109# a_1139_21# a_1081_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X38 a_n2471_n1009# a_n2561_n1097# a_n2619_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X39 a_n4543_n1009# a_n4633_n1097# a_n4691_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X40 a_n695_109# a_n785_21# a_n843_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X41 a_3301_n1009# a_3211_n1097# a_3153_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X42 a_2265_109# a_2175_21# a_2117_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X43 a_n2323_109# a_n2413_21# a_n2471_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X44 a_4189_109# a_4099_21# a_4041_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X45 a_n4247_109# a_n4337_21# a_n4395_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X46 a_n5283_109# a_n5373_21# a_n5431_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X47 a_1377_109# a_1287_21# a_1229_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X48 a_n4247_n1009# a_n4337_n1097# a_n4395_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X49 a_n1435_109# a_n1525_21# a_n1583_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X50 a_n2175_n1009# a_n2265_n1097# a_n2323_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X51 a_n3359_109# a_n3449_21# a_n3507_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X52 a_n3655_n1009# a_n3745_n1097# a_n3803_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X53 a_n2471_109# a_n2561_21# a_n2619_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X54 a_n695_n1009# a_n785_n1097# a_n843_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X55 a_n1583_n1009# a_n1673_n1097# a_n1731_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X56 a_637_109# a_547_21# a_489_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X57 a_2413_n1009# a_2323_n1097# a_2265_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X58 a_n4395_109# a_n4485_21# a_n4543_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X59 a_3893_n1009# a_3803_n1097# a_3745_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X60 a_1821_n1009# a_1731_n1097# a_1673_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X61 a_3893_109# a_3803_21# a_3745_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X62 a_n1583_109# a_n1673_21# a_n1731_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X63 a_n3507_109# a_n3597_21# a_n3655_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X64 a_785_109# a_695_21# a_637_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X65 a_n3359_n1009# a_n3449_n1097# a_n3507_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X66 a_3005_109# a_2915_21# a_2857_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X67 a_n399_n1009# a_n489_n1097# a_n547_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X68 a_n1287_n1009# a_n1377_n1097# a_n1435_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X69 a_n4839_n1009# a_n4929_n1097# a_n4987_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X70 a_2117_n1009# a_2027_n1097# a_1969_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X71 a_341_n1009# a_251_n1097# a_193_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X72 a_n2767_n1009# a_n2857_n1097# a_n2915_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X73 a_4929_109# a_4839_21# a_4781_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X74 a_4041_109# a_3951_21# a_3893_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X75 a_n103_109# a_n193_21# a_n251_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X76 a_3597_n1009# a_3507_n1097# a_3449_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X77 a_1525_n1009# a_1435_n1097# a_1377_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X78 a_3005_n1009# a_2915_n1097# a_2857_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X79 a_5077_109# a_4987_21# a_4929_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X80 a_1229_n1009# a_1139_n1097# a_1081_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X81 a_n1879_n1009# a_n1969_n1097# a_n2027_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X82 a_2709_n1009# a_2619_n1097# a_2561_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X83 a_n5283_n1009# a_n5373_n1097# a_n5431_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X84 a_933_n1009# a_843_n1097# a_785_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X85 a_n4691_n1009# a_n4781_n1097# a_n4839_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X86 a_5521_n1009# a_5431_n1097# a_5373_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.45
X87 a_3301_109# a_3211_21# a_3153_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X88 a_5225_109# a_5135_21# a_5077_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X89 a_n991_109# a_n1081_21# a_n1139_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X90 a_n843_109# a_n933_21# a_n991_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X91 a_2413_109# a_2323_21# a_2265_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X92 a_n4987_n1009# a_n5077_n1097# a_n5135_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X93 a_637_n1009# a_547_n1097# a_489_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X94 a_4337_109# a_4247_21# a_4189_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X95 a_n4395_n1009# a_n4485_n1097# a_n4543_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X96 a_5225_n1009# a_5135_n1097# a_5077_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X97 a_3153_n1009# a_3063_n1097# a_3005_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X98 a_n3803_n1009# a_n3893_n1097# a_n3951_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X99 a_5373_109# a_5283_21# a_5225_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X100 a_n5431_109# a_n5521_21# a_n5579_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.45
X101 a_1525_109# a_1435_21# a_1377_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X102 a_4633_n1009# a_4543_n1097# a_4485_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X103 a_2561_n1009# a_2471_n1097# a_2413_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X104 a_4041_n1009# a_3951_n1097# a_3893_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X105 a_3449_109# a_3359_21# a_3301_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X106 a_2561_109# a_2471_21# a_2413_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X107 a_4485_109# a_4395_21# a_4337_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X108 a_n4543_109# a_n4633_21# a_n4691_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X109 a_n4099_n1009# a_n4189_n1097# a_n4247_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X110 a_1673_109# a_1583_21# a_1525_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X111 a_n3507_n1009# a_n3597_n1097# a_n3655_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X112 a_n2619_109# a_n2709_21# a_n2767_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X113 a_n1731_109# a_n1821_21# a_n1879_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X114 a_4337_n1009# a_4247_n1097# a_4189_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X115 a_2265_n1009# a_2175_n1097# a_2117_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X116 a_n3655_109# a_n3745_21# a_n3803_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X117 a_3745_n1009# a_3655_n1097# a_3597_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X118 a_933_109# a_843_21# a_785_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X119 a_1673_n1009# a_1583_n1097# a_1525_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X120 a_n4691_109# a_n4781_21# a_n4839_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X121 a_n251_109# a_n341_21# a_n399_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X122 a_n2767_109# a_n2857_21# a_n2915_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X123 a_n3803_109# a_n3893_21# a_n3951_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X124 a_1081_109# a_991_21# a_933_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X125 a_3449_n1009# a_3359_n1097# a_3301_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X126 a_4929_n1009# a_4839_n1097# a_4781_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X127 a_1377_n1009# a_1287_n1097# a_1229_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X128 a_n1879_109# a_n1969_21# a_n2027_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X129 a_2857_n1009# a_2767_n1097# a_2709_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X130 a_1081_n1009# a_991_n1097# a_933_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X131 a_n2915_109# a_n3005_21# a_n3063_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X132 a_193_109# a_103_21# a_45_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X133 a_n3951_109# a_n4041_21# a_n4099_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X134 a_n399_109# a_n489_21# a_n547_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X135 a_n3211_n1009# a_n3301_n1097# a_n3359_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X136 a_n251_n1009# a_n341_n1097# a_n399_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X137 a_n2027_109# a_n2117_21# a_n2175_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X138 a_785_n1009# a_695_n1097# a_637_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X139 a_1969_n1009# a_1879_n1097# a_1821_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X140 a_n3063_109# a_n3153_21# a_n3211_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X141 a_5373_n1009# a_5283_n1097# a_5225_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X142 a_341_109# a_251_21# a_193_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X143 a_n4987_109# a_n5077_21# a_n5135_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X144 a_4781_n1009# a_4691_n1097# a_4633_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X145 a_n1139_109# a_n1229_21# a_n1287_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X146 a_n2915_n1009# a_n3005_n1097# a_n3063_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X147 a_n2175_109# a_n2265_21# a_n2323_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X148 a_5521_109# a_5431_21# a_5373_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.45
X149 a_n2323_n1009# a_n2413_n1097# a_n2471_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
.ends

.subckt opamp_v1 iref vin_n vin_p vout vdd vss a_4019_n9933#
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[0] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[1] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[2] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__nfet_01v8_8HUREQ_0 vbn vbn vbn vbn vbn vss vbn vss vss vbn vbn vbn
+ vbn vbn vss vbn vbn vss vbn vss vbn vbn vbn vbn vbn vbn vss vbn vbn vbn vbn vbn
+ vbn vbn vbn vbn vss vss vbn vbn vbn vbn vbn vss vss vbn vbn vbn vbn vss vbn vss
+ vss vbn vbn vbn vss vbn vbn vbn vss vss vbn sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__nfet_01v8_8HUREQ_1 voe1 vbn vbn vbn vbn vss vbn vss vss vbn voe1 voe1
+ vbn vbn vss vbn voe1 vss voe1 vss voe1 vbn vbn vbn voe1 vbn vss vbn vbn vbn vbn
+ voe1 voe1 vbn voe1 vbn vss vss vbn vbn vbn voe1 voe1 vss vss voe1 vbn vbn vbn vss
+ vbn vss vss vbn voe1 voe1 vss voe1 vbn vbn vss vss vbn sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_0 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_1 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_2 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_1 w_4660_n6791# w_4660_n6791# iref vdd iref iref w_4660_n6791#
+ iref vdd iref iref vdd vdd iref vdd iref w_4660_n6791# iref iref w_4660_n6791# iref
+ iref vdd w_4660_n6791# iref vdd w_4660_n6791# vdd w_4660_n6791# iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__pfet_01v8_YC9MKB_0 iref iref iref vdd iref iref iref iref vdd iref
+ iref vdd vdd iref vdd iref iref iref iref iref iref iref vdd iref iref vdd iref
+ vdd iref iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_3 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_2 w_4660_n6791# w_4660_n6791# iref vdd iref iref w_4660_n6791#
+ iref vdd iref iref vdd vdd iref vdd iref w_4660_n6791# iref iref w_4660_n6791# iref
+ iref vdd w_4660_n6791# iref vdd w_4660_n6791# vdd w_4660_n6791# iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_4 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_5 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__nfet_01v8_GQFJAV_0 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_1 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_2 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_3 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_4 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_5 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__pfet_01v8_YCMRKB_0 vin_p w_4660_n6791# vin_p voe1 voe1 vin_p vin_p
+ vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791# vin_p vin_p vin_p vin_p
+ vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 w_4660_n6791#
+ vin_p w_4660_n6791# vin_p vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p voe1 vin_p
+ voe1 vin_p vin_p voe1 w_4660_n6791# voe1 vin_p vin_p w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 vin_p vin_p w_4660_n6791# voe1 voe1
+ w_4660_n6791# voe1 w_4660_n6791# w_4660_n6791# vin_p w_4660_n6791# vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 voe1 w_4660_n6791# vin_p vin_p voe1 voe1 voe1
+ w_4660_n6791# voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791#
+ vin_p voe1 vin_p vin_p w_4660_n6791# voe1 vin_p voe1 voe1 vin_p vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p voe1 voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p
+ vin_p vin_p w_4660_n6791# w_4660_n6791# w_4660_n6791# vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p w_4660_n6791# voe1 vin_p voe1 w_4660_n6791# vin_p vin_p
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 vin_p voe1 voe1 vin_p
+ vin_p w_4660_n6791# vin_p vin_p vin_p voe1 voe1 voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p w_4660_n6791# voe1 w_4660_n6791# vin_p voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p vin_p w_4660_n6791# vin_p vin_p vin_p vin_p vin_p w_4660_n6791# w_4660_n6791#
+ vin_p vin_p voe1 voe1 voe1 vin_p sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_1 vin_n w_4660_n6791# vin_n vbn vbn vin_n vin_n vin_n
+ vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vin_n vin_n vin_n vin_n
+ w_4660_n6791# vbn vin_n w_4660_n6791# w_4660_n6791# vbn vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vin_n
+ vbn vin_n vin_n vbn w_4660_n6791# vbn vin_n vin_n w_4660_n6791# w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# vbn vin_n vbn vin_n vin_n w_4660_n6791# vbn vbn w_4660_n6791# vbn
+ w_4660_n6791# w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vbn w_4660_n6791# vin_n vin_n vbn vbn vbn w_4660_n6791# vbn
+ vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vbn vin_n
+ vin_n w_4660_n6791# vbn vin_n vbn vbn vin_n vin_n vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vbn vin_n w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n vbn vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n
+ w_4660_n6791# vbn vin_n vbn w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vin_n vin_n vin_n vbn vin_n vbn vbn vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vbn vbn w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# vbn w_4660_n6791#
+ vin_n vbn w_4660_n6791# vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vbn vbn vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_2 vin_n w_4660_n6791# vin_n vbn vbn vin_n vin_n vin_n
+ vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vin_n vin_n vin_n vin_n
+ w_4660_n6791# vbn vin_n w_4660_n6791# w_4660_n6791# vbn vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vin_n
+ vbn vin_n vin_n vbn w_4660_n6791# vbn vin_n vin_n w_4660_n6791# w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# vbn vin_n vbn vin_n vin_n w_4660_n6791# vbn vbn w_4660_n6791# vbn
+ w_4660_n6791# w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vbn w_4660_n6791# vin_n vin_n vbn vbn vbn w_4660_n6791# vbn
+ vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vbn vin_n
+ vin_n w_4660_n6791# vbn vin_n vbn vbn vin_n vin_n vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vbn vin_n w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n vbn vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n
+ w_4660_n6791# vbn vin_n vbn w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vin_n vin_n vin_n vbn vin_n vbn vbn vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vbn vbn w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# vbn w_4660_n6791#
+ vin_n vbn w_4660_n6791# vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vbn vbn vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__nfet_01v8_8JUMX6_0 vss vout voe1 vout vss voe1 voe1 vout vout voe1
+ vss voe1 voe1 vss vout voe1 vss vss voe1 voe1 vout voe1 vout vss voe1 voe1 vss voe1
+ vss voe1 vout voe1 voe1 vss voe1 voe1 vout voe1 vout voe1 vout voe1 vss voe1 voe1
+ voe1 voe1 voe1 vout voe1 vss vss voe1 voe1 voe1 vout vout vout vout voe1 voe1 voe1
+ vss voe1 voe1 voe1 voe1 vss vout vout voe1 voe1 vout vss vout vout vout vss voe1
+ vss vout vss voe1 vss vout vss voe1 vout vss vout vout voe1 voe1 vss vss vss voe1
+ vout voe1 voe1 vout vss voe1 vss vss voe1 vout vss vss voe1 vout vout voe1 voe1
+ vss voe1 voe1 vss vout vout vss voe1 vout voe1 vss vout voe1 vss voe1 voe1 voe1
+ vss vout voe1 vout vss vout vout vout voe1 voe1 vss voe1 vss voe1 voe1 voe1 voe1
+ vss vout voe1 voe1 voe1 vout voe1 voe1 voe1 voe1 voe1 vss vss vss voe1 voe1 voe1
+ voe1 voe1 voe1 vss voe1 vout voe1 vss voe1 voe1 voe1 voe1 voe1 vout voe1 voe1 voe1
+ vss voe1 vout voe1 voe1 vout vss vout voe1 vout vss vss vss voe1 voe1 voe1 vout
+ vout voe1 voe1 vout vss voe1 vss vout voe1 voe1 vss vss vout vss vout voe1 vss vout
+ vss vss voe1 voe1 voe1 vss vout vss voe1 voe1 vss vss voe1 voe1 voe1 vout voe1 vout
+ voe1 vout voe1 vss vss voe1 voe1 voe1 voe1 voe1 vout vout voe1 voe1 vss vss vout
+ vss vss voe1 voe1 vss voe1 voe1 vss vout voe1 vout vout vss voe1 vss vss voe1 voe1
+ voe1 vout vout voe1 vss vout voe1 voe1 voe1 vout vout voe1 voe1 vss voe1 vout voe1
+ voe1 vout vout voe1 voe1 voe1 vout vss vout voe1 vss voe1 voe1 voe1 voe1 voe1 sky130_fd_pr__nfet_01v8_8JUMX6
Xsky130_fd_pr__pfet_01v8_YCMRKB_3 vin_p w_4660_n6791# vin_p voe1 voe1 vin_p vin_p
+ vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791# vin_p vin_p vin_p vin_p
+ vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 w_4660_n6791#
+ vin_p w_4660_n6791# vin_p vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p voe1 vin_p
+ voe1 vin_p vin_p voe1 w_4660_n6791# voe1 vin_p vin_p w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 vin_p vin_p w_4660_n6791# voe1 voe1
+ w_4660_n6791# voe1 w_4660_n6791# w_4660_n6791# vin_p w_4660_n6791# vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 voe1 w_4660_n6791# vin_p vin_p voe1 voe1 voe1
+ w_4660_n6791# voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791#
+ vin_p voe1 vin_p vin_p w_4660_n6791# voe1 vin_p voe1 voe1 vin_p vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p voe1 voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p
+ vin_p vin_p w_4660_n6791# w_4660_n6791# w_4660_n6791# vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p w_4660_n6791# voe1 vin_p voe1 w_4660_n6791# vin_p vin_p
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 vin_p voe1 voe1 vin_p
+ vin_p w_4660_n6791# vin_p vin_p vin_p voe1 voe1 voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p w_4660_n6791# voe1 w_4660_n6791# vin_p voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p vin_p w_4660_n6791# vin_p vin_p vin_p vin_p vin_p w_4660_n6791# w_4660_n6791#
+ vin_p vin_p voe1 voe1 voe1 vin_p sky130_fd_pr__pfet_01v8_YCMRKB
.ends

.subckt opamp_wrapper AOUT OUT_IB AMP_IB ARRAY_OUT VSS VDD
Xopamp_v1_0 opamp_v1_0/iref AOUT ARRAY_OUT AOUT VDD VSS VSS opamp_v1
X0 ARRAY_OUT OUT_IB VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=31.9 pd=27 as=11.5 ps=22.3 w=10 l=0.15
X1 opamp_v1_0/iref AMP_IB VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=34.4 pd=27.7 as=11.5 ps=22.3 w=10 l=0.15
.ends

.subckt bias VDD NB1 NB2 OUT_IB AMP_IB GND SF_IB
X0 NB1 NB1 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.35 ps=2.7 w=1 l=1.2
X1 NB2 NB2 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.35 pd=2.7 as=0.35 ps=2.7 w=1 l=1.2
X2 AMP_IB AMP_IB GND GND sky130_fd_pr__nfet_01v8_lvt ad=5.6 pd=17.4 as=5.2 ps=17.3 w=8 l=2
X3 OUT_IB OUT_IB GND GND sky130_fd_pr__nfet_01v8_lvt ad=5.6 pd=17.4 as=5.2 ps=17.3 w=8 l=2
X4 SF_IB SF_IB VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0.55 pd=3.1 as=0.45 ps=2.9 w=1 l=1
.ends

.subckt sky130_fd_pr__res_generic_m3_3NNQKJ m3_n50_n107# m3_n50_50#
R0 m3_n50_50# m3_n50_n107# sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xpixel_array_0 io_analog[7] io_analog[8] io_analog[4] vccd1 io_analog[6] io_analog[9]
+ io_in[20] io_in[21] io_in[22] pixel_array_0/PIX0_IN io_analog[10] pixel_array_0/PIX1_IN
+ pixel_array_0/PIX2_IN pixel_array_0/PIX3_IN pixel_array_0/PIX4_IN pixel_array_0/PIX5_IN
+ pixel_array_0/PIX6_IN pixel_array_0/PIX_OUT0 pixel_array_0/PIX7_IN pixel_array_0/PIX_OUT1
+ pixel_array_0/PIX8_IN pixel_array_0/PIX_OUT2 pixel_array_0/ARRAY_OUT io_in[23] io_in[24]
+ io_in[15] vssd1 io_analog[5] pixel_array
Xarray_SR_0 vccd1 io_in[7] io_in[8] io_in[9] io_in[6] io_analog[9] array_SR_0/ARRAY_OUT
+ io_analog[5] io_analog[4] io_analog[7] io_analog[8] io_analog[6] io_in[19] io_analog[10]
+ io_in[16] io_in[18] io_in[17] vssd1 array_SR
Xopamp_wrapper_0 io_analog[0] io_analog[3] io_analog[2] array_SR_0/ARRAY_OUT vssd1
+ vccd1 opamp_wrapper
Xopamp_wrapper_1 io_analog[1] io_analog[3] io_analog[2] pixel_array_0/ARRAY_OUT vssd1
+ vccd1 opamp_wrapper
Xbias_1 vccd1 io_analog[5] io_analog[4] io_analog[3] io_analog[2] vssd1 io_analog[6]
+ bias
Xsky130_fd_pr__res_generic_m3_3NNQKJ_0 vccd1 io_oeb[9] sky130_fd_pr__res_generic_m3_3NNQKJ
Xsky130_fd_pr__res_generic_m3_3NNQKJ_1 io_oeb[15] vccd1 sky130_fd_pr__res_generic_m3_3NNQKJ
R0 io_oeb[21] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R1 vccd1 io_oeb[6] sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R2 vccd1 io_oeb[8] sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R3 io_oeb[19] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R4 io_oeb[17] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R5 io_oeb[24] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R6 vccd1 io_oeb[7] sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R7 io_oeb[23] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R8 io_oeb[16] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R9 io_oeb[20] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R10 io_oeb[22] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
R11 io_oeb[18] vccd1 sky130_fd_pr__res_generic_m3 w=0.5 l=0.5
.ends

