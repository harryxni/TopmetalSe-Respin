magic
tech sky130A
timestamp 1757709129
<< metal1 >>
rect 151254 162266 151354 162269
rect 151254 160679 151354 162166
rect 151963 160679 152123 160682
rect 151254 160519 151963 160679
rect 54 159961 154 160155
rect 151254 160049 151354 160519
rect 151963 160516 152123 160519
rect 51 159861 54 159961
rect 154 159861 157 159961
rect 51 159850 157 159861
rect 54 159725 154 159850
rect 151963 159179 152123 159182
rect 151268 159019 151963 159179
rect 151963 159016 152123 159019
rect 54 158461 154 158655
rect 51 158361 54 158461
rect 154 158361 157 158461
rect 51 158350 157 158361
rect 54 158225 154 158350
rect 151963 157679 152123 157682
rect 151268 157519 151963 157679
rect 151963 157516 152123 157519
rect 54 156961 154 157155
rect 51 156861 54 156961
rect 154 156861 157 156961
rect 51 156850 157 156861
rect 54 156725 154 156850
rect 151963 156179 152123 156182
rect 151268 156019 151963 156179
rect 151963 156016 152123 156019
rect 54 155461 154 155655
rect 51 155361 54 155461
rect 154 155361 157 155461
rect 51 155350 157 155361
rect 54 155225 154 155350
rect 151963 154679 152123 154682
rect 151268 154519 151963 154679
rect 151963 154516 152123 154519
rect 54 153961 154 154155
rect 51 153861 54 153961
rect 154 153861 157 153961
rect 51 153850 157 153861
rect 54 153725 154 153850
rect 151963 153179 152123 153182
rect 151268 153019 151963 153179
rect 151963 153016 152123 153019
rect 54 152461 154 152655
rect 51 152361 54 152461
rect 154 152361 157 152461
rect 51 152350 157 152361
rect 54 152225 154 152350
rect 151963 151679 152123 151682
rect 151268 151519 151963 151679
rect 151963 151516 152123 151519
rect 54 150961 154 151155
rect 51 150861 54 150961
rect 154 150861 157 150961
rect 51 150850 157 150861
rect 54 150725 154 150850
rect 151963 150179 152123 150182
rect 151268 150019 151963 150179
rect 151963 150016 152123 150019
rect 54 149461 154 149655
rect 51 149361 54 149461
rect 154 149361 157 149461
rect 51 149350 157 149361
rect 54 149225 154 149350
rect 151963 148679 152123 148682
rect 151268 148519 151963 148679
rect 151963 148516 152123 148519
rect 54 147961 154 148155
rect 51 147861 54 147961
rect 154 147861 157 147961
rect 51 147850 157 147861
rect 54 147725 154 147850
rect 151963 147179 152123 147182
rect 151268 147019 151963 147179
rect 151963 147016 152123 147019
rect 54 146461 154 146655
rect 51 146361 54 146461
rect 154 146361 157 146461
rect 51 146350 157 146361
rect 54 146225 154 146350
rect 151963 145679 152123 145682
rect 151268 145519 151963 145679
rect 151963 145516 152123 145519
rect 54 144961 154 145155
rect 51 144861 54 144961
rect 154 144861 157 144961
rect 51 144850 157 144861
rect 54 144725 154 144850
rect 151963 144179 152123 144182
rect 151268 144019 151963 144179
rect 151963 144016 152123 144019
rect 54 143461 154 143655
rect 51 143361 54 143461
rect 154 143361 157 143461
rect 51 143350 157 143361
rect 54 143225 154 143350
rect 151963 142679 152123 142682
rect 151268 142519 151963 142679
rect 151963 142516 152123 142519
rect 54 141961 154 142155
rect 51 141861 54 141961
rect 154 141861 157 141961
rect 51 141850 157 141861
rect 54 141725 154 141850
rect 151963 141179 152123 141182
rect 151268 141019 151963 141179
rect 151963 141016 152123 141019
rect 54 140461 154 140655
rect 51 140361 54 140461
rect 154 140361 157 140461
rect 51 140350 157 140361
rect 54 140225 154 140350
rect 151963 139679 152123 139682
rect 151268 139519 151963 139679
rect 151963 139516 152123 139519
rect 54 138961 154 139155
rect 51 138861 54 138961
rect 154 138861 157 138961
rect 51 138850 157 138861
rect 54 138725 154 138850
rect 151963 138179 152123 138182
rect 151268 138019 151963 138179
rect 151963 138016 152123 138019
rect 54 137461 154 137655
rect 51 137361 54 137461
rect 154 137361 157 137461
rect 51 137350 157 137361
rect 54 137225 154 137350
rect 151963 136679 152123 136682
rect 151268 136519 151963 136679
rect 151963 136516 152123 136519
rect 54 135961 154 136155
rect 51 135861 54 135961
rect 154 135861 157 135961
rect 51 135850 157 135861
rect 54 135725 154 135850
rect 151963 135179 152123 135182
rect 151268 135019 151963 135179
rect 151963 135016 152123 135019
rect 54 134461 154 134655
rect 51 134361 54 134461
rect 154 134361 157 134461
rect 51 134350 157 134361
rect 54 134225 154 134350
rect 151963 133679 152123 133682
rect 151268 133519 151963 133679
rect 151963 133516 152123 133519
rect 54 132961 154 133155
rect 51 132861 54 132961
rect 154 132861 157 132961
rect 51 132850 157 132861
rect 54 132725 154 132850
rect 151963 132179 152123 132182
rect 151268 132019 151963 132179
rect 151963 132016 152123 132019
rect 54 131461 154 131655
rect 51 131361 54 131461
rect 154 131361 157 131461
rect 51 131350 157 131361
rect 54 131225 154 131350
rect 151963 130679 152123 130682
rect 151268 130519 151963 130679
rect 151963 130516 152123 130519
rect 54 129961 154 130155
rect 51 129861 54 129961
rect 154 129861 157 129961
rect 51 129850 157 129861
rect 54 129725 154 129850
rect 151963 129179 152123 129182
rect 151268 129019 151963 129179
rect 151963 129016 152123 129019
rect 54 128461 154 128655
rect 51 128361 54 128461
rect 154 128361 157 128461
rect 51 128350 157 128361
rect 54 128225 154 128350
rect 151963 127679 152123 127682
rect 151268 127519 151963 127679
rect 151963 127516 152123 127519
rect 54 126961 154 127155
rect 51 126861 54 126961
rect 154 126861 157 126961
rect 51 126850 157 126861
rect 54 126725 154 126850
rect 151963 126179 152123 126182
rect 151268 126019 151963 126179
rect 151963 126016 152123 126019
rect 54 125461 154 125655
rect 51 125361 54 125461
rect 154 125361 157 125461
rect 51 125350 157 125361
rect 54 125225 154 125350
rect 151963 124679 152123 124682
rect 151268 124519 151963 124679
rect 151963 124516 152123 124519
rect 54 123961 154 124155
rect 51 123861 54 123961
rect 154 123861 157 123961
rect 51 123850 157 123861
rect 54 123725 154 123850
rect 151963 123179 152123 123182
rect 151268 123019 151963 123179
rect 151963 123016 152123 123019
rect 54 122461 154 122655
rect 51 122361 54 122461
rect 154 122361 157 122461
rect 51 122350 157 122361
rect 54 122225 154 122350
rect 151963 121679 152123 121682
rect 151268 121519 151963 121679
rect 151963 121516 152123 121519
rect 54 120961 154 121155
rect 51 120861 54 120961
rect 154 120861 157 120961
rect 51 120850 157 120861
rect 54 120725 154 120850
rect 151963 120179 152123 120182
rect 151268 120019 151963 120179
rect 151963 120016 152123 120019
rect 54 119461 154 119655
rect 51 119361 54 119461
rect 154 119361 157 119461
rect 51 119350 157 119361
rect 54 119225 154 119350
rect 151963 118679 152123 118682
rect 151268 118519 151963 118679
rect 151963 118516 152123 118519
rect 54 117961 154 118155
rect 51 117861 54 117961
rect 154 117861 157 117961
rect 51 117850 157 117861
rect 54 117725 154 117850
rect 151963 117179 152123 117182
rect 151268 117019 151963 117179
rect 151963 117016 152123 117019
rect 54 116461 154 116655
rect 51 116361 54 116461
rect 154 116361 157 116461
rect 51 116350 157 116361
rect 54 116225 154 116350
rect 151963 115679 152123 115682
rect 151268 115519 151963 115679
rect 151963 115516 152123 115519
rect 54 114961 154 115155
rect 51 114861 54 114961
rect 154 114861 157 114961
rect 51 114850 157 114861
rect 54 114725 154 114850
rect 151963 114179 152123 114182
rect 151268 114019 151963 114179
rect 151963 114016 152123 114019
rect 54 113461 154 113655
rect 51 113361 54 113461
rect 154 113361 157 113461
rect 51 113350 157 113361
rect 54 113225 154 113350
rect 151963 112679 152123 112682
rect 151268 112519 151963 112679
rect 151963 112516 152123 112519
rect 54 111961 154 112155
rect 51 111861 54 111961
rect 154 111861 157 111961
rect 51 111850 157 111861
rect 54 111725 154 111850
rect 151963 111179 152123 111182
rect 151268 111019 151963 111179
rect 151963 111016 152123 111019
rect 54 110461 154 110655
rect 51 110361 54 110461
rect 154 110361 157 110461
rect 51 110350 157 110361
rect 54 110225 154 110350
rect 151963 109679 152123 109682
rect 151268 109519 151963 109679
rect 151963 109516 152123 109519
rect 54 108961 154 109155
rect 51 108861 54 108961
rect 154 108861 157 108961
rect 51 108850 157 108861
rect 54 108725 154 108850
rect 151963 108179 152123 108182
rect 151268 108019 151963 108179
rect 151963 108016 152123 108019
rect 54 107461 154 107655
rect 51 107361 54 107461
rect 154 107361 157 107461
rect 51 107350 157 107361
rect 54 107225 154 107350
rect 151963 106679 152123 106682
rect 151268 106519 151963 106679
rect 151963 106516 152123 106519
rect 54 105961 154 106155
rect 51 105861 54 105961
rect 154 105861 157 105961
rect 51 105850 157 105861
rect 54 105725 154 105850
rect 151963 105179 152123 105182
rect 151268 105019 151963 105179
rect 151963 105016 152123 105019
rect 54 104461 154 104655
rect 51 104361 54 104461
rect 154 104361 157 104461
rect 51 104350 157 104361
rect 54 104225 154 104350
rect 151963 103679 152123 103682
rect 151268 103519 151963 103679
rect 151963 103516 152123 103519
rect 54 102961 154 103155
rect 51 102861 54 102961
rect 154 102861 157 102961
rect 51 102850 157 102861
rect 54 102725 154 102850
rect 151963 102179 152123 102182
rect 151268 102019 151963 102179
rect 151963 102016 152123 102019
rect 54 101461 154 101655
rect 51 101361 54 101461
rect 154 101361 157 101461
rect 51 101350 157 101361
rect 54 101225 154 101350
rect 151963 100679 152123 100682
rect 151268 100519 151963 100679
rect 151963 100516 152123 100519
rect 54 99961 154 100155
rect 51 99861 54 99961
rect 154 99861 157 99961
rect 51 99850 157 99861
rect 54 99725 154 99850
rect 151963 99179 152123 99182
rect 151268 99019 151963 99179
rect 151963 99016 152123 99019
rect 54 98461 154 98655
rect 51 98361 54 98461
rect 154 98361 157 98461
rect 51 98350 157 98361
rect 54 98225 154 98350
rect 151963 97679 152123 97682
rect 151268 97519 151963 97679
rect 151963 97516 152123 97519
rect 54 96961 154 97155
rect 51 96861 54 96961
rect 154 96861 157 96961
rect 51 96850 157 96861
rect 54 96725 154 96850
rect 151963 96179 152123 96182
rect 151268 96019 151963 96179
rect 151963 96016 152123 96019
rect 54 95461 154 95655
rect 51 95361 54 95461
rect 154 95361 157 95461
rect 51 95350 157 95361
rect 54 95225 154 95350
rect 151963 94679 152123 94682
rect 151268 94519 151963 94679
rect 151963 94516 152123 94519
rect 54 93961 154 94155
rect 51 93861 54 93961
rect 154 93861 157 93961
rect 51 93850 157 93861
rect 54 93725 154 93850
rect 151963 93179 152123 93182
rect 151268 93019 151963 93179
rect 151963 93016 152123 93019
rect 54 92461 154 92655
rect 51 92361 54 92461
rect 154 92361 157 92461
rect 51 92350 157 92361
rect 54 92225 154 92350
rect 151963 91679 152123 91682
rect 151268 91519 151963 91679
rect 151963 91516 152123 91519
rect 54 90961 154 91155
rect 51 90861 54 90961
rect 154 90861 157 90961
rect 51 90850 157 90861
rect 54 90725 154 90850
rect 151963 90179 152123 90182
rect 151268 90019 151963 90179
rect 151963 90016 152123 90019
rect 54 89461 154 89655
rect 51 89361 54 89461
rect 154 89361 157 89461
rect 51 89350 157 89361
rect 54 89225 154 89350
rect 151963 88679 152123 88682
rect 151268 88519 151963 88679
rect 151963 88516 152123 88519
rect 54 87961 154 88155
rect 51 87861 54 87961
rect 154 87861 157 87961
rect 51 87850 157 87861
rect 54 87725 154 87850
rect 151963 87179 152123 87182
rect 151268 87019 151963 87179
rect 151963 87016 152123 87019
rect 54 86461 154 86655
rect 51 86361 54 86461
rect 154 86361 157 86461
rect 51 86350 157 86361
rect 54 86225 154 86350
rect 151963 85679 152123 85682
rect 151268 85519 151963 85679
rect 151963 85516 152123 85519
rect 54 84961 154 85155
rect 51 84861 54 84961
rect 154 84861 157 84961
rect 51 84850 157 84861
rect 54 84725 154 84850
rect 151963 84179 152123 84182
rect 151268 84019 151963 84179
rect 151963 84016 152123 84019
rect 54 83461 154 83655
rect 51 83361 54 83461
rect 154 83361 157 83461
rect 51 83350 157 83361
rect 54 83225 154 83350
rect 151963 82679 152123 82682
rect 151268 82519 151963 82679
rect 151963 82516 152123 82519
rect 54 81961 154 82155
rect 51 81861 54 81961
rect 154 81861 157 81961
rect 51 81850 157 81861
rect 54 81725 154 81850
rect 151963 81179 152123 81182
rect 151268 81019 151963 81179
rect 151963 81016 152123 81019
rect 54 80461 154 80655
rect 51 80361 54 80461
rect 154 80361 157 80461
rect 51 80350 157 80361
rect 54 80225 154 80350
rect 151963 79679 152123 79682
rect 151268 79519 151963 79679
rect 151963 79516 152123 79519
rect 54 78961 154 79155
rect 51 78861 54 78961
rect 154 78861 157 78961
rect 51 78850 157 78861
rect 54 78725 154 78850
rect 151963 78179 152123 78182
rect 151268 78019 151963 78179
rect 151963 78016 152123 78019
rect 54 77461 154 77655
rect 51 77361 54 77461
rect 154 77361 157 77461
rect 51 77350 157 77361
rect 54 77225 154 77350
rect 151963 76679 152123 76682
rect 151268 76519 151963 76679
rect 151963 76516 152123 76519
rect 54 75961 154 76155
rect 51 75861 54 75961
rect 154 75861 157 75961
rect 51 75850 157 75861
rect 54 75725 154 75850
rect 151963 75179 152123 75182
rect 151268 75019 151963 75179
rect 151963 75016 152123 75019
rect 54 74461 154 74655
rect 51 74361 54 74461
rect 154 74361 157 74461
rect 51 74350 157 74361
rect 54 74225 154 74350
rect 151963 73679 152123 73682
rect 151268 73519 151963 73679
rect 151963 73516 152123 73519
rect 54 72961 154 73155
rect 51 72861 54 72961
rect 154 72861 157 72961
rect 51 72850 157 72861
rect 54 72725 154 72850
rect 151963 72179 152123 72182
rect 151268 72019 151963 72179
rect 151963 72016 152123 72019
rect 54 71461 154 71655
rect 51 71361 54 71461
rect 154 71361 157 71461
rect 51 71350 157 71361
rect 54 71225 154 71350
rect 151963 70679 152123 70682
rect 151268 70519 151963 70679
rect 151963 70516 152123 70519
rect 54 69961 154 70155
rect 51 69861 54 69961
rect 154 69861 157 69961
rect 51 69850 157 69861
rect 54 69725 154 69850
rect 151963 69179 152123 69182
rect 151268 69019 151963 69179
rect 151963 69016 152123 69019
rect 54 68461 154 68655
rect 51 68361 54 68461
rect 154 68361 157 68461
rect 51 68350 157 68361
rect 54 68225 154 68350
rect 151963 67679 152123 67682
rect 151268 67519 151963 67679
rect 151963 67516 152123 67519
rect 54 66961 154 67155
rect 51 66861 54 66961
rect 154 66861 157 66961
rect 51 66850 157 66861
rect 54 66725 154 66850
rect 151963 66179 152123 66182
rect 151268 66019 151963 66179
rect 151963 66016 152123 66019
rect 54 65461 154 65655
rect 51 65361 54 65461
rect 154 65361 157 65461
rect 51 65350 157 65361
rect 54 65225 154 65350
rect 151963 64679 152123 64682
rect 151268 64519 151963 64679
rect 151963 64516 152123 64519
rect 54 63961 154 64155
rect 51 63861 54 63961
rect 154 63861 157 63961
rect 51 63850 157 63861
rect 54 63725 154 63850
rect 151963 63179 152123 63182
rect 151268 63019 151963 63179
rect 151963 63016 152123 63019
rect 54 62461 154 62655
rect 51 62361 54 62461
rect 154 62361 157 62461
rect 51 62350 157 62361
rect 54 62225 154 62350
rect 151963 61679 152123 61682
rect 151268 61519 151963 61679
rect 151963 61516 152123 61519
rect 54 60961 154 61155
rect 51 60861 54 60961
rect 154 60861 157 60961
rect 51 60850 157 60861
rect 54 60725 154 60850
rect 151963 60179 152123 60182
rect 151268 60019 151963 60179
rect 151963 60016 152123 60019
rect 54 59461 154 59655
rect 51 59361 54 59461
rect 154 59361 157 59461
rect 51 59350 157 59361
rect 54 59225 154 59350
rect 151963 58679 152123 58682
rect 151268 58519 151963 58679
rect 151963 58516 152123 58519
rect 54 57961 154 58155
rect 51 57861 54 57961
rect 154 57861 157 57961
rect 51 57850 157 57861
rect 54 57725 154 57850
rect 151963 57179 152123 57182
rect 151268 57019 151963 57179
rect 151963 57016 152123 57019
rect 54 56461 154 56655
rect 51 56361 54 56461
rect 154 56361 157 56461
rect 51 56350 157 56361
rect 54 56225 154 56350
rect 151963 55679 152123 55682
rect 151268 55519 151963 55679
rect 151963 55516 152123 55519
rect 54 54961 154 55155
rect 51 54861 54 54961
rect 154 54861 157 54961
rect 51 54850 157 54861
rect 54 54725 154 54850
rect 151963 54179 152123 54182
rect 151268 54019 151963 54179
rect 151963 54016 152123 54019
rect 54 53461 154 53655
rect 51 53361 54 53461
rect 154 53361 157 53461
rect 51 53350 157 53361
rect 54 53225 154 53350
rect 151963 52679 152123 52682
rect 151268 52519 151963 52679
rect 151963 52516 152123 52519
rect 54 51961 154 52155
rect 51 51861 54 51961
rect 154 51861 157 51961
rect 51 51850 157 51861
rect 54 51725 154 51850
rect 151963 51179 152123 51182
rect 151268 51019 151963 51179
rect 151963 51016 152123 51019
rect 54 50461 154 50655
rect 51 50361 54 50461
rect 154 50361 157 50461
rect 51 50350 157 50361
rect 54 50225 154 50350
rect 151963 49679 152123 49682
rect 151268 49519 151963 49679
rect 151963 49516 152123 49519
rect 54 48961 154 49155
rect 51 48861 54 48961
rect 154 48861 157 48961
rect 51 48850 157 48861
rect 54 48725 154 48850
rect 151963 48179 152123 48182
rect 151268 48019 151963 48179
rect 151963 48016 152123 48019
rect 54 47461 154 47655
rect 51 47361 54 47461
rect 154 47361 157 47461
rect 51 47350 157 47361
rect 54 47225 154 47350
rect 151963 46679 152123 46682
rect 151268 46519 151963 46679
rect 151963 46516 152123 46519
rect 54 45961 154 46155
rect 51 45861 54 45961
rect 154 45861 157 45961
rect 51 45850 157 45861
rect 54 45725 154 45850
rect 151963 45179 152123 45182
rect 151268 45019 151963 45179
rect 151963 45016 152123 45019
rect 54 44461 154 44655
rect 51 44361 54 44461
rect 154 44361 157 44461
rect 51 44350 157 44361
rect 54 44225 154 44350
rect 151963 43679 152123 43682
rect 151268 43519 151963 43679
rect 151963 43516 152123 43519
rect 54 42961 154 43155
rect 51 42861 54 42961
rect 154 42861 157 42961
rect 51 42850 157 42861
rect 54 42725 154 42850
rect 151963 42179 152123 42182
rect 151268 42019 151963 42179
rect 151963 42016 152123 42019
rect 54 41461 154 41655
rect 51 41361 54 41461
rect 154 41361 157 41461
rect 51 41350 157 41361
rect 54 41225 154 41350
rect 151963 40679 152123 40682
rect 151268 40519 151963 40679
rect 151963 40516 152123 40519
rect 54 39961 154 40155
rect 51 39861 54 39961
rect 154 39861 157 39961
rect 51 39850 157 39861
rect 54 39725 154 39850
rect 151963 39179 152123 39182
rect 151268 39019 151963 39179
rect 151963 39016 152123 39019
rect 54 38461 154 38655
rect 51 38361 54 38461
rect 154 38361 157 38461
rect 51 38350 157 38361
rect 54 38225 154 38350
rect 151963 37679 152123 37682
rect 151268 37519 151963 37679
rect 151963 37516 152123 37519
rect 54 36961 154 37155
rect 51 36861 54 36961
rect 154 36861 157 36961
rect 51 36850 157 36861
rect 54 36725 154 36850
rect 151963 36179 152123 36182
rect 151268 36019 151963 36179
rect 151963 36016 152123 36019
rect 54 35461 154 35655
rect 51 35361 54 35461
rect 154 35361 157 35461
rect 51 35350 157 35361
rect 54 35225 154 35350
rect 151963 34679 152123 34682
rect 151268 34519 151963 34679
rect 151963 34516 152123 34519
rect 54 33961 154 34155
rect 51 33861 54 33961
rect 154 33861 157 33961
rect 51 33850 157 33861
rect 54 33725 154 33850
rect 151963 33179 152123 33182
rect 151268 33019 151963 33179
rect 151963 33016 152123 33019
rect 54 32461 154 32655
rect 51 32361 54 32461
rect 154 32361 157 32461
rect 51 32350 157 32361
rect 54 32225 154 32350
rect 151963 31679 152123 31682
rect 151268 31519 151963 31679
rect 151963 31516 152123 31519
rect 54 30961 154 31155
rect 51 30861 54 30961
rect 154 30861 157 30961
rect 51 30850 157 30861
rect 54 30725 154 30850
rect 151963 30179 152123 30182
rect 151268 30019 151963 30179
rect 151963 30016 152123 30019
rect 54 29461 154 29655
rect 51 29361 54 29461
rect 154 29361 157 29461
rect 51 29350 157 29361
rect 54 29225 154 29350
rect 151963 28679 152123 28682
rect 151268 28519 151963 28679
rect 151963 28516 152123 28519
rect 54 27961 154 28155
rect 51 27861 54 27961
rect 154 27861 157 27961
rect 51 27850 157 27861
rect 54 27725 154 27850
rect 151963 27179 152123 27182
rect 151268 27019 151963 27179
rect 151963 27016 152123 27019
rect 54 26461 154 26655
rect 51 26361 54 26461
rect 154 26361 157 26461
rect 51 26350 157 26361
rect 54 26225 154 26350
rect 151963 25679 152123 25682
rect 151268 25519 151963 25679
rect 151963 25516 152123 25519
rect 54 24961 154 25155
rect 51 24861 54 24961
rect 154 24861 157 24961
rect 51 24850 157 24861
rect 54 24725 154 24850
rect 151963 24179 152123 24182
rect 151268 24019 151963 24179
rect 151963 24016 152123 24019
rect 54 23461 154 23655
rect 51 23361 54 23461
rect 154 23361 157 23461
rect 51 23350 157 23361
rect 54 23225 154 23350
rect 151963 22679 152123 22682
rect 151268 22519 151963 22679
rect 151963 22516 152123 22519
rect 54 21961 154 22155
rect 51 21861 54 21961
rect 154 21861 157 21961
rect 51 21850 157 21861
rect 54 21725 154 21850
rect 151963 21179 152123 21182
rect 151268 21019 151963 21179
rect 151963 21016 152123 21019
rect 54 20461 154 20655
rect 51 20361 54 20461
rect 154 20361 157 20461
rect 51 20350 157 20361
rect 54 20225 154 20350
rect 151963 19679 152123 19682
rect 151268 19519 151963 19679
rect 151963 19516 152123 19519
rect 54 18961 154 19155
rect 51 18861 54 18961
rect 154 18861 157 18961
rect 51 18850 157 18861
rect 54 18725 154 18850
rect 151963 18179 152123 18182
rect 151268 18019 151963 18179
rect 151963 18016 152123 18019
rect 54 17461 154 17655
rect 51 17361 54 17461
rect 154 17361 157 17461
rect 51 17350 157 17361
rect 54 17225 154 17350
rect 151963 16679 152123 16682
rect 151268 16519 151963 16679
rect 151963 16516 152123 16519
rect 54 15961 154 16155
rect 51 15861 54 15961
rect 154 15861 157 15961
rect 51 15850 157 15861
rect 54 15725 154 15850
rect 151963 15179 152123 15182
rect 151268 15019 151963 15179
rect 151963 15016 152123 15019
rect 54 14461 154 14655
rect 51 14361 54 14461
rect 154 14361 157 14461
rect 51 14350 157 14361
rect 54 14225 154 14350
rect 151963 13679 152123 13682
rect 151268 13519 151963 13679
rect 151963 13516 152123 13519
rect 54 12961 154 13155
rect 51 12861 54 12961
rect 154 12861 157 12961
rect 51 12850 157 12861
rect 54 12725 154 12850
rect 151963 12179 152123 12182
rect 151268 12019 151963 12179
rect 151963 12016 152123 12019
rect 54 11461 154 11655
rect 51 11361 54 11461
rect 154 11361 157 11461
rect 51 11350 157 11361
rect 54 11225 154 11350
rect 151963 10679 152123 10682
rect 151268 10519 151963 10679
rect 151963 10516 152123 10519
rect 54 9950 154 10404
rect 151254 10204 151414 10304
rect 51 9850 157 9950
rect 54 8973 154 9850
rect 1829 9220 1832 9380
rect 1992 9220 1995 9380
rect 9041 9220 9044 9380
rect 9204 9220 9207 9380
rect 16454 9220 16457 9380
rect 16617 9220 16620 9380
rect 32125 9220 32128 9380
rect 32288 9220 32291 9380
rect 60836 9220 60839 9380
rect 60999 9220 61002 9380
rect 83771 9220 83774 9380
rect 83934 9220 83937 9380
rect 90271 9220 90274 9380
rect 90434 9220 90437 9380
rect 94771 9220 94774 9380
rect 94934 9220 94937 9380
rect 99271 9220 99274 9380
rect 99434 9220 99437 9380
rect 102271 9220 102274 9380
rect 102434 9220 102437 9380
rect 105771 9220 105774 9380
rect 105934 9220 105937 9380
rect 111771 9220 111774 9380
rect 111934 9220 111937 9380
rect 116271 9220 116274 9380
rect 116434 9220 116437 9380
rect 119271 9220 119274 9380
rect 119434 9220 119437 9380
rect 125271 9220 125274 9380
rect 125434 9220 125437 9380
rect 131971 9220 131974 9380
rect 132134 9220 132137 9380
rect 134971 9220 134974 9380
rect 135134 9220 135137 9380
rect 136471 9220 136474 9380
rect 136634 9220 136637 9380
rect 137971 9220 137974 9380
rect 138134 9220 138137 9380
rect 140971 9220 140974 9380
rect 141134 9220 141137 9380
rect 142971 9220 142974 9380
rect 143134 9220 143137 9380
rect 146971 9220 146974 9380
rect 147134 9220 147137 9380
rect 148471 9220 148474 9380
rect 148634 9220 148637 9380
rect 149971 9220 149974 9380
rect 150134 9220 150137 9380
rect 151471 9220 151474 9380
rect 151634 9220 151637 9380
rect -3102 8873 -3099 8973
rect -2999 8873 154 8973
rect 1832 8969 1992 9220
rect 9044 8969 9204 9220
rect 16457 8969 16617 9220
rect 32128 8969 32288 9220
rect 60839 8969 60999 9220
rect 83774 8969 83934 9220
rect 90274 8969 90434 9220
rect 94774 8969 94934 9220
rect 99274 8969 99434 9220
rect 102274 8969 102434 9220
rect 105774 8969 105934 9220
rect 111774 8969 111934 9220
rect 116274 8969 116434 9220
rect 119274 8969 119434 9220
rect 125274 8969 125434 9220
rect 131974 8969 132134 9220
rect 134974 8969 135134 9220
rect 136474 8969 136634 9220
rect 137974 8969 138134 9220
rect 140974 8969 141134 9220
rect 142974 8969 143134 9220
rect 146974 8969 147134 9220
rect 148474 8969 148634 9220
rect 149974 8969 150134 9220
rect 151474 9129 151634 9220
rect 54 7794 154 8873
rect 151473 8208 151634 9129
rect 151473 8044 151634 8047
rect 54 7691 154 7694
<< via1 >>
rect 151254 162166 151354 162266
rect 151963 160519 152123 160679
rect 54 159861 154 159961
rect 151963 159019 152123 159179
rect 54 158361 154 158461
rect 151963 157519 152123 157679
rect 54 156861 154 156961
rect 151963 156019 152123 156179
rect 54 155361 154 155461
rect 151963 154519 152123 154679
rect 54 153861 154 153961
rect 151963 153019 152123 153179
rect 54 152361 154 152461
rect 151963 151519 152123 151679
rect 54 150861 154 150961
rect 151963 150019 152123 150179
rect 54 149361 154 149461
rect 151963 148519 152123 148679
rect 54 147861 154 147961
rect 151963 147019 152123 147179
rect 54 146361 154 146461
rect 151963 145519 152123 145679
rect 54 144861 154 144961
rect 151963 144019 152123 144179
rect 54 143361 154 143461
rect 151963 142519 152123 142679
rect 54 141861 154 141961
rect 151963 141019 152123 141179
rect 54 140361 154 140461
rect 151963 139519 152123 139679
rect 54 138861 154 138961
rect 151963 138019 152123 138179
rect 54 137361 154 137461
rect 151963 136519 152123 136679
rect 54 135861 154 135961
rect 151963 135019 152123 135179
rect 54 134361 154 134461
rect 151963 133519 152123 133679
rect 54 132861 154 132961
rect 151963 132019 152123 132179
rect 54 131361 154 131461
rect 151963 130519 152123 130679
rect 54 129861 154 129961
rect 151963 129019 152123 129179
rect 54 128361 154 128461
rect 151963 127519 152123 127679
rect 54 126861 154 126961
rect 151963 126019 152123 126179
rect 54 125361 154 125461
rect 151963 124519 152123 124679
rect 54 123861 154 123961
rect 151963 123019 152123 123179
rect 54 122361 154 122461
rect 151963 121519 152123 121679
rect 54 120861 154 120961
rect 151963 120019 152123 120179
rect 54 119361 154 119461
rect 151963 118519 152123 118679
rect 54 117861 154 117961
rect 151963 117019 152123 117179
rect 54 116361 154 116461
rect 151963 115519 152123 115679
rect 54 114861 154 114961
rect 151963 114019 152123 114179
rect 54 113361 154 113461
rect 151963 112519 152123 112679
rect 54 111861 154 111961
rect 151963 111019 152123 111179
rect 54 110361 154 110461
rect 151963 109519 152123 109679
rect 54 108861 154 108961
rect 151963 108019 152123 108179
rect 54 107361 154 107461
rect 151963 106519 152123 106679
rect 54 105861 154 105961
rect 151963 105019 152123 105179
rect 54 104361 154 104461
rect 151963 103519 152123 103679
rect 54 102861 154 102961
rect 151963 102019 152123 102179
rect 54 101361 154 101461
rect 151963 100519 152123 100679
rect 54 99861 154 99961
rect 151963 99019 152123 99179
rect 54 98361 154 98461
rect 151963 97519 152123 97679
rect 54 96861 154 96961
rect 151963 96019 152123 96179
rect 54 95361 154 95461
rect 151963 94519 152123 94679
rect 54 93861 154 93961
rect 151963 93019 152123 93179
rect 54 92361 154 92461
rect 151963 91519 152123 91679
rect 54 90861 154 90961
rect 151963 90019 152123 90179
rect 54 89361 154 89461
rect 151963 88519 152123 88679
rect 54 87861 154 87961
rect 151963 87019 152123 87179
rect 54 86361 154 86461
rect 151963 85519 152123 85679
rect 54 84861 154 84961
rect 151963 84019 152123 84179
rect 54 83361 154 83461
rect 151963 82519 152123 82679
rect 54 81861 154 81961
rect 151963 81019 152123 81179
rect 54 80361 154 80461
rect 151963 79519 152123 79679
rect 54 78861 154 78961
rect 151963 78019 152123 78179
rect 54 77361 154 77461
rect 151963 76519 152123 76679
rect 54 75861 154 75961
rect 151963 75019 152123 75179
rect 54 74361 154 74461
rect 151963 73519 152123 73679
rect 54 72861 154 72961
rect 151963 72019 152123 72179
rect 54 71361 154 71461
rect 151963 70519 152123 70679
rect 54 69861 154 69961
rect 151963 69019 152123 69179
rect 54 68361 154 68461
rect 151963 67519 152123 67679
rect 54 66861 154 66961
rect 151963 66019 152123 66179
rect 54 65361 154 65461
rect 151963 64519 152123 64679
rect 54 63861 154 63961
rect 151963 63019 152123 63179
rect 54 62361 154 62461
rect 151963 61519 152123 61679
rect 54 60861 154 60961
rect 151963 60019 152123 60179
rect 54 59361 154 59461
rect 151963 58519 152123 58679
rect 54 57861 154 57961
rect 151963 57019 152123 57179
rect 54 56361 154 56461
rect 151963 55519 152123 55679
rect 54 54861 154 54961
rect 151963 54019 152123 54179
rect 54 53361 154 53461
rect 151963 52519 152123 52679
rect 54 51861 154 51961
rect 151963 51019 152123 51179
rect 54 50361 154 50461
rect 151963 49519 152123 49679
rect 54 48861 154 48961
rect 151963 48019 152123 48179
rect 54 47361 154 47461
rect 151963 46519 152123 46679
rect 54 45861 154 45961
rect 151963 45019 152123 45179
rect 54 44361 154 44461
rect 151963 43519 152123 43679
rect 54 42861 154 42961
rect 151963 42019 152123 42179
rect 54 41361 154 41461
rect 151963 40519 152123 40679
rect 54 39861 154 39961
rect 151963 39019 152123 39179
rect 54 38361 154 38461
rect 151963 37519 152123 37679
rect 54 36861 154 36961
rect 151963 36019 152123 36179
rect 54 35361 154 35461
rect 151963 34519 152123 34679
rect 54 33861 154 33961
rect 151963 33019 152123 33179
rect 54 32361 154 32461
rect 151963 31519 152123 31679
rect 54 30861 154 30961
rect 151963 30019 152123 30179
rect 54 29361 154 29461
rect 151963 28519 152123 28679
rect 54 27861 154 27961
rect 151963 27019 152123 27179
rect 54 26361 154 26461
rect 151963 25519 152123 25679
rect 54 24861 154 24961
rect 151963 24019 152123 24179
rect 54 23361 154 23461
rect 151963 22519 152123 22679
rect 54 21861 154 21961
rect 151963 21019 152123 21179
rect 54 20361 154 20461
rect 151963 19519 152123 19679
rect 54 18861 154 18961
rect 151963 18019 152123 18179
rect 54 17361 154 17461
rect 151963 16519 152123 16679
rect 54 15861 154 15961
rect 151963 15019 152123 15179
rect 54 14361 154 14461
rect 151963 13519 152123 13679
rect 54 12861 154 12961
rect 151963 12019 152123 12179
rect 54 11361 154 11461
rect 151963 10519 152123 10679
rect 1832 9220 1992 9380
rect 9044 9220 9204 9380
rect 16457 9220 16617 9380
rect 32128 9220 32288 9380
rect 60839 9220 60999 9380
rect 83774 9220 83934 9380
rect 90274 9220 90434 9380
rect 94774 9220 94934 9380
rect 99274 9220 99434 9380
rect 102274 9220 102434 9380
rect 105774 9220 105934 9380
rect 111774 9220 111934 9380
rect 116274 9220 116434 9380
rect 119274 9220 119434 9380
rect 125274 9220 125434 9380
rect 131974 9220 132134 9380
rect 134974 9220 135134 9380
rect 136474 9220 136634 9380
rect 137974 9220 138134 9380
rect 140974 9220 141134 9380
rect 142974 9220 143134 9380
rect 146974 9220 147134 9380
rect 148474 9220 148634 9380
rect 149974 9220 150134 9380
rect 151474 9220 151634 9380
rect -3099 8873 -2999 8973
rect 151473 8047 151634 8208
rect 54 7694 154 7794
<< metal2 >>
rect -4083 162690 -813 162745
rect -2590 161221 -1016 161266
rect -2566 159701 -1201 159729
rect -2584 158183 -1371 158211
rect -2574 156619 -1551 156647
rect -1767 155129 -1722 155137
rect -2574 155101 -1722 155129
rect -2569 153583 -1966 153611
rect -2579 152019 -2171 152047
rect -2199 151169 -2171 152019
rect -1994 151974 -1966 153583
rect -1767 153474 -1722 155101
rect -1579 154974 -1551 156619
rect -1399 156474 -1371 158183
rect -1229 157965 -1201 159701
rect -1061 159474 -1016 161221
rect -868 160419 -813 162690
rect 679 160619 734 163560
rect 1059 160709 1114 163498
rect 151254 162266 151354 162271
rect 151251 162166 151254 162266
rect 151354 162166 151357 162266
rect 151254 162162 151354 162166
rect 151965 160679 152120 160681
rect 151960 160519 151963 160679
rect 152123 160519 152126 160679
rect 151965 160517 152120 160519
rect -868 160364 -391 160419
rect 54 159961 154 159964
rect 49 159861 54 159961
rect 154 159861 158 159961
rect 54 159858 154 159861
rect -1061 159429 -401 159474
rect 151965 159179 152120 159181
rect 151960 159019 151963 159179
rect 152123 159019 152126 159179
rect 151965 159017 152120 159019
rect 54 158461 154 158464
rect 49 158361 54 158461
rect 154 158361 158 158461
rect 54 158358 154 158361
rect -1229 157937 -289 157965
rect 151965 157679 152120 157681
rect 151960 157519 151963 157679
rect 152123 157519 152126 157679
rect 151965 157517 152120 157519
rect 54 156961 154 156964
rect 49 156861 54 156961
rect 154 156861 158 156961
rect 54 156858 154 156861
rect -1399 156446 -311 156474
rect 151965 156179 152120 156181
rect 151960 156019 151963 156179
rect 152123 156019 152126 156179
rect 151965 156017 152120 156019
rect 54 155461 154 155464
rect 49 155361 54 155461
rect 154 155361 158 155461
rect 54 155358 154 155361
rect -1582 154929 -377 154974
rect 151965 154679 152120 154681
rect 151960 154519 151963 154679
rect 152123 154519 152126 154679
rect 151965 154517 152120 154519
rect 54 153961 154 153964
rect 49 153861 54 153961
rect 154 153861 158 153961
rect 54 153858 154 153861
rect -1767 153429 -401 153474
rect 151965 153179 152120 153181
rect 151960 153019 151963 153179
rect 152123 153019 152126 153179
rect 151965 153017 152120 153019
rect 54 152461 154 152464
rect 49 152361 54 152461
rect 154 152361 158 152461
rect 54 152358 154 152361
rect -2002 151929 -387 151974
rect 151965 151679 152120 151681
rect 151960 151519 151963 151679
rect 152123 151519 152126 151679
rect 151965 151517 152120 151519
rect -2199 151141 -346 151169
rect -742 150529 -502 150532
rect -2564 150501 -502 150529
rect -742 150487 -502 150501
rect -2574 148983 -771 149011
rect -817 147474 -772 148983
rect -547 148974 -502 150487
rect -417 150429 -372 151141
rect 54 150961 154 150964
rect 49 150861 54 150961
rect 154 150861 158 150961
rect 54 150858 154 150861
rect 151965 150179 152120 150181
rect 151960 150019 151963 150179
rect 152123 150019 152126 150179
rect 151965 150017 152120 150019
rect 54 149461 154 149464
rect 49 149361 54 149461
rect 154 149361 158 149461
rect 54 149358 154 149361
rect -547 148929 -372 148974
rect 151965 148679 152120 148681
rect 151960 148519 151963 148679
rect 152123 148519 152126 148679
rect 151965 148517 152120 148519
rect 54 147961 154 147964
rect 49 147861 54 147961
rect 154 147861 158 147961
rect 54 147858 154 147861
rect -2574 147419 -1076 147447
rect -817 147429 -362 147474
rect -1547 145929 -1502 146027
rect -1104 145959 -1076 147419
rect 151965 147179 152120 147181
rect 151960 147019 151963 147179
rect 152123 147019 152126 147179
rect 151965 147017 152120 147019
rect 54 146461 154 146464
rect 49 146361 54 146461
rect 154 146361 158 146461
rect 54 146358 154 146361
rect -1104 145931 -226 145959
rect -2574 145901 -1502 145929
rect -1547 144474 -1502 145901
rect 151965 145679 152120 145681
rect 151960 145519 151963 145679
rect 152123 145519 152126 145679
rect 151965 145517 152120 145519
rect 54 144961 154 144964
rect 49 144861 54 144961
rect 154 144861 158 144961
rect 54 144858 154 144861
rect -1547 144429 -392 144474
rect -1957 144365 -1912 144407
rect -2574 144337 -1912 144365
rect -1957 142974 -1912 144337
rect 151965 144179 152120 144181
rect 151960 144019 151963 144179
rect 152123 144019 152126 144179
rect 151965 144017 152120 144019
rect 54 143461 154 143464
rect 49 143361 54 143461
rect 154 143361 158 143461
rect 54 143358 154 143361
rect -1957 142929 -382 142974
rect -2569 142819 -2116 142847
rect -2144 142044 -2116 142819
rect 151965 142679 152120 142681
rect 151960 142519 151963 142679
rect 152123 142519 152126 142679
rect 151965 142517 152120 142519
rect -552 142044 -507 142052
rect -2144 142016 -481 142044
rect -552 141474 -507 142016
rect 54 141961 154 141964
rect 49 141861 54 141961
rect 154 141861 158 141961
rect 54 141858 154 141861
rect -552 141429 -401 141474
rect -1102 141329 -1057 141382
rect -2579 141301 -1057 141329
rect -1102 139974 -1057 141301
rect 151965 141179 152120 141181
rect 151960 141019 151963 141179
rect 152123 141019 152126 141179
rect 151965 141017 152120 141019
rect 54 140461 154 140464
rect 49 140361 54 140461
rect 154 140361 158 140461
rect 54 140358 154 140361
rect -1102 139929 -401 139974
rect -2609 139737 -981 139765
rect -1027 138474 -982 139737
rect 151965 139679 152120 139681
rect 151960 139519 151963 139679
rect 152123 139519 152126 139679
rect 151965 139517 152120 139519
rect 54 138961 154 138964
rect 49 138861 54 138961
rect 154 138861 158 138961
rect 54 138858 154 138861
rect -1027 138429 -392 138474
rect -446 138247 -401 138262
rect -2594 138219 -401 138247
rect -446 136929 -401 138219
rect 151965 138179 152120 138181
rect 151960 138019 151963 138179
rect 152123 138019 152126 138179
rect 151965 138017 152120 138019
rect 54 137461 154 137464
rect 49 137361 54 137461
rect 154 137361 158 137461
rect 54 137358 154 137361
rect -1982 136729 -1937 136792
rect -2614 136701 -1937 136729
rect -1982 135474 -1937 136701
rect 151965 136679 152120 136681
rect 151960 136519 151963 136679
rect 152123 136519 152126 136679
rect 151965 136517 152120 136519
rect 54 135961 154 135964
rect 49 135861 54 135961
rect 154 135861 158 135961
rect 54 135858 154 135861
rect -1982 135429 -401 135474
rect 151965 135179 152120 135181
rect -2584 135137 -2291 135165
rect -2319 133974 -2291 135137
rect 151960 135019 151963 135179
rect 152123 135019 152126 135179
rect 151965 135017 152120 135019
rect 54 134461 154 134464
rect 49 134361 54 134461
rect 154 134361 158 134461
rect 54 134358 154 134361
rect -2319 133941 -401 133974
rect -2307 133929 -401 133941
rect -2142 133647 -2097 133712
rect 151965 133679 152120 133681
rect -2574 133619 -2097 133647
rect -2142 132474 -2097 133619
rect 151960 133519 151963 133679
rect 152123 133519 152126 133679
rect 151965 133517 152120 133519
rect 54 132961 154 132964
rect 49 132861 54 132961
rect 154 132861 158 132961
rect 54 132858 154 132861
rect -2142 132429 -401 132474
rect 151965 132179 152120 132181
rect -2574 132055 -966 132083
rect -994 130974 -966 132055
rect 151960 132019 151963 132179
rect 152123 132019 152126 132179
rect 151965 132017 152120 132019
rect 54 131461 154 131464
rect 49 131361 54 131461
rect 154 131361 158 131461
rect 54 131358 154 131361
rect -994 130929 -401 130974
rect -994 130906 -966 130929
rect 151965 130679 152120 130681
rect -2589 130537 -546 130565
rect -574 129474 -546 130537
rect 151960 130519 151963 130679
rect 152123 130519 152126 130679
rect 151965 130517 152120 130519
rect 54 129961 154 129964
rect 49 129861 54 129961
rect 154 129861 158 129961
rect 54 129858 154 129861
rect -574 129429 -387 129474
rect -574 129411 -546 129429
rect 151965 129179 152120 129181
rect -2609 129019 -556 129047
rect 151960 129019 151963 129179
rect 152123 129019 152126 129179
rect -584 127974 -556 129019
rect 151965 129017 152120 129019
rect 54 128461 154 128464
rect 49 128361 54 128461
rect 154 128361 158 128461
rect 54 128358 154 128361
rect -584 127929 -401 127974
rect -584 127921 -556 127929
rect 151965 127679 152120 127681
rect 151960 127519 151963 127679
rect 152123 127519 152126 127679
rect 151965 127517 152120 127519
rect -2584 127455 -586 127483
rect -614 126474 -586 127455
rect 54 126961 154 126964
rect 49 126861 54 126961
rect 154 126861 158 126961
rect 54 126858 154 126861
rect -614 126429 -401 126474
rect -614 126426 -586 126429
rect 151965 126179 152120 126181
rect 151960 126019 151963 126179
rect 152123 126019 152126 126179
rect 151965 126017 152120 126019
rect -2604 125937 -701 125965
rect -729 124974 -701 125937
rect 54 125461 154 125464
rect 49 125361 54 125461
rect 154 125361 158 125461
rect 54 125358 154 125361
rect -729 124946 -397 124974
rect -717 124929 -397 124946
rect 151965 124679 152120 124681
rect -442 124447 -397 124542
rect 151960 124519 151963 124679
rect 152123 124519 152126 124679
rect 151965 124517 152120 124519
rect -2564 124419 -396 124447
rect -442 123429 -397 124419
rect 54 123961 154 123964
rect 49 123861 54 123961
rect 154 123861 158 123961
rect 54 123858 154 123861
rect 151965 123179 152120 123181
rect 151960 123019 151963 123179
rect 152123 123019 152126 123179
rect 151965 123017 152120 123019
rect -446 122883 -401 122942
rect -2634 122855 -401 122883
rect -446 121929 -401 122855
rect 54 122461 154 122464
rect 49 122361 54 122461
rect 154 122361 158 122461
rect 54 122358 154 122361
rect 151965 121679 152120 121681
rect 151960 121519 151963 121679
rect 152123 121519 152126 121679
rect 151965 121517 152120 121519
rect -2614 121337 -416 121365
rect -444 120426 -416 121337
rect 54 120961 154 120964
rect 49 120861 54 120961
rect 154 120861 158 120961
rect 54 120858 154 120861
rect 151965 120179 152120 120181
rect 151960 120019 151963 120179
rect 152123 120019 152126 120179
rect 151965 120017 152120 120019
rect -2579 119819 -406 119847
rect -434 118946 -406 119819
rect 54 119461 154 119464
rect 49 119361 54 119461
rect 154 119361 158 119461
rect 54 119358 154 119361
rect 151965 118679 152120 118681
rect 151960 118519 151963 118679
rect 152123 118519 152126 118679
rect 151965 118517 152120 118519
rect -446 118283 -401 118362
rect -2594 118255 -401 118283
rect -446 117429 -401 118255
rect 54 117961 154 117964
rect 49 117861 54 117961
rect 154 117861 158 117961
rect 54 117858 154 117861
rect 151965 117179 152120 117181
rect 151960 117019 151963 117179
rect 152123 117019 152126 117179
rect 151965 117017 152120 117019
rect -2584 116737 -446 116765
rect -474 115926 -446 116737
rect 54 116461 154 116464
rect 49 116361 54 116461
rect 154 116361 158 116461
rect 54 116358 154 116361
rect 151965 115679 152120 115681
rect 151960 115519 151963 115679
rect 152123 115519 152126 115679
rect 151965 115517 152120 115519
rect -2584 114474 -2556 115201
rect 54 114961 154 114964
rect 49 114861 54 114961
rect 154 114861 158 114961
rect 54 114858 154 114861
rect -2584 114446 -392 114474
rect -2577 114429 -392 114446
rect 151965 114179 152120 114181
rect 151960 114019 151963 114179
rect 152123 114019 152126 114179
rect 151965 114017 152120 114019
rect -2569 113655 -306 113683
rect -417 112929 -372 113655
rect 54 113461 154 113464
rect 49 113361 54 113461
rect 154 113361 158 113461
rect 54 113358 154 113361
rect 151965 112679 152120 112681
rect 151960 112519 151963 112679
rect 152123 112519 152126 112679
rect 151965 112517 152120 112519
rect -2597 112132 -401 112177
rect -446 111429 -401 112132
rect 54 111961 154 111964
rect 49 111861 54 111961
rect 154 111861 158 111961
rect 54 111858 154 111861
rect 151965 111179 152120 111181
rect 151960 111019 151963 111179
rect 152123 111019 152126 111179
rect 151965 111017 152120 111019
rect -2574 110573 -404 110601
rect -432 109941 -404 110573
rect 54 110461 154 110464
rect 49 110361 54 110461
rect 154 110361 158 110461
rect 54 110358 154 110361
rect 151965 109679 152120 109681
rect 151960 109519 151963 109679
rect 152123 109519 152126 109679
rect 151965 109517 152120 109519
rect -404 109089 -376 109101
rect -2564 109061 -376 109089
rect -404 108436 -376 109061
rect 54 108961 154 108964
rect 49 108861 54 108961
rect 154 108861 158 108961
rect 54 108858 154 108861
rect 151965 108179 152120 108181
rect 151960 108019 151963 108179
rect 152123 108019 152126 108179
rect 151965 108017 152120 108019
rect -2564 107541 -376 107569
rect -404 106929 -376 107541
rect 54 107461 154 107464
rect 49 107361 54 107461
rect 154 107361 158 107461
rect 54 107358 154 107361
rect 151965 106679 152120 106681
rect 151960 106519 151963 106679
rect 152123 106519 152126 106679
rect 151965 106517 152120 106519
rect -2567 105957 -401 106002
rect 54 105961 154 105964
rect -446 105429 -401 105957
rect 49 105861 54 105961
rect 154 105861 158 105961
rect 54 105858 154 105861
rect 151965 105179 152120 105181
rect 151960 105019 151963 105179
rect 152123 105019 152126 105179
rect 151965 105017 152120 105019
rect -2564 104455 -366 104483
rect 54 104461 154 104464
rect -446 103936 -366 104455
rect 49 104361 54 104461
rect 154 104361 158 104461
rect 54 104358 154 104361
rect -446 103929 -382 103936
rect 151965 103679 152120 103681
rect 151960 103519 151963 103679
rect 152123 103519 152126 103679
rect 151965 103517 152120 103519
rect 54 102961 154 102964
rect -2584 102891 -401 102919
rect -429 102421 -401 102891
rect 49 102861 54 102961
rect 154 102861 158 102961
rect 54 102858 154 102861
rect 151965 102179 152120 102181
rect 151960 102019 151963 102179
rect 152123 102019 152126 102179
rect 151965 102017 152120 102019
rect 54 101461 154 101464
rect -2579 101373 -381 101401
rect -442 100929 -397 101373
rect 49 101361 54 101461
rect 154 101361 158 101461
rect 54 101358 154 101361
rect 151965 100679 152120 100681
rect 151960 100519 151963 100679
rect 152123 100519 152126 100679
rect 151965 100517 152120 100519
rect 54 99961 154 99964
rect -2604 99855 -361 99883
rect 49 99861 54 99961
rect 154 99861 158 99961
rect 54 99858 154 99861
rect -389 99426 -361 99855
rect 151965 99179 152120 99181
rect 151960 99019 151963 99179
rect 152123 99019 152126 99179
rect 151965 99017 152120 99019
rect 54 98461 154 98464
rect 49 98361 54 98461
rect 154 98361 158 98461
rect 54 98358 154 98361
rect -2572 98291 -601 98319
rect -629 97974 -601 98291
rect -629 97929 -396 97974
rect -629 97902 -601 97929
rect 151965 97679 152120 97681
rect 151960 97519 151963 97679
rect 152123 97519 152126 97679
rect 151965 97517 152120 97519
rect 54 96961 154 96964
rect 49 96861 54 96961
rect 154 96861 158 96961
rect 54 96858 154 96861
rect -2572 96776 -2445 96821
rect -2490 96474 -2445 96776
rect -2490 96429 -391 96474
rect 151965 96179 152120 96181
rect 151960 96019 151963 96179
rect 152123 96019 152126 96179
rect 151965 96017 152120 96019
rect 54 95461 154 95464
rect 49 95361 54 95461
rect 154 95361 158 95461
rect 54 95358 154 95361
rect -2567 95255 -368 95283
rect -396 94903 -368 95255
rect 151965 94679 152120 94681
rect 151960 94519 151963 94679
rect 152123 94519 152126 94679
rect 151965 94517 152120 94519
rect 54 93961 154 93964
rect 49 93861 54 93961
rect 154 93861 158 93961
rect 54 93858 154 93861
rect -2570 93474 -2525 93730
rect -2570 93429 -396 93474
rect 151965 93179 152120 93181
rect 151960 93019 151963 93179
rect 152123 93019 152126 93179
rect 151965 93017 152120 93019
rect 54 92461 154 92464
rect 49 92361 54 92461
rect 154 92361 158 92461
rect 54 92358 154 92361
rect -2570 91974 -2525 92212
rect -2570 91929 -289 91974
rect 151965 91679 152120 91681
rect 151960 91519 151963 91679
rect 152123 91519 152126 91679
rect 151965 91517 152120 91519
rect 54 90961 154 90964
rect 49 90861 54 90961
rect 154 90861 158 90961
rect 54 90858 154 90861
rect -2592 90474 -2547 90669
rect -2592 90429 -401 90474
rect 151965 90179 152120 90181
rect 151960 90019 151963 90179
rect 152123 90019 152126 90179
rect 151965 90017 152120 90019
rect 54 89461 154 89464
rect 49 89361 54 89461
rect 154 89361 158 89461
rect 54 89358 154 89361
rect -2584 88974 -2539 89117
rect -2584 88929 -286 88974
rect 151965 88679 152120 88681
rect 151960 88519 151963 88679
rect 152123 88519 152126 88679
rect 151965 88517 152120 88519
rect 54 87961 154 87964
rect 49 87861 54 87961
rect 154 87861 158 87961
rect 54 87858 154 87861
rect -2564 87474 -2536 87601
rect -2564 87429 -345 87474
rect -2564 87395 -2536 87429
rect 151965 87179 152120 87181
rect 151960 87019 151963 87179
rect 152123 87019 152126 87179
rect 151965 87017 152120 87019
rect 54 86461 154 86464
rect 49 86361 54 86461
rect 154 86361 158 86461
rect 54 86358 154 86361
rect -2604 85974 -2559 86032
rect -2604 85929 -391 85974
rect 151965 85679 152120 85681
rect 151960 85519 151963 85679
rect 152123 85519 152126 85679
rect 151965 85517 152120 85519
rect 54 84961 154 84964
rect 49 84861 54 84961
rect 154 84861 158 84961
rect 54 84858 154 84861
rect -2578 84474 -2533 84540
rect -2578 84429 -401 84474
rect 151965 84179 152120 84181
rect 151960 84019 151963 84179
rect 152123 84019 152126 84179
rect 151965 84017 152120 84019
rect 54 83461 154 83464
rect 49 83361 54 83461
rect 154 83361 158 83461
rect 54 83358 154 83361
rect -2572 82974 -2527 83016
rect -2572 82929 -365 82974
rect 151965 82679 152120 82681
rect 151960 82519 151963 82679
rect 152123 82519 152126 82679
rect 151965 82517 152120 82519
rect 54 81961 154 81964
rect 49 81861 54 81961
rect 154 81861 158 81961
rect 54 81858 154 81861
rect -2572 81429 -385 81474
rect 151965 81179 152120 81181
rect 151960 81019 151963 81179
rect 152123 81019 152126 81179
rect 151965 81017 152120 81019
rect 54 80461 154 80464
rect 49 80361 54 80461
rect 154 80361 158 80461
rect 54 80358 154 80361
rect -2961 79929 -399 79974
rect -2961 79889 -408 79929
rect 151965 79679 152120 79681
rect 151960 79519 151963 79679
rect 152123 79519 152126 79679
rect 151965 79517 152120 79519
rect 54 78961 154 78964
rect 49 78861 54 78961
rect 154 78861 158 78961
rect 54 78858 154 78861
rect -413 78450 -368 78474
rect -2581 78428 -368 78450
rect -2584 78371 -368 78428
rect 151965 78179 152120 78181
rect 151960 78019 151963 78179
rect 152123 78019 152126 78179
rect 151965 78017 152120 78019
rect 54 77461 154 77464
rect 49 77361 54 77461
rect 154 77361 158 77461
rect 54 77358 154 77361
rect -441 76839 -396 76974
rect -2567 76794 -396 76839
rect 151965 76679 152120 76681
rect 151960 76519 151963 76679
rect 152123 76519 152126 76679
rect 151965 76517 152120 76519
rect 54 75961 154 75964
rect 49 75861 54 75961
rect 154 75861 158 75961
rect 54 75858 154 75861
rect -2621 75292 -2505 75329
rect -446 75292 -401 75474
rect -2621 75284 -401 75292
rect -2550 75247 -401 75284
rect 151965 75179 152120 75181
rect 151960 75019 151963 75179
rect 152123 75019 152126 75179
rect 151965 75017 152120 75019
rect 54 74461 154 74464
rect 49 74361 54 74461
rect 154 74361 158 74461
rect 54 74358 154 74361
rect -2561 73714 -2516 73777
rect -441 73714 -396 73974
rect -2561 73669 -396 73714
rect 151965 73679 152120 73681
rect 151960 73519 151963 73679
rect 152123 73519 152126 73679
rect 151965 73517 152120 73519
rect 54 72961 154 72964
rect 49 72861 54 72961
rect 154 72861 158 72961
rect 54 72858 154 72861
rect -441 72284 -396 72474
rect -2589 72239 -396 72284
rect -2589 72208 -419 72239
rect 151965 72179 152120 72181
rect 151960 72019 151963 72179
rect 152123 72019 152126 72179
rect 151965 72017 152120 72019
rect 54 71461 154 71464
rect 49 71361 54 71461
rect 154 71361 158 71461
rect 54 71358 154 71361
rect -433 70752 -388 70974
rect -2570 70707 -388 70752
rect -2570 70676 -408 70707
rect 151965 70679 152120 70681
rect 151960 70519 151963 70679
rect 152123 70519 152126 70679
rect 151965 70517 152120 70519
rect 54 69961 154 69964
rect 49 69861 54 69961
rect 154 69861 158 69961
rect 54 69858 154 69861
rect -430 69169 -385 69474
rect 151965 69179 152120 69181
rect -2589 69124 -385 69169
rect 151960 69019 151963 69179
rect 152123 69019 152126 69179
rect 151965 69017 152120 69019
rect 54 68461 154 68464
rect 49 68361 54 68461
rect 154 68361 158 68461
rect 54 68358 154 68361
rect -446 67670 -401 67974
rect 151965 67679 152120 67681
rect -2595 67625 -401 67670
rect -2567 67591 -402 67625
rect 151960 67519 151963 67679
rect 152123 67519 152126 67679
rect 151965 67517 152120 67519
rect 54 66961 154 66964
rect 49 66861 54 66961
rect 154 66861 158 66961
rect 54 66858 154 66861
rect -424 66184 -379 66474
rect -2587 66139 -379 66184
rect 151965 66179 152120 66181
rect -2587 66093 -2542 66139
rect 151960 66019 151963 66179
rect 152123 66019 152126 66179
rect 151965 66017 152120 66019
rect 54 65461 154 65464
rect 49 65361 54 65461
rect 154 65361 158 65461
rect 54 65358 154 65361
rect -440 64542 -395 64974
rect 151965 64679 152120 64681
rect -2593 64468 -395 64542
rect 151960 64519 151963 64679
rect 152123 64519 152126 64679
rect 151965 64517 152120 64519
rect 54 63961 154 63964
rect 49 63861 54 63961
rect 154 63861 158 63961
rect 54 63858 154 63861
rect -426 63042 -381 63474
rect 151965 63179 152120 63181
rect -2599 62969 -381 63042
rect 151960 63019 151963 63179
rect 152123 63019 152126 63179
rect 151965 63017 152120 63019
rect 54 62461 154 62464
rect 49 62361 54 62461
rect 154 62361 158 62461
rect 54 62358 154 62361
rect -446 61488 -401 61974
rect 151965 61679 152120 61681
rect 151960 61519 151963 61679
rect 152123 61519 152126 61679
rect 151965 61517 152120 61519
rect -2570 61395 -401 61488
rect 54 60961 154 60964
rect 49 60861 54 60961
rect 154 60861 158 60961
rect 54 60858 154 60861
rect -2564 60474 -2536 60579
rect -2570 60429 -381 60474
rect -2564 59927 -2536 60429
rect 151965 60179 152120 60181
rect 151960 60019 151963 60179
rect 152123 60019 152126 60179
rect 151965 60017 152120 60019
rect 54 59461 154 59464
rect 49 59361 54 59461
rect 154 59361 158 59461
rect 54 59358 154 59361
rect -2593 58929 -401 58974
rect -2593 58387 -2548 58929
rect 151965 58679 152120 58681
rect 151960 58519 151963 58679
rect 152123 58519 152126 58679
rect 151965 58517 152120 58519
rect 54 57961 154 57964
rect 49 57861 54 57961
rect 154 57861 158 57961
rect 54 57858 154 57861
rect -2579 57429 -307 57474
rect -2579 56825 -2534 57429
rect 151965 57179 152120 57181
rect 151960 57019 151963 57179
rect 152123 57019 152126 57179
rect 151965 57017 152120 57019
rect 54 56461 154 56464
rect 49 56361 54 56461
rect 154 56361 158 56461
rect 54 56358 154 56361
rect -2596 55929 -384 55974
rect -2596 55316 -2551 55929
rect 151965 55679 152120 55681
rect 151960 55519 151963 55679
rect 152123 55519 152126 55679
rect 151965 55517 152120 55519
rect 54 54961 154 54964
rect 49 54861 54 54961
rect 154 54861 158 54961
rect 54 54858 154 54861
rect -2562 54429 -401 54474
rect -2562 53811 -2517 54429
rect 151965 54179 152120 54181
rect 151960 54019 151963 54179
rect 152123 54019 152126 54179
rect 151965 54017 152120 54019
rect 54 53461 154 53464
rect 49 53361 54 53461
rect 154 53361 158 53461
rect 54 53358 154 53361
rect -418 52294 -373 52974
rect 151965 52679 152120 52681
rect 151960 52519 151963 52679
rect 152123 52519 152126 52679
rect 151965 52517 152120 52519
rect -2582 52249 -373 52294
rect -2582 52245 -384 52249
rect 54 51961 154 51964
rect 49 51861 54 51961
rect 154 51861 158 51961
rect 54 51858 154 51861
rect -446 50774 -401 51474
rect 151965 51179 152120 51181
rect 151960 51019 151963 51179
rect 152123 51019 152126 51179
rect 151965 51017 152120 51019
rect -2587 50729 -401 50774
rect -446 50629 -401 50729
rect 54 50461 154 50464
rect 49 50361 54 50461
rect 154 50361 158 50461
rect 54 50358 154 50361
rect -446 49214 -401 49974
rect 151965 49679 152120 49681
rect 151960 49519 151963 49679
rect 152123 49519 152126 49679
rect 151965 49517 152120 49519
rect -2604 49169 -401 49214
rect -446 49038 -401 49169
rect 54 48961 154 48964
rect 49 48861 54 48961
rect 154 48861 158 48961
rect 54 48858 154 48861
rect -440 47698 -395 48474
rect 151965 48179 152120 48181
rect 151960 48019 151963 48179
rect 152123 48019 152126 48179
rect 151965 48017 152120 48019
rect -2590 47653 -395 47698
rect -440 47504 -395 47653
rect 54 47461 154 47464
rect 49 47361 54 47461
rect 154 47361 158 47461
rect 54 47358 154 47361
rect -435 46158 -390 46974
rect 151965 46679 152120 46681
rect 151960 46519 151963 46679
rect 152123 46519 152126 46679
rect 151965 46517 152120 46519
rect -2616 46113 -390 46158
rect -435 45956 -390 46113
rect 54 45961 154 45964
rect 49 45861 54 45961
rect 154 45861 158 45961
rect 54 45858 154 45861
rect -426 44604 -381 45474
rect 151965 45179 152120 45181
rect 151960 45019 151963 45179
rect 152123 45019 152126 45179
rect 151965 45017 152120 45019
rect -2596 44559 -381 44604
rect -426 44508 -381 44559
rect 54 44461 154 44464
rect 49 44361 54 44461
rect 154 44361 158 44461
rect 54 44358 154 44361
rect -418 43099 -373 43974
rect 151965 43679 152120 43681
rect 151960 43519 151963 43679
rect 152123 43519 152126 43679
rect 151965 43517 152120 43519
rect -2564 43054 -373 43099
rect -418 42988 -373 43054
rect 54 42961 154 42964
rect 49 42861 54 42961
rect 154 42861 158 42961
rect 54 42858 154 42861
rect -398 41576 -353 42474
rect 151965 42179 152120 42181
rect 151960 42019 151963 42179
rect 152123 42019 152126 42179
rect 151965 42017 152120 42019
rect -2610 41531 -353 41576
rect -398 41360 -353 41531
rect 54 41461 154 41464
rect 49 41361 54 41461
rect 154 41361 158 41461
rect 54 41358 154 41361
rect -440 40011 -395 40974
rect 151965 40679 152120 40681
rect 151960 40519 151963 40679
rect 152123 40519 152126 40679
rect 151965 40517 152120 40519
rect -2601 39966 -395 40011
rect -440 39763 -395 39966
rect 54 39961 154 39964
rect 49 39861 54 39961
rect 154 39861 158 39961
rect 54 39858 154 39861
rect -429 38474 -384 39474
rect 151965 39179 152120 39181
rect 151960 39019 151963 39179
rect 152123 39019 152126 39179
rect 151965 39017 152120 39019
rect -2604 38429 -384 38474
rect 54 38461 154 38464
rect -429 38195 -384 38429
rect 49 38361 54 38461
rect 154 38361 158 38461
rect 54 38358 154 38361
rect -2582 36886 -2537 37029
rect -395 36886 -350 37974
rect 151965 37679 152120 37681
rect 151960 37519 151963 37679
rect 152123 37519 152126 37679
rect 151965 37517 152120 37519
rect 54 36961 154 36964
rect -2582 36841 -350 36886
rect 49 36861 54 36961
rect 154 36861 158 36961
rect 54 36858 154 36861
rect -395 36738 -350 36841
rect -415 35398 -370 36474
rect 151965 36179 152120 36181
rect 151960 36019 151963 36179
rect 152123 36019 152126 36179
rect 151965 36017 152120 36019
rect 54 35461 154 35464
rect -2576 35353 -370 35398
rect 49 35361 54 35461
rect 154 35361 158 35461
rect 54 35358 154 35361
rect -415 35290 -370 35353
rect -2584 33827 -2539 33887
rect -446 33827 -401 34974
rect 151965 34679 152120 34681
rect 151960 34519 151963 34679
rect 152123 34519 152126 34679
rect 151965 34517 152120 34519
rect 54 33961 154 33964
rect 49 33861 54 33961
rect 154 33861 158 33961
rect 54 33858 154 33861
rect -2584 33782 -401 33827
rect -446 33685 -401 33782
rect -304 32309 -276 33462
rect 151965 33179 152120 33181
rect 151960 33019 151963 33179
rect 152123 33019 152126 33179
rect 151965 33017 152120 33019
rect 54 32461 154 32464
rect 49 32361 54 32461
rect 154 32361 158 32461
rect 54 32358 154 32361
rect -2613 32281 -276 32309
rect -2604 31929 -321 31974
rect -2604 30677 -2559 31929
rect 151965 31679 152120 31681
rect 151960 31519 151963 31679
rect 152123 31519 152126 31679
rect 151965 31517 152120 31519
rect 54 30961 154 30964
rect 49 30861 54 30961
rect 154 30861 158 30961
rect 54 30858 154 30861
rect -2621 30429 -350 30474
rect -2621 29189 -2576 30429
rect 151965 30179 152120 30181
rect 151960 30019 151963 30179
rect 152123 30019 152126 30179
rect 151965 30017 152120 30019
rect 54 29461 154 29464
rect 49 29361 54 29461
rect 154 29361 158 29461
rect 54 29358 154 29361
rect -2607 28929 -387 28974
rect -2607 27612 -2562 28929
rect 151965 28679 152120 28681
rect 151960 28519 151963 28679
rect 152123 28519 152126 28679
rect 151965 28517 152120 28519
rect 54 27961 154 27964
rect 49 27861 54 27961
rect 154 27861 158 27961
rect 54 27858 154 27861
rect -2621 27429 -387 27474
rect -2621 26158 -2576 27429
rect 151965 27179 152120 27181
rect 151960 27019 151963 27179
rect 152123 27019 152126 27179
rect 151965 27017 152120 27019
rect 54 26461 154 26464
rect 49 26361 54 26461
rect 154 26361 158 26461
rect 54 26358 154 26361
rect -161 24673 -133 26089
rect 151965 25679 152120 25681
rect 151960 25519 151963 25679
rect 152123 25519 152126 25679
rect 151965 25517 152120 25519
rect 54 24961 154 24964
rect 49 24861 54 24961
rect 154 24861 158 24961
rect 54 24858 154 24861
rect -2573 24645 -133 24673
rect -2613 24429 -244 24474
rect -2613 22985 -2568 24429
rect 151965 24179 152120 24181
rect 151960 24019 151963 24179
rect 152123 24019 152126 24179
rect 151965 24017 152120 24019
rect 54 23461 154 23464
rect 49 23361 54 23461
rect 154 23361 158 23461
rect 54 23358 154 23361
rect -1770 22929 -401 22974
rect -1770 21591 -1725 22929
rect 151965 22679 152120 22681
rect 151960 22519 151963 22679
rect 152123 22519 152126 22679
rect 151965 22517 152120 22519
rect 54 21961 154 21964
rect 49 21861 54 21961
rect 154 21861 158 21961
rect 54 21858 154 21861
rect -2594 21563 -1671 21591
rect -1770 21245 -1725 21563
rect -1180 21474 -1152 21595
rect -1229 21429 -401 21474
rect -1180 20027 -1152 21429
rect 151965 21179 152120 21181
rect 151960 21019 151963 21179
rect 152123 21019 152126 21179
rect 151965 21017 152120 21019
rect 54 20461 154 20464
rect 49 20361 54 20461
rect 154 20361 158 20461
rect 54 20358 154 20361
rect -2628 19999 -1152 20027
rect -375 19221 -330 19974
rect 151965 19679 152120 19681
rect 151960 19519 151963 19679
rect 152123 19519 152126 19679
rect 151965 19517 152120 19519
rect -995 19193 -248 19221
rect -995 18509 -967 19193
rect -375 19140 -330 19193
rect 54 18961 154 18964
rect 49 18861 54 18961
rect 154 18861 158 18961
rect 54 18858 154 18861
rect -2565 18481 -967 18509
rect -231 17782 -186 18474
rect 151965 18179 152120 18181
rect 151960 18019 151963 18179
rect 152123 18019 152126 18179
rect 151965 18017 152120 18019
rect -1217 17754 -186 17782
rect -1217 16991 -1189 17754
rect -231 17627 -186 17754
rect 54 17461 154 17464
rect 49 17361 54 17461
rect 154 17361 158 17461
rect 54 17358 154 17361
rect -2572 16963 -1189 16991
rect -386 16425 -358 17279
rect 151965 16679 152120 16681
rect 151960 16519 151963 16679
rect 152123 16519 152126 16679
rect 151965 16517 152120 16519
rect -1649 16397 -358 16425
rect -1649 15427 -1621 16397
rect 54 15961 154 15964
rect 49 15861 54 15961
rect 154 15861 158 15961
rect 54 15858 154 15861
rect -2587 15399 -1621 15427
rect -360 14870 -315 15474
rect 151965 15179 152120 15181
rect 151960 15019 151963 15179
rect 152123 15019 152126 15179
rect 151965 15017 152120 15019
rect -1452 14842 -292 14870
rect -1452 13909 -1424 14842
rect -360 14692 -292 14842
rect -360 14630 -315 14692
rect 54 14461 154 14464
rect 49 14361 54 14461
rect 154 14361 158 14461
rect 54 14358 154 14361
rect -2587 13881 -1424 13909
rect -378 13450 -333 13974
rect 151965 13679 152120 13681
rect 151960 13519 151963 13679
rect 152123 13519 152126 13679
rect 151965 13517 152120 13519
rect -1296 13422 -314 13450
rect -1296 12391 -1268 13422
rect -378 13295 -333 13422
rect 54 12961 154 12964
rect 49 12861 54 12961
rect 154 12861 158 12961
rect 54 12858 154 12861
rect -2594 12363 -1268 12391
rect -382 11955 -337 12474
rect 151965 12179 152120 12181
rect 151960 12019 151963 12179
rect 152123 12019 152126 12179
rect 151965 12017 152120 12019
rect -2622 11927 -229 11955
rect -2622 10799 -2594 11927
rect -382 11759 -337 11927
rect 54 11461 154 11464
rect 49 11361 54 11461
rect 154 11361 158 11461
rect 54 11358 154 11361
rect -2008 10929 -368 10974
rect -2008 9309 -1963 10929
rect 151965 10679 152120 10681
rect 151960 10519 151963 10679
rect 152123 10519 152126 10679
rect 151965 10517 152120 10519
rect 151424 9736 151514 9739
rect 151424 9646 153682 9736
rect 151424 9639 151514 9646
rect 19156 9607 19281 9613
rect 9925 9594 10050 9601
rect 9925 9489 9937 9594
rect 10042 9489 10050 9594
rect 14542 9531 14652 9535
rect 6895 9465 7020 9475
rect 9925 9472 10050 9489
rect 12954 9503 13113 9514
rect 6825 9462 7020 9465
rect 3735 9443 3860 9455
rect 2658 9392 2783 9405
rect 2259 9390 2783 9392
rect 1832 9380 1992 9383
rect -2590 9255 -1902 9309
rect -2590 9248 -1963 9255
rect 1158 9220 1283 9233
rect 1830 9222 1832 9377
rect 1992 9222 1994 9377
rect 2259 9285 2666 9390
rect 2771 9285 2783 9390
rect 3735 9338 3743 9443
rect 3848 9338 3860 9443
rect 3735 9326 3860 9338
rect 5346 9415 5471 9429
rect 2259 9282 2783 9285
rect 749 9217 1283 9220
rect 749 9112 1166 9217
rect 1271 9112 1283 9217
rect 1832 9217 1992 9220
rect 749 9110 1283 9112
rect -3099 8973 -2999 8978
rect -3099 8869 -2999 8873
rect 749 8278 859 9110
rect 1158 9104 1283 9110
rect 2259 8215 2369 9282
rect 2658 9276 2783 9282
rect 3741 8228 3851 9326
rect 5346 9310 5358 9415
rect 5463 9310 5471 9415
rect 5346 9300 5471 9310
rect 6825 9357 6903 9462
rect 7008 9357 7020 9462
rect 6825 9346 7020 9357
rect 8450 9406 8575 9412
rect 5355 8263 5465 9300
rect 6825 8225 6935 9346
rect 8450 9301 8458 9406
rect 8563 9301 8575 9406
rect 9044 9380 9204 9383
rect 8450 9283 8575 9301
rect 8455 8347 8565 9283
rect 9042 9222 9044 9377
rect 9204 9222 9206 9377
rect 9044 9217 9204 9220
rect 8373 8237 8565 8347
rect 9934 8241 10044 9472
rect 12954 9398 12974 9503
rect 13079 9398 13113 9503
rect 14537 9421 14542 9526
rect 14652 9421 14656 9526
rect 17649 9525 17792 9533
rect 16166 9493 16271 9495
rect 16062 9491 16274 9493
rect 12954 9381 13113 9398
rect 11436 9327 11594 9336
rect 11436 9222 11451 9327
rect 11556 9222 11594 9327
rect 11436 9203 11594 9222
rect 11448 8228 11558 9203
rect 12971 8225 13081 9381
rect 14542 8241 14652 9421
rect 16062 9386 16166 9491
rect 16271 9386 16274 9491
rect 17649 9420 17666 9525
rect 17771 9420 17792 9525
rect 19156 9502 19166 9607
rect 19271 9502 19281 9607
rect 28297 9579 28422 9589
rect 19156 9484 19281 9502
rect 23659 9563 23784 9572
rect 17649 9414 17792 9420
rect 16062 9383 16274 9386
rect 16062 9381 16271 9383
rect 16062 8263 16172 9381
rect 16457 9380 16617 9383
rect 16455 9222 16457 9377
rect 16617 9222 16619 9377
rect 16457 9217 16617 9220
rect 17664 8624 17774 9414
rect 17598 8514 17774 8624
rect 17598 8241 17708 8514
rect 19164 8256 19274 9484
rect 22160 9459 22285 9468
rect 20659 9434 20784 9446
rect 20659 9329 20666 9434
rect 20771 9329 20784 9434
rect 22160 9354 22166 9459
rect 22271 9354 22285 9459
rect 23659 9458 23666 9563
rect 23771 9458 23784 9563
rect 26760 9519 26885 9532
rect 23659 9443 23784 9458
rect 25250 9503 25375 9511
rect 22160 9339 22285 9354
rect 20659 9317 20784 9329
rect 20664 8228 20774 9317
rect 22164 8212 22274 9339
rect 23664 8816 23774 9443
rect 25250 9398 25260 9503
rect 25365 9398 25375 9503
rect 26760 9414 26771 9519
rect 26876 9414 26885 9519
rect 28297 9474 28310 9579
rect 28415 9474 28422 9579
rect 87183 9565 87293 9568
rect 37526 9513 37673 9522
rect 54450 9514 54560 9516
rect 34277 9476 34382 9478
rect 28297 9460 28422 9474
rect 34275 9474 34629 9476
rect 26760 9403 26885 9414
rect 25250 9382 25375 9398
rect 23664 8706 23867 8816
rect 23757 8253 23867 8706
rect 25258 8237 25368 9382
rect 26768 8905 26878 9403
rect 26768 8795 26944 8905
rect 26834 8253 26944 8795
rect 28307 8222 28417 9460
rect 29804 9433 29929 9443
rect 32868 9438 33005 9446
rect 29804 9431 30000 9433
rect 29804 9326 29817 9431
rect 29922 9326 30000 9431
rect 29804 9314 30000 9326
rect 29890 8247 30000 9314
rect 31310 9395 31435 9401
rect 31310 9393 31498 9395
rect 31310 9288 31318 9393
rect 31423 9288 31498 9393
rect 32128 9380 32288 9383
rect 31310 9272 31498 9288
rect 31388 8234 31498 9272
rect 32126 9222 32128 9377
rect 32288 9222 32290 9377
rect 32868 9333 32873 9438
rect 32978 9333 33005 9438
rect 34275 9369 34277 9474
rect 34382 9369 34629 9474
rect 37526 9408 37541 9513
rect 37646 9408 37673 9513
rect 48226 9435 48336 9438
rect 45206 9416 45316 9419
rect 37526 9391 37673 9408
rect 34275 9366 34629 9369
rect 34277 9364 34382 9366
rect 32868 9305 33005 9333
rect 32128 9217 32288 9220
rect 32973 8249 33001 9305
rect 34519 8253 34629 9366
rect 35964 9260 36074 9262
rect 35962 9155 35966 9260
rect 36071 9155 36076 9260
rect 35964 8503 36074 9155
rect 35964 8393 36139 8503
rect 36029 8253 36139 8393
rect 37539 8208 37649 9391
rect 40595 9353 40705 9355
rect 40593 9248 40597 9353
rect 40702 9248 40707 9353
rect 45204 9311 45208 9416
rect 45313 9311 45318 9416
rect 46778 9394 46888 9397
rect 39051 9041 39156 9043
rect 39049 9038 39159 9041
rect 39049 8933 39051 9038
rect 39156 8933 39159 9038
rect 39049 8577 39159 8933
rect 39049 8467 39226 8577
rect 39116 8246 39226 8467
rect 40595 8239 40705 9248
rect 43667 9155 43777 9157
rect 43665 9050 43670 9155
rect 43775 9050 43779 9155
rect 42137 8990 42247 8992
rect 42135 8885 42139 8990
rect 42244 8885 42249 8990
rect 42137 8246 42247 8885
rect 43667 8190 43777 9050
rect 45206 8220 45316 9311
rect 46776 9289 46780 9394
rect 46885 9289 46890 9394
rect 48224 9330 48229 9435
rect 48334 9330 48338 9435
rect 54448 9409 54453 9514
rect 54558 9409 54562 9514
rect 78921 9496 79031 9499
rect 57476 9490 57586 9492
rect 55974 9465 56084 9468
rect 52837 9375 52947 9378
rect 51355 9368 51465 9370
rect 46778 8224 46888 9289
rect 48226 8513 48336 9330
rect 51353 9263 51358 9368
rect 51463 9263 51467 9368
rect 52835 9270 52840 9375
rect 52945 9270 52949 9375
rect 49801 9251 49906 9253
rect 49798 9248 49908 9251
rect 49798 9143 49801 9248
rect 49906 9143 49908 9248
rect 48226 8403 48407 8513
rect 48297 8239 48407 8403
rect 49798 8257 49908 9143
rect 51355 8205 51465 9263
rect 52837 8498 52947 9270
rect 52837 8388 53007 8498
rect 52897 8231 53007 8388
rect 54450 8227 54560 9409
rect 55972 9360 55976 9465
rect 56081 9360 56086 9465
rect 57474 9385 57479 9490
rect 57584 9385 57588 9490
rect 58980 9486 59101 9496
rect 55974 8257 56084 9360
rect 57476 8226 57586 9385
rect 58980 9381 58986 9486
rect 59091 9381 59101 9486
rect 63620 9469 63730 9471
rect 58980 9373 59101 9381
rect 60564 9430 60691 9439
rect 58984 8952 59094 9373
rect 60564 9325 60577 9430
rect 60682 9325 60691 9430
rect 62059 9426 62169 9430
rect 62057 9421 62059 9423
rect 60839 9380 60999 9383
rect 60564 9307 60691 9325
rect 58984 8842 59184 8952
rect 59074 8241 59184 8842
rect 60575 8230 60685 9307
rect 60837 9222 60839 9377
rect 60999 9222 61001 9377
rect 62054 9316 62059 9421
rect 62169 9421 62171 9423
rect 62169 9316 62173 9421
rect 63618 9364 63623 9469
rect 63728 9364 63732 9469
rect 66706 9433 66816 9438
rect 66704 9428 66706 9431
rect 65125 9404 65235 9407
rect 60839 9217 60999 9220
rect 62059 8276 62169 9316
rect 63620 8230 63730 9364
rect 65123 9299 65127 9404
rect 65232 9299 65237 9404
rect 66701 9323 66706 9428
rect 66816 9428 66818 9431
rect 66816 9323 66820 9428
rect 77396 9427 77506 9429
rect 72789 9419 72899 9422
rect 74377 9419 74487 9422
rect 71299 9332 71409 9334
rect 65125 8238 65235 9299
rect 66706 8230 66816 9323
rect 69776 9298 69886 9300
rect 69774 9193 69778 9298
rect 69883 9193 69888 9298
rect 71297 9227 71302 9332
rect 71407 9227 71411 9332
rect 72787 9314 72791 9419
rect 72896 9314 72901 9419
rect 74375 9314 74379 9419
rect 74484 9314 74489 9419
rect 75886 9385 75996 9387
rect 68233 9118 68343 9121
rect 68231 9013 68236 9118
rect 68341 9013 68345 9118
rect 68233 8200 68343 9013
rect 69776 8242 69886 9193
rect 71299 8234 71409 9227
rect 72789 8473 72899 9314
rect 72789 8363 72959 8473
rect 72849 8226 72959 8363
rect 74377 8203 74487 9314
rect 75884 9280 75888 9385
rect 75993 9280 75998 9385
rect 77394 9322 77398 9427
rect 77503 9322 77508 9427
rect 78919 9391 78924 9496
rect 79029 9391 79033 9496
rect 87181 9460 87185 9565
rect 87290 9460 87295 9565
rect 152692 9547 152802 9550
rect 145166 9478 145271 9480
rect 145164 9475 146809 9478
rect 114829 9467 114939 9470
rect 75886 8186 75996 9280
rect 77396 8807 77506 9322
rect 77396 8697 77583 8807
rect 77473 8232 77583 8697
rect 78921 8519 79031 9391
rect 83774 9380 83934 9383
rect 80443 9377 80553 9379
rect 80441 9272 80445 9377
rect 80550 9272 80555 9377
rect 80443 8596 80553 9272
rect 81621 9230 81726 9232
rect 81619 9227 82159 9230
rect 81619 9122 81621 9227
rect 81726 9122 82159 9227
rect 83772 9222 83774 9377
rect 83934 9222 83936 9377
rect 86533 9242 86668 9267
rect 83774 9217 83934 9220
rect 81619 9120 82159 9122
rect 81621 9118 81726 9120
rect 82049 8844 82159 9120
rect 86533 9137 86543 9242
rect 86648 9137 86668 9242
rect 86533 9119 86668 9137
rect 82966 9087 83071 9089
rect 82964 9085 83661 9087
rect 82964 8980 82966 9085
rect 83071 8980 83661 9085
rect 82964 8977 83661 8980
rect 82966 8975 83071 8977
rect 82026 8666 82159 8844
rect 78921 8409 79112 8519
rect 80443 8486 80622 8596
rect 79002 8247 79112 8409
rect 80512 8270 80622 8486
rect 82026 8220 82136 8666
rect 83551 8220 83661 8977
rect 86541 8803 86651 9119
rect 84434 8711 84539 8713
rect 84431 8708 85241 8711
rect 84431 8603 84434 8708
rect 84539 8603 85241 8708
rect 86541 8693 86755 8803
rect 84431 8601 85241 8603
rect 84434 8599 84539 8601
rect 85131 8251 85241 8601
rect 86645 8232 86755 8693
rect 87183 8780 87293 9460
rect 88155 9406 88282 9411
rect 88155 9404 89606 9406
rect 88155 9299 88166 9404
rect 88271 9299 89606 9404
rect 90274 9380 90434 9383
rect 94774 9380 94934 9383
rect 99274 9380 99434 9383
rect 102274 9380 102434 9383
rect 105774 9380 105934 9383
rect 111774 9380 111934 9383
rect 88155 9296 89606 9299
rect 88155 9289 88282 9296
rect 87183 8670 88334 8780
rect 88224 8228 88334 8670
rect 89496 8645 89606 9296
rect 90272 9222 90274 9377
rect 90434 9222 90436 9377
rect 94772 9222 94774 9377
rect 94934 9222 94936 9377
rect 99272 9222 99274 9377
rect 99434 9222 99436 9377
rect 102272 9222 102274 9377
rect 102434 9222 102436 9377
rect 103166 9228 103271 9230
rect 103164 9225 104350 9228
rect 90274 9217 90434 9220
rect 94774 9217 94934 9220
rect 99274 9217 99434 9220
rect 102274 9217 102434 9220
rect 103164 9120 103166 9225
rect 103271 9120 104350 9225
rect 105772 9222 105774 9377
rect 105934 9222 105936 9377
rect 107666 9282 107771 9284
rect 107664 9279 109808 9282
rect 105774 9217 105934 9220
rect 107664 9174 107666 9279
rect 107771 9174 109808 9279
rect 111772 9222 111774 9377
rect 111934 9222 111936 9377
rect 114827 9362 114831 9467
rect 114936 9362 114941 9467
rect 116274 9380 116434 9383
rect 119274 9380 119434 9383
rect 125274 9380 125434 9383
rect 131974 9380 132134 9383
rect 134974 9380 135134 9383
rect 136474 9380 136634 9383
rect 137974 9380 138134 9383
rect 140974 9380 141134 9383
rect 142974 9380 143134 9383
rect 111774 9217 111934 9220
rect 113597 9212 113707 9214
rect 107664 9172 109808 9174
rect 107666 9170 107771 9172
rect 103164 9118 104350 9120
rect 103166 9116 103271 9118
rect 92666 9018 92771 9020
rect 92664 9016 94063 9018
rect 91236 8927 91346 8930
rect 91234 8822 91239 8927
rect 91344 8822 91348 8927
rect 92664 8911 92666 9016
rect 92771 8911 94063 9016
rect 100457 8976 100567 8978
rect 98396 8962 98506 8965
rect 92664 8908 94063 8911
rect 92666 8906 92771 8908
rect 89496 8535 89852 8645
rect 89742 8247 89852 8535
rect 91236 8240 91346 8822
rect 92007 8576 92112 8578
rect 92005 8574 92937 8576
rect 92005 8469 92007 8574
rect 92112 8469 92937 8574
rect 92005 8466 92937 8469
rect 92007 8464 92112 8466
rect 92827 8228 92937 8466
rect 93953 8442 94063 8908
rect 98394 8857 98399 8962
rect 98504 8857 98508 8962
rect 100455 8871 100460 8976
rect 100565 8871 100569 8976
rect 103499 8873 103609 8876
rect 94166 8830 94271 8832
rect 94164 8827 95938 8830
rect 94164 8722 94166 8827
rect 94271 8722 95938 8827
rect 94164 8720 95938 8722
rect 94166 8718 94271 8720
rect 93953 8332 94420 8442
rect 94310 8224 94420 8332
rect 95828 8243 95938 8720
rect 96735 8510 96840 8512
rect 98396 8510 98506 8857
rect 96732 8507 97525 8510
rect 96732 8402 96735 8507
rect 96840 8402 97525 8507
rect 96732 8400 97525 8402
rect 98396 8400 99068 8510
rect 96735 8398 96840 8400
rect 97415 8226 97525 8400
rect 98958 8190 99068 8400
rect 100457 8235 100567 8871
rect 103497 8768 103502 8873
rect 103607 8768 103611 8873
rect 101004 8447 101109 8449
rect 101001 8445 102128 8447
rect 101001 8340 101004 8445
rect 101109 8340 102128 8445
rect 101001 8337 102128 8340
rect 101004 8335 101109 8337
rect 102018 8257 102128 8337
rect 103499 8261 103609 8768
rect 104240 8545 104350 9118
rect 106577 9047 106687 9049
rect 106575 8942 106580 9047
rect 106685 8942 106689 9047
rect 104240 8435 105215 8545
rect 105105 8253 105215 8435
rect 106577 8217 106687 8942
rect 106954 8635 107059 8637
rect 106952 8632 108248 8635
rect 106952 8527 106954 8632
rect 107059 8527 108248 8632
rect 106952 8525 108248 8527
rect 106954 8523 107059 8525
rect 108138 8186 108248 8525
rect 109698 8217 109808 9172
rect 113595 9107 113599 9212
rect 113704 9107 113709 9212
rect 110666 8856 110771 8858
rect 110664 8853 112860 8856
rect 110664 8748 110666 8853
rect 110771 8748 112860 8853
rect 110664 8746 112860 8748
rect 110666 8744 110771 8746
rect 110346 8614 110451 8616
rect 110344 8612 111341 8614
rect 110344 8507 110346 8612
rect 110451 8507 111341 8612
rect 110344 8504 111341 8507
rect 110346 8502 110451 8504
rect 111231 8213 111341 8504
rect 112750 8249 112860 8746
rect 113597 8762 113707 9107
rect 113597 8652 114419 8762
rect 114309 8240 114419 8652
rect 114829 8717 114939 9362
rect 116272 9222 116274 9377
rect 116434 9222 116436 9377
rect 116666 9345 116771 9347
rect 116664 9342 118801 9345
rect 116664 9237 116666 9342
rect 116771 9340 118801 9342
rect 116771 9237 118974 9340
rect 116664 9235 118974 9237
rect 116666 9233 116771 9235
rect 118678 9230 118974 9235
rect 116274 9217 116434 9220
rect 117325 9149 117520 9152
rect 117323 9044 117327 9149
rect 117432 9044 117520 9149
rect 117325 9042 117520 9044
rect 114829 8607 115938 8717
rect 115828 8271 115938 8607
rect 117410 8253 117520 9042
rect 118864 8980 118974 9230
rect 119272 9222 119274 9377
rect 119434 9222 119436 9377
rect 121166 9285 121271 9287
rect 121164 9283 122544 9285
rect 120836 9265 120946 9267
rect 119274 9217 119434 9220
rect 120834 9160 120838 9265
rect 120943 9160 120948 9265
rect 121164 9178 121166 9283
rect 121271 9178 122544 9283
rect 125272 9222 125274 9377
rect 125434 9222 125436 9377
rect 127166 9350 127271 9352
rect 127164 9348 128768 9350
rect 126962 9252 127072 9255
rect 125274 9217 125434 9220
rect 121164 9175 122544 9178
rect 121166 9173 121271 9175
rect 120458 9005 120568 9008
rect 118853 8889 118974 8980
rect 120456 8900 120460 9005
rect 120565 8900 120570 9005
rect 118853 8213 118963 8889
rect 120458 8242 120568 8900
rect 120836 8607 120946 9160
rect 120836 8497 122075 8607
rect 121965 8160 122075 8497
rect 122434 8493 122544 9175
rect 126960 9147 126965 9252
rect 127070 9147 127074 9252
rect 127164 9243 127166 9348
rect 127271 9243 128768 9348
rect 127164 9240 128768 9243
rect 127166 9238 127271 9240
rect 124822 8930 124962 8941
rect 124822 8928 126673 8930
rect 124822 8823 124836 8928
rect 124941 8823 126673 8928
rect 124822 8820 126673 8823
rect 124822 8811 124962 8820
rect 124358 8539 124463 8541
rect 124355 8536 125134 8539
rect 122434 8383 123636 8493
rect 124355 8431 124358 8536
rect 124463 8431 125134 8536
rect 124355 8429 125134 8431
rect 124358 8427 124463 8429
rect 123526 8260 123636 8383
rect 125024 8210 125134 8429
rect 126563 8260 126673 8820
rect 126962 8677 127072 9147
rect 128658 8679 128768 9240
rect 131972 9222 131974 9377
rect 132134 9222 132136 9377
rect 134516 9278 134626 9280
rect 131974 9217 132134 9220
rect 134514 9173 134518 9278
rect 134623 9173 134628 9278
rect 134972 9222 134974 9377
rect 135134 9222 135136 9377
rect 136472 9222 136474 9377
rect 136634 9222 136636 9377
rect 137972 9222 137974 9377
rect 138134 9222 138136 9377
rect 139838 9347 139948 9349
rect 139836 9242 139840 9347
rect 139945 9242 139950 9347
rect 134974 9217 135134 9220
rect 136474 9217 136634 9220
rect 137974 9217 138134 9220
rect 130524 9063 130629 9065
rect 130522 9060 132824 9063
rect 130522 8955 130524 9060
rect 130629 8955 132824 9060
rect 132937 8982 133042 8984
rect 130522 8953 132824 8955
rect 130524 8951 130629 8953
rect 129683 8679 129793 8693
rect 126962 8567 128208 8677
rect 128658 8569 129804 8679
rect 130029 8623 130134 8625
rect 130026 8621 131303 8623
rect 128098 8219 128208 8567
rect 129683 8253 129793 8569
rect 130026 8516 130029 8621
rect 130134 8516 131303 8621
rect 130026 8513 131303 8516
rect 130029 8511 130134 8513
rect 131193 8240 131303 8513
rect 132714 8219 132824 8953
rect 132935 8979 133689 8982
rect 132935 8874 132937 8979
rect 133042 8874 133689 8979
rect 132935 8872 133689 8874
rect 132937 8870 133042 8872
rect 133579 8685 133689 8872
rect 133579 8575 134376 8685
rect 133579 8574 133689 8575
rect 134266 8194 134376 8575
rect 134516 8545 134626 9173
rect 134666 9134 134771 9136
rect 134664 9132 137406 9134
rect 134664 9027 134666 9132
rect 134771 9027 137406 9132
rect 139439 9101 139549 9103
rect 134664 9024 137406 9027
rect 134666 9022 134771 9024
rect 134516 8435 135905 8545
rect 135795 8203 135905 8435
rect 137296 8251 137406 9024
rect 139437 8996 139441 9101
rect 139546 8996 139551 9101
rect 138846 8789 138956 8791
rect 138844 8684 138849 8789
rect 138954 8684 138958 8789
rect 138846 8241 138956 8684
rect 139439 8573 139549 8996
rect 139838 8958 139948 9242
rect 140972 9222 140974 9377
rect 141134 9222 141136 9377
rect 142972 9222 142974 9377
rect 143134 9222 143136 9377
rect 145164 9370 145166 9475
rect 145271 9370 146809 9475
rect 152690 9442 152695 9547
rect 152800 9442 152804 9547
rect 146974 9380 147134 9383
rect 148474 9380 148634 9383
rect 149974 9380 150134 9383
rect 151474 9380 151634 9383
rect 145164 9368 146809 9370
rect 145166 9366 145271 9368
rect 140974 9217 141134 9220
rect 142974 9217 143134 9220
rect 146203 9111 146313 9114
rect 142166 9069 142271 9071
rect 142164 9066 143911 9069
rect 142164 8961 142166 9066
rect 142271 8961 143911 9066
rect 146201 9006 146206 9111
rect 146311 9006 146315 9111
rect 142164 8959 143911 8961
rect 139838 8848 142056 8958
rect 142166 8957 142271 8959
rect 139439 8463 140485 8573
rect 140375 8182 140485 8463
rect 141946 8227 142056 8848
rect 143464 8754 143574 8756
rect 143462 8649 143467 8754
rect 143572 8649 143576 8754
rect 143464 8223 143574 8649
rect 143801 8490 143911 8959
rect 143801 8380 145093 8490
rect 144983 8244 145093 8380
rect 146203 8462 146313 9006
rect 146699 8677 146809 9368
rect 146972 9222 146974 9377
rect 147134 9222 147136 9377
rect 148472 9222 148474 9377
rect 148634 9222 148636 9377
rect 149972 9222 149974 9377
rect 150134 9222 150136 9377
rect 151472 9222 151474 9377
rect 151634 9222 151636 9377
rect 146974 9217 147134 9220
rect 148474 9217 148634 9220
rect 149974 9217 150134 9220
rect 151474 9217 151634 9220
rect 149629 8859 149739 8862
rect 149627 8754 149631 8859
rect 149736 8754 149741 8859
rect 146699 8567 148203 8677
rect 146203 8352 146653 8462
rect 146543 8223 146653 8352
rect 148093 8230 148203 8567
rect 149629 8445 149739 8754
rect 150128 8553 150233 8555
rect 149573 8335 149739 8445
rect 150125 8550 151250 8553
rect 150125 8445 150128 8550
rect 150233 8445 151250 8550
rect 150125 8443 151250 8445
rect 150128 8441 150233 8443
rect 149573 8199 149683 8335
rect 151140 8255 151250 8443
rect 152692 8252 152802 9442
rect 151473 8208 151634 8212
rect 151470 8047 151473 8208
rect 151634 8047 151637 8208
rect 151473 8042 151634 8047
rect 9044 7856 9204 7860
rect 1832 7847 1992 7851
rect 54 7794 154 7798
rect 51 7694 54 7794
rect 154 7694 157 7794
rect 54 7689 154 7694
rect 1829 7687 1832 7847
rect 1992 7687 1995 7847
rect 9041 7696 9044 7856
rect 9204 7696 9207 7856
rect 60839 7855 60999 7859
rect 83774 7856 83934 7860
rect 90274 7856 90434 7860
rect 94774 7856 94934 7860
rect 99274 7856 99434 7860
rect 102274 7856 102434 7860
rect 105774 7856 105934 7860
rect 111774 7856 111934 7860
rect 116274 7856 116434 7860
rect 119274 7856 119434 7860
rect 125274 7856 125434 7860
rect 131974 7856 132134 7860
rect 134974 7856 135134 7860
rect 136474 7856 136634 7860
rect 137974 7856 138134 7860
rect 140974 7856 141134 7860
rect 142974 7856 143134 7860
rect 146974 7856 147134 7860
rect 148474 7856 148634 7860
rect 149974 7856 150134 7860
rect 151474 7856 151634 7860
rect 16457 7844 16617 7848
rect 32128 7848 32288 7852
rect 9044 7691 9204 7696
rect 1832 7682 1992 7687
rect 16454 7684 16457 7844
rect 16617 7684 16620 7844
rect 32125 7688 32128 7848
rect 32288 7688 32291 7848
rect 60836 7695 60839 7855
rect 60999 7695 61002 7855
rect 83771 7696 83774 7856
rect 83934 7696 83937 7856
rect 90271 7696 90274 7856
rect 90434 7696 90437 7856
rect 94771 7696 94774 7856
rect 94934 7696 94937 7856
rect 99271 7696 99274 7856
rect 99434 7696 99437 7856
rect 102271 7696 102274 7856
rect 102434 7696 102437 7856
rect 105771 7696 105774 7856
rect 105934 7696 105937 7856
rect 111771 7696 111774 7856
rect 111934 7696 111937 7856
rect 116271 7696 116274 7856
rect 116434 7696 116437 7856
rect 119271 7696 119274 7856
rect 119434 7696 119437 7856
rect 125271 7696 125274 7856
rect 125434 7696 125437 7856
rect 131971 7696 131974 7856
rect 132134 7696 132137 7856
rect 134971 7696 134974 7856
rect 135134 7696 135137 7856
rect 136471 7696 136474 7856
rect 136634 7696 136637 7856
rect 137971 7696 137974 7856
rect 138134 7696 138137 7856
rect 140971 7696 140974 7856
rect 141134 7696 141137 7856
rect 142971 7696 142974 7856
rect 143134 7696 143137 7856
rect 146971 7696 146974 7856
rect 147134 7696 147137 7856
rect 148471 7696 148474 7856
rect 148634 7696 148637 7856
rect 149971 7696 149974 7856
rect 150134 7696 150137 7856
rect 151471 7696 151474 7856
rect 151634 7696 151637 7856
rect 60839 7690 60999 7695
rect 83774 7691 83934 7696
rect 90274 7691 90434 7696
rect 94774 7691 94934 7696
rect 99274 7691 99434 7696
rect 102274 7691 102434 7696
rect 105774 7691 105934 7696
rect 111774 7691 111934 7696
rect 116274 7691 116434 7696
rect 119274 7691 119434 7696
rect 125274 7691 125434 7696
rect 131974 7691 132134 7696
rect 134974 7691 135134 7696
rect 136474 7691 136634 7696
rect 137974 7691 138134 7696
rect 140974 7691 141134 7696
rect 142974 7691 143134 7696
rect 146974 7691 147134 7696
rect 148474 7691 148634 7696
rect 149974 7691 150134 7696
rect 151474 7691 151634 7696
rect 16457 7679 16617 7684
rect 32128 7683 32288 7688
<< via2 >>
rect 151254 162166 151354 162266
rect 151965 160521 152120 160676
rect 54 159861 154 159961
rect 151965 159021 152120 159176
rect 54 158361 154 158461
rect 151965 157521 152120 157676
rect 54 156861 154 156961
rect 151965 156021 152120 156176
rect 54 155361 154 155461
rect 151965 154521 152120 154676
rect 54 153861 154 153961
rect 151965 153021 152120 153176
rect 54 152361 154 152461
rect 151965 151521 152120 151676
rect 54 150861 154 150961
rect 151965 150021 152120 150176
rect 54 149361 154 149461
rect 151965 148521 152120 148676
rect 54 147861 154 147961
rect 151965 147021 152120 147176
rect 54 146361 154 146461
rect 151965 145521 152120 145676
rect 54 144861 154 144961
rect 151965 144021 152120 144176
rect 54 143361 154 143461
rect 151965 142521 152120 142676
rect 54 141861 154 141961
rect 151965 141021 152120 141176
rect 54 140361 154 140461
rect 151965 139521 152120 139676
rect 54 138861 154 138961
rect 151965 138021 152120 138176
rect 54 137361 154 137461
rect 151965 136521 152120 136676
rect 54 135861 154 135961
rect 151965 135021 152120 135176
rect 54 134361 154 134461
rect 151965 133521 152120 133676
rect 54 132861 154 132961
rect 151965 132021 152120 132176
rect 54 131361 154 131461
rect 151965 130521 152120 130676
rect 54 129861 154 129961
rect 151965 129021 152120 129176
rect 54 128361 154 128461
rect 151965 127521 152120 127676
rect 54 126861 154 126961
rect 151965 126021 152120 126176
rect 54 125361 154 125461
rect 151965 124521 152120 124676
rect 54 123861 154 123961
rect 151965 123021 152120 123176
rect 54 122361 154 122461
rect 151965 121521 152120 121676
rect 54 120861 154 120961
rect 151965 120021 152120 120176
rect 54 119361 154 119461
rect 151965 118521 152120 118676
rect 54 117861 154 117961
rect 151965 117021 152120 117176
rect 54 116361 154 116461
rect 151965 115521 152120 115676
rect 54 114861 154 114961
rect 151965 114021 152120 114176
rect 54 113361 154 113461
rect 151965 112521 152120 112676
rect 54 111861 154 111961
rect 151965 111021 152120 111176
rect 54 110361 154 110461
rect 151965 109521 152120 109676
rect 54 108861 154 108961
rect 151965 108021 152120 108176
rect 54 107361 154 107461
rect 151965 106521 152120 106676
rect 54 105861 154 105961
rect 151965 105021 152120 105176
rect 54 104361 154 104461
rect 151965 103521 152120 103676
rect 54 102861 154 102961
rect 151965 102021 152120 102176
rect 54 101361 154 101461
rect 151965 100521 152120 100676
rect 54 99861 154 99961
rect 151965 99021 152120 99176
rect 54 98361 154 98461
rect 151965 97521 152120 97676
rect 54 96861 154 96961
rect 151965 96021 152120 96176
rect 54 95361 154 95461
rect 151965 94521 152120 94676
rect 54 93861 154 93961
rect 151965 93021 152120 93176
rect 54 92361 154 92461
rect 151965 91521 152120 91676
rect 54 90861 154 90961
rect 151965 90021 152120 90176
rect 54 89361 154 89461
rect 151965 88521 152120 88676
rect 54 87861 154 87961
rect 151965 87021 152120 87176
rect 54 86361 154 86461
rect 151965 85521 152120 85676
rect 54 84861 154 84961
rect 151965 84021 152120 84176
rect 54 83361 154 83461
rect 151965 82521 152120 82676
rect 54 81861 154 81961
rect 151965 81021 152120 81176
rect 54 80361 154 80461
rect 151965 79521 152120 79676
rect 54 78861 154 78961
rect 151965 78021 152120 78176
rect 54 77361 154 77461
rect 151965 76521 152120 76676
rect 54 75861 154 75961
rect 151965 75021 152120 75176
rect 54 74361 154 74461
rect 151965 73521 152120 73676
rect 54 72861 154 72961
rect 151965 72021 152120 72176
rect 54 71361 154 71461
rect 151965 70521 152120 70676
rect 54 69861 154 69961
rect 151965 69021 152120 69176
rect 54 68361 154 68461
rect 151965 67521 152120 67676
rect 54 66861 154 66961
rect 151965 66021 152120 66176
rect 54 65361 154 65461
rect 151965 64521 152120 64676
rect 54 63861 154 63961
rect 151965 63021 152120 63176
rect 54 62361 154 62461
rect 151965 61521 152120 61676
rect 54 60861 154 60961
rect 151965 60021 152120 60176
rect 54 59361 154 59461
rect 151965 58521 152120 58676
rect 54 57861 154 57961
rect 151965 57021 152120 57176
rect 54 56361 154 56461
rect 151965 55521 152120 55676
rect 54 54861 154 54961
rect 151965 54021 152120 54176
rect 54 53361 154 53461
rect 151965 52521 152120 52676
rect 54 51861 154 51961
rect 151965 51021 152120 51176
rect 54 50361 154 50461
rect 151965 49521 152120 49676
rect 54 48861 154 48961
rect 151965 48021 152120 48176
rect 54 47361 154 47461
rect 151965 46521 152120 46676
rect 54 45861 154 45961
rect 151965 45021 152120 45176
rect 54 44361 154 44461
rect 151965 43521 152120 43676
rect 54 42861 154 42961
rect 151965 42021 152120 42176
rect 54 41361 154 41461
rect 151965 40521 152120 40676
rect 54 39861 154 39961
rect 151965 39021 152120 39176
rect 54 38361 154 38461
rect 151965 37521 152120 37676
rect 54 36861 154 36961
rect 151965 36021 152120 36176
rect 54 35361 154 35461
rect 151965 34521 152120 34676
rect 54 33861 154 33961
rect 151965 33021 152120 33176
rect 54 32361 154 32461
rect 151965 31521 152120 31676
rect 54 30861 154 30961
rect 151965 30021 152120 30176
rect 54 29361 154 29461
rect 151965 28521 152120 28676
rect 54 27861 154 27961
rect 151965 27021 152120 27176
rect 54 26361 154 26461
rect 151965 25521 152120 25676
rect 54 24861 154 24961
rect 151965 24021 152120 24176
rect 54 23361 154 23461
rect 151965 22521 152120 22676
rect 54 21861 154 21961
rect 151965 21021 152120 21176
rect 54 20361 154 20461
rect 151965 19521 152120 19676
rect 54 18861 154 18961
rect 151965 18021 152120 18176
rect 54 17361 154 17461
rect 151965 16521 152120 16676
rect 54 15861 154 15961
rect 151965 15021 152120 15176
rect 54 14361 154 14461
rect 151965 13521 152120 13676
rect 54 12861 154 12961
rect 151965 12021 152120 12176
rect 54 11361 154 11461
rect 151965 10521 152120 10676
rect 9937 9489 10042 9594
rect 1834 9222 1989 9377
rect 2666 9285 2771 9390
rect 3743 9338 3848 9443
rect 1166 9112 1271 9217
rect -3099 8873 -2999 8973
rect 5358 9310 5463 9415
rect 6903 9357 7008 9462
rect 8458 9301 8563 9406
rect 9046 9222 9201 9377
rect 12974 9398 13079 9503
rect 14542 9421 14652 9531
rect 11451 9222 11556 9327
rect 16166 9386 16271 9491
rect 17666 9420 17771 9525
rect 19166 9502 19271 9607
rect 16459 9222 16614 9377
rect 20666 9329 20771 9434
rect 22166 9354 22271 9459
rect 23666 9458 23771 9563
rect 25260 9398 25365 9503
rect 26771 9414 26876 9519
rect 28310 9474 28415 9579
rect 29817 9326 29922 9431
rect 31318 9288 31423 9393
rect 32130 9222 32285 9377
rect 32873 9333 32978 9438
rect 34277 9369 34382 9474
rect 37541 9408 37646 9513
rect 35966 9155 36071 9260
rect 40597 9248 40702 9353
rect 45208 9311 45313 9416
rect 39051 8933 39156 9038
rect 43670 9050 43775 9155
rect 42139 8885 42244 8990
rect 46780 9289 46885 9394
rect 48229 9330 48334 9435
rect 54453 9409 54558 9514
rect 51358 9263 51463 9368
rect 52840 9270 52945 9375
rect 49801 9143 49906 9248
rect 55976 9360 56081 9465
rect 57479 9385 57584 9490
rect 58986 9381 59091 9486
rect 60577 9325 60682 9430
rect 60841 9222 60996 9377
rect 62059 9316 62169 9426
rect 63623 9364 63728 9469
rect 65127 9299 65232 9404
rect 66706 9323 66816 9433
rect 69778 9193 69883 9298
rect 71302 9227 71407 9332
rect 72791 9314 72896 9419
rect 74379 9314 74484 9419
rect 68236 9013 68341 9118
rect 75888 9280 75993 9385
rect 77398 9322 77503 9427
rect 78924 9391 79029 9496
rect 87185 9460 87290 9565
rect 80445 9272 80550 9377
rect 81621 9122 81726 9227
rect 83776 9222 83931 9377
rect 86543 9137 86648 9242
rect 82966 8980 83071 9085
rect 84434 8603 84539 8708
rect 88166 9299 88271 9404
rect 90276 9222 90431 9377
rect 94776 9222 94931 9377
rect 99276 9222 99431 9377
rect 102276 9222 102431 9377
rect 103166 9120 103271 9225
rect 105776 9222 105931 9377
rect 107666 9174 107771 9279
rect 111776 9222 111931 9377
rect 114831 9362 114936 9467
rect 91239 8822 91344 8927
rect 92666 8911 92771 9016
rect 92007 8469 92112 8574
rect 98399 8857 98504 8962
rect 100460 8871 100565 8976
rect 94166 8722 94271 8827
rect 96735 8402 96840 8507
rect 103502 8768 103607 8873
rect 101004 8340 101109 8445
rect 106580 8942 106685 9047
rect 106954 8527 107059 8632
rect 113599 9107 113704 9212
rect 110666 8748 110771 8853
rect 110346 8507 110451 8612
rect 116276 9222 116431 9377
rect 116666 9237 116771 9342
rect 117327 9044 117432 9149
rect 119276 9222 119431 9377
rect 120838 9160 120943 9265
rect 121166 9178 121271 9283
rect 125276 9222 125431 9377
rect 120460 8900 120565 9005
rect 126965 9147 127070 9252
rect 127166 9243 127271 9348
rect 124836 8823 124941 8928
rect 124358 8431 124463 8536
rect 131976 9222 132131 9377
rect 134518 9173 134623 9278
rect 134976 9222 135131 9377
rect 136476 9222 136631 9377
rect 137976 9222 138131 9377
rect 139840 9242 139945 9347
rect 130524 8955 130629 9060
rect 130029 8516 130134 8621
rect 132937 8874 133042 8979
rect 134666 9027 134771 9132
rect 139441 8996 139546 9101
rect 138849 8684 138954 8789
rect 140976 9222 141131 9377
rect 142976 9222 143131 9377
rect 145166 9370 145271 9475
rect 152695 9442 152800 9547
rect 142166 8961 142271 9066
rect 146206 9006 146311 9111
rect 143467 8649 143572 8754
rect 146976 9222 147131 9377
rect 148476 9222 148631 9377
rect 149976 9222 150131 9377
rect 151476 9222 151631 9377
rect 149631 8754 149736 8859
rect 150128 8445 150233 8550
rect 151473 8047 151634 8208
rect 54 7694 154 7794
rect 1832 7687 1992 7847
rect 9044 7696 9204 7856
rect 16457 7684 16617 7844
rect 32128 7688 32288 7848
rect 60839 7695 60999 7855
rect 83774 7696 83934 7856
rect 90274 7696 90434 7856
rect 94774 7696 94934 7856
rect 99274 7696 99434 7856
rect 102274 7696 102434 7856
rect 105774 7696 105934 7856
rect 111774 7696 111934 7856
rect 116274 7696 116434 7856
rect 119274 7696 119434 7856
rect 125274 7696 125434 7856
rect 131974 7696 132134 7856
rect 134974 7696 135134 7856
rect 136474 7696 136634 7856
rect 137974 7696 138134 7856
rect 140974 7696 141134 7856
rect 142974 7696 143134 7856
rect 146974 7696 147134 7856
rect 148474 7696 148634 7856
rect 149974 7696 150134 7856
rect 151474 7696 151634 7856
<< metal3 >>
rect 454 161140 499 163683
rect 151251 162269 151356 162272
rect 151251 162166 151254 162169
rect 151354 162166 151356 162169
rect 151251 162164 151356 162166
rect 151963 160679 152122 160681
rect 151963 160678 152123 160679
rect 151963 160519 151963 160678
rect 152122 160519 152123 160678
rect 151963 160519 152123 160519
rect 151963 160516 152122 160519
rect 51 159961 156 159963
rect -1006 159861 -1003 159961
rect -903 159861 54 159961
rect 154 159861 156 159961
rect 51 159858 156 159861
rect 151963 159179 152122 159181
rect 151963 159178 152123 159179
rect 151963 159019 151963 159178
rect 152122 159019 152123 159178
rect 151963 159019 152123 159019
rect 151963 159016 152122 159019
rect 51 158461 156 158463
rect -1006 158361 -1003 158461
rect -903 158361 54 158461
rect 154 158361 156 158461
rect 51 158358 156 158361
rect 151963 157679 152122 157681
rect 151963 157678 152123 157679
rect 151963 157519 151963 157678
rect 152122 157519 152123 157678
rect 151963 157519 152123 157519
rect 151963 157516 152122 157519
rect 51 156961 156 156963
rect -1006 156861 -1003 156961
rect -903 156861 54 156961
rect 154 156861 156 156961
rect 51 156858 156 156861
rect 151963 156179 152122 156181
rect 151963 156178 152123 156179
rect 151963 156019 151963 156178
rect 152122 156019 152123 156178
rect 151963 156019 152123 156019
rect 151963 156016 152122 156019
rect 51 155461 156 155463
rect -1006 155361 -1003 155461
rect -903 155361 54 155461
rect 154 155361 156 155461
rect 51 155358 156 155361
rect 151963 154679 152122 154681
rect 151963 154678 152123 154679
rect 151963 154519 151963 154678
rect 152122 154519 152123 154678
rect 151963 154519 152123 154519
rect 151963 154516 152122 154519
rect 51 153961 156 153963
rect -1006 153861 -1003 153961
rect -903 153861 54 153961
rect 154 153861 156 153961
rect 51 153858 156 153861
rect 151963 153179 152122 153181
rect 151963 153178 152123 153179
rect 151963 153019 151963 153178
rect 152122 153019 152123 153178
rect 151963 153019 152123 153019
rect 151963 153016 152122 153019
rect 51 152461 156 152463
rect -1006 152361 -1003 152461
rect -903 152361 54 152461
rect 154 152361 156 152461
rect 51 152358 156 152361
rect 151963 151679 152122 151681
rect 151963 151678 152123 151679
rect 151963 151519 151963 151678
rect 152122 151519 152123 151678
rect 151963 151519 152123 151519
rect 151963 151516 152122 151519
rect 51 150961 156 150963
rect -1006 150861 -1003 150961
rect -903 150861 54 150961
rect 154 150861 156 150961
rect 51 150858 156 150861
rect 151963 150179 152122 150181
rect 151963 150178 152123 150179
rect 151963 150019 151963 150178
rect 152122 150019 152123 150178
rect 151963 150019 152123 150019
rect 151963 150016 152122 150019
rect 51 149461 156 149463
rect -1006 149361 -1003 149461
rect -903 149361 54 149461
rect 154 149361 156 149461
rect 51 149358 156 149361
rect 151963 148679 152122 148681
rect 151963 148678 152123 148679
rect 151963 148519 151963 148678
rect 152122 148519 152123 148678
rect 151963 148519 152123 148519
rect 151963 148516 152122 148519
rect 51 147961 156 147963
rect -1006 147861 -1003 147961
rect -903 147861 54 147961
rect 154 147861 156 147961
rect 51 147858 156 147861
rect 151963 147179 152122 147181
rect 151963 147178 152123 147179
rect 151963 147019 151963 147178
rect 152122 147019 152123 147178
rect 151963 147019 152123 147019
rect 151963 147016 152122 147019
rect 51 146461 156 146463
rect -1006 146361 -1003 146461
rect -903 146361 54 146461
rect 154 146361 156 146461
rect 51 146358 156 146361
rect 151963 145679 152122 145681
rect 151963 145678 152123 145679
rect 151963 145519 151963 145678
rect 152122 145519 152123 145678
rect 151963 145519 152123 145519
rect 151963 145516 152122 145519
rect 51 144961 156 144963
rect -1006 144861 -1003 144961
rect -903 144861 54 144961
rect 154 144861 156 144961
rect 51 144858 156 144861
rect 151963 144179 152122 144181
rect 151963 144178 152123 144179
rect 151963 144019 151963 144178
rect 152122 144019 152123 144178
rect 151963 144019 152123 144019
rect 151963 144016 152122 144019
rect 51 143461 156 143463
rect -1006 143361 -1003 143461
rect -903 143361 54 143461
rect 154 143361 156 143461
rect 51 143358 156 143361
rect 151963 142679 152122 142681
rect 151963 142678 152123 142679
rect 151963 142519 151963 142678
rect 152122 142519 152123 142678
rect 151963 142519 152123 142519
rect 151963 142516 152122 142519
rect 51 141961 156 141963
rect -1006 141861 -1003 141961
rect -903 141861 54 141961
rect 154 141861 156 141961
rect 51 141858 156 141861
rect 151963 141179 152122 141181
rect 151963 141178 152123 141179
rect 151963 141019 151963 141178
rect 152122 141019 152123 141178
rect 151963 141019 152123 141019
rect 151963 141016 152122 141019
rect 51 140461 156 140463
rect -1006 140361 -1003 140461
rect -903 140361 54 140461
rect 154 140361 156 140461
rect 51 140358 156 140361
rect 151963 139679 152122 139681
rect 151963 139678 152123 139679
rect 151963 139519 151963 139678
rect 152122 139519 152123 139678
rect 151963 139519 152123 139519
rect 151963 139516 152122 139519
rect 51 138961 156 138963
rect -1006 138861 -1003 138961
rect -903 138861 54 138961
rect 154 138861 156 138961
rect 51 138858 156 138861
rect 151963 138179 152122 138181
rect 151963 138178 152123 138179
rect 151963 138019 151963 138178
rect 152122 138019 152123 138178
rect 151963 138019 152123 138019
rect 151963 138016 152122 138019
rect 51 137461 156 137463
rect -1006 137361 -1003 137461
rect -903 137361 54 137461
rect 154 137361 156 137461
rect 51 137358 156 137361
rect 151963 136679 152122 136681
rect 151963 136678 152123 136679
rect 151963 136519 151963 136678
rect 152122 136519 152123 136678
rect 151963 136519 152123 136519
rect 151963 136516 152122 136519
rect 51 135961 156 135963
rect -1006 135861 -1003 135961
rect -903 135861 54 135961
rect 154 135861 156 135961
rect 51 135858 156 135861
rect 151963 135179 152122 135181
rect 151963 135178 152123 135179
rect 151963 135019 151963 135178
rect 152122 135019 152123 135178
rect 151963 135019 152123 135019
rect 151963 135016 152122 135019
rect 51 134461 156 134463
rect -1006 134361 -1003 134461
rect -903 134361 54 134461
rect 154 134361 156 134461
rect 51 134358 156 134361
rect 151963 133679 152122 133681
rect 151963 133678 152123 133679
rect 151963 133519 151963 133678
rect 152122 133519 152123 133678
rect 151963 133519 152123 133519
rect 151963 133516 152122 133519
rect 51 132961 156 132963
rect -1006 132861 -1003 132961
rect -903 132861 54 132961
rect 154 132861 156 132961
rect 51 132858 156 132861
rect 151963 132179 152122 132181
rect 151963 132178 152123 132179
rect 151963 132019 151963 132178
rect 152122 132019 152123 132178
rect 151963 132019 152123 132019
rect 151963 132016 152122 132019
rect 51 131461 156 131463
rect -1006 131361 -1003 131461
rect -903 131361 54 131461
rect 154 131361 156 131461
rect 51 131358 156 131361
rect 151963 130679 152122 130681
rect 151963 130678 152123 130679
rect 151963 130519 151963 130678
rect 152122 130519 152123 130678
rect 151963 130519 152123 130519
rect 151963 130516 152122 130519
rect 51 129961 156 129963
rect -1006 129861 -1003 129961
rect -903 129861 54 129961
rect 154 129861 156 129961
rect 51 129858 156 129861
rect 151963 129179 152122 129181
rect 151963 129178 152123 129179
rect 151963 129019 151963 129178
rect 152122 129019 152123 129178
rect 151963 129019 152123 129019
rect 151963 129016 152122 129019
rect 51 128461 156 128463
rect -1006 128361 -1003 128461
rect -903 128361 54 128461
rect 154 128361 156 128461
rect 51 128358 156 128361
rect 151963 127679 152122 127681
rect 151963 127678 152123 127679
rect 151963 127519 151963 127678
rect 152122 127519 152123 127678
rect 151963 127519 152123 127519
rect 151963 127516 152122 127519
rect 51 126961 156 126963
rect -1006 126861 -1003 126961
rect -903 126861 54 126961
rect 154 126861 156 126961
rect 51 126858 156 126861
rect 151963 126179 152122 126181
rect 151963 126178 152123 126179
rect 151963 126019 151963 126178
rect 152122 126019 152123 126178
rect 151963 126019 152123 126019
rect 151963 126016 152122 126019
rect 51 125461 156 125463
rect -1006 125361 -1003 125461
rect -903 125361 54 125461
rect 154 125361 156 125461
rect 51 125358 156 125361
rect 151963 124679 152122 124681
rect 151963 124678 152123 124679
rect 151963 124519 151963 124678
rect 152122 124519 152123 124678
rect 151963 124519 152123 124519
rect 151963 124516 152122 124519
rect 51 123961 156 123963
rect -1006 123861 -1003 123961
rect -903 123861 54 123961
rect 154 123861 156 123961
rect 51 123858 156 123861
rect 151963 123179 152122 123181
rect 151963 123178 152123 123179
rect 151963 123019 151963 123178
rect 152122 123019 152123 123178
rect 151963 123019 152123 123019
rect 151963 123016 152122 123019
rect 51 122461 156 122463
rect -1006 122361 -1003 122461
rect -903 122361 54 122461
rect 154 122361 156 122461
rect 51 122358 156 122361
rect 151963 121679 152122 121681
rect 151963 121678 152123 121679
rect 151963 121519 151963 121678
rect 152122 121519 152123 121678
rect 151963 121519 152123 121519
rect 151963 121516 152122 121519
rect 51 120961 156 120963
rect -1006 120861 -1003 120961
rect -903 120861 54 120961
rect 154 120861 156 120961
rect 51 120858 156 120861
rect 151963 120179 152122 120181
rect 151963 120178 152123 120179
rect 151963 120019 151963 120178
rect 152122 120019 152123 120178
rect 151963 120019 152123 120019
rect 151963 120016 152122 120019
rect 51 119461 156 119463
rect -1006 119361 -1003 119461
rect -903 119361 54 119461
rect 154 119361 156 119461
rect 51 119358 156 119361
rect 151963 118679 152122 118681
rect 151963 118678 152123 118679
rect 151963 118519 151963 118678
rect 152122 118519 152123 118678
rect 151963 118519 152123 118519
rect 151963 118516 152122 118519
rect 51 117961 156 117963
rect -1006 117861 -1003 117961
rect -903 117861 54 117961
rect 154 117861 156 117961
rect 51 117858 156 117861
rect 151963 117179 152122 117181
rect 151963 117178 152123 117179
rect 151963 117019 151963 117178
rect 152122 117019 152123 117178
rect 151963 117019 152123 117019
rect 151963 117016 152122 117019
rect 51 116461 156 116463
rect -1006 116361 -1003 116461
rect -903 116361 54 116461
rect 154 116361 156 116461
rect 51 116358 156 116361
rect 151963 115679 152122 115681
rect 151963 115678 152123 115679
rect 151963 115519 151963 115678
rect 152122 115519 152123 115678
rect 151963 115519 152123 115519
rect 151963 115516 152122 115519
rect 51 114961 156 114963
rect -1006 114861 -1003 114961
rect -903 114861 54 114961
rect 154 114861 156 114961
rect 51 114858 156 114861
rect 151963 114179 152122 114181
rect 151963 114178 152123 114179
rect 151963 114019 151963 114178
rect 152122 114019 152123 114178
rect 151963 114019 152123 114019
rect 151963 114016 152122 114019
rect 51 113461 156 113463
rect -1006 113361 -1003 113461
rect -903 113361 54 113461
rect 154 113361 156 113461
rect 51 113358 156 113361
rect 151963 112679 152122 112681
rect 151963 112678 152123 112679
rect 151963 112519 151963 112678
rect 152122 112519 152123 112678
rect 151963 112519 152123 112519
rect 151963 112516 152122 112519
rect 51 111961 156 111963
rect -1006 111861 -1003 111961
rect -903 111861 54 111961
rect 154 111861 156 111961
rect 51 111858 156 111861
rect 151963 111179 152122 111181
rect 151963 111178 152123 111179
rect 151963 111019 151963 111178
rect 152122 111019 152123 111178
rect 151963 111019 152123 111019
rect 151963 111016 152122 111019
rect 51 110461 156 110463
rect -1006 110361 -1003 110461
rect -903 110361 54 110461
rect 154 110361 156 110461
rect 51 110358 156 110361
rect 151963 109679 152122 109681
rect 151963 109678 152123 109679
rect 151963 109519 151963 109678
rect 152122 109519 152123 109678
rect 151963 109519 152123 109519
rect 151963 109516 152122 109519
rect 51 108961 156 108963
rect -1006 108861 -1003 108961
rect -903 108861 54 108961
rect 154 108861 156 108961
rect 51 108858 156 108861
rect 151963 108179 152122 108181
rect 151963 108178 152123 108179
rect 151963 108019 151963 108178
rect 152122 108019 152123 108178
rect 151963 108019 152123 108019
rect 151963 108016 152122 108019
rect 51 107461 156 107463
rect -1006 107361 -1003 107461
rect -903 107361 54 107461
rect 154 107361 156 107461
rect 51 107358 156 107361
rect 151963 106679 152122 106681
rect 151963 106678 152123 106679
rect 151963 106519 151963 106678
rect 152122 106519 152123 106678
rect 151963 106519 152123 106519
rect 151963 106516 152122 106519
rect 51 105961 156 105963
rect -1006 105861 -1003 105961
rect -903 105861 54 105961
rect 154 105861 156 105961
rect 51 105858 156 105861
rect 151963 105179 152122 105181
rect 151963 105178 152123 105179
rect 151963 105019 151963 105178
rect 152122 105019 152123 105178
rect 151963 105019 152123 105019
rect 151963 105016 152122 105019
rect 51 104461 156 104463
rect -1006 104361 -1003 104461
rect -903 104361 54 104461
rect 154 104361 156 104461
rect 51 104358 156 104361
rect 151963 103679 152122 103681
rect 151963 103678 152123 103679
rect 151963 103519 151963 103678
rect 152122 103519 152123 103678
rect 151963 103519 152123 103519
rect 151963 103516 152122 103519
rect 51 102961 156 102963
rect -1006 102861 -1003 102961
rect -903 102861 54 102961
rect 154 102861 156 102961
rect 51 102858 156 102861
rect 151963 102179 152122 102181
rect 151963 102178 152123 102179
rect 151963 102019 151963 102178
rect 152122 102019 152123 102178
rect 151963 102019 152123 102019
rect 151963 102016 152122 102019
rect 51 101461 156 101463
rect -1006 101361 -1003 101461
rect -903 101361 54 101461
rect 154 101361 156 101461
rect 51 101358 156 101361
rect 151963 100679 152122 100681
rect 151963 100678 152123 100679
rect 151963 100519 151963 100678
rect 152122 100519 152123 100678
rect 151963 100519 152123 100519
rect 151963 100516 152122 100519
rect 51 99961 156 99963
rect -1006 99861 -1003 99961
rect -903 99861 54 99961
rect 154 99861 156 99961
rect 51 99858 156 99861
rect 151963 99179 152122 99181
rect 151963 99178 152123 99179
rect 151963 99019 151963 99178
rect 152122 99019 152123 99178
rect 151963 99019 152123 99019
rect 151963 99016 152122 99019
rect 51 98461 156 98463
rect -1006 98361 -1003 98461
rect -903 98361 54 98461
rect 154 98361 156 98461
rect 51 98358 156 98361
rect 151963 97679 152122 97681
rect 151963 97678 152123 97679
rect 151963 97519 151963 97678
rect 152122 97519 152123 97678
rect 151963 97519 152123 97519
rect 151963 97516 152122 97519
rect 51 96961 156 96963
rect -1006 96861 -1003 96961
rect -903 96861 54 96961
rect 154 96861 156 96961
rect 51 96858 156 96861
rect 151963 96179 152122 96181
rect 151963 96178 152123 96179
rect 151963 96019 151963 96178
rect 152122 96019 152123 96178
rect 151963 96019 152123 96019
rect 151963 96016 152122 96019
rect 51 95461 156 95463
rect -1006 95361 -1003 95461
rect -903 95361 54 95461
rect 154 95361 156 95461
rect 51 95358 156 95361
rect 151963 94679 152122 94681
rect 151963 94678 152123 94679
rect 151963 94519 151963 94678
rect 152122 94519 152123 94678
rect 151963 94519 152123 94519
rect 151963 94516 152122 94519
rect 51 93961 156 93963
rect -1006 93861 -1003 93961
rect -903 93861 54 93961
rect 154 93861 156 93961
rect 51 93858 156 93861
rect 151963 93179 152122 93181
rect 151963 93178 152123 93179
rect 151963 93019 151963 93178
rect 152122 93019 152123 93178
rect 151963 93019 152123 93019
rect 151963 93016 152122 93019
rect 51 92461 156 92463
rect -1006 92361 -1003 92461
rect -903 92361 54 92461
rect 154 92361 156 92461
rect 51 92358 156 92361
rect 151963 91679 152122 91681
rect 151963 91678 152123 91679
rect 151963 91519 151963 91678
rect 152122 91519 152123 91678
rect 151963 91519 152123 91519
rect 151963 91516 152122 91519
rect 51 90961 156 90963
rect -1006 90861 -1003 90961
rect -903 90861 54 90961
rect 154 90861 156 90961
rect 51 90858 156 90861
rect 151963 90179 152122 90181
rect 151963 90178 152123 90179
rect 151963 90019 151963 90178
rect 152122 90019 152123 90178
rect 151963 90019 152123 90019
rect 151963 90016 152122 90019
rect 51 89461 156 89463
rect -1006 89361 -1003 89461
rect -903 89361 54 89461
rect 154 89361 156 89461
rect 51 89358 156 89361
rect 151963 88679 152122 88681
rect 151963 88678 152123 88679
rect 151963 88519 151963 88678
rect 152122 88519 152123 88678
rect 151963 88519 152123 88519
rect 151963 88516 152122 88519
rect 51 87961 156 87963
rect -1006 87861 -1003 87961
rect -903 87861 54 87961
rect 154 87861 156 87961
rect 51 87858 156 87861
rect 151963 87179 152122 87181
rect 151963 87178 152123 87179
rect 151963 87019 151963 87178
rect 152122 87019 152123 87178
rect 151963 87019 152123 87019
rect 151963 87016 152122 87019
rect 51 86461 156 86463
rect -1006 86361 -1003 86461
rect -903 86361 54 86461
rect 154 86361 156 86461
rect 51 86358 156 86361
rect 151963 85679 152122 85681
rect 151963 85678 152123 85679
rect 151963 85519 151963 85678
rect 152122 85519 152123 85678
rect 151963 85519 152123 85519
rect 151963 85516 152122 85519
rect 51 84961 156 84963
rect -1006 84861 -1003 84961
rect -903 84861 54 84961
rect 154 84861 156 84961
rect 51 84858 156 84861
rect 151963 84179 152122 84181
rect 151963 84178 152123 84179
rect 151963 84019 151963 84178
rect 152122 84019 152123 84178
rect 151963 84019 152123 84019
rect 151963 84016 152122 84019
rect 51 83461 156 83463
rect -1006 83361 -1003 83461
rect -903 83361 54 83461
rect 154 83361 156 83461
rect 51 83358 156 83361
rect 151963 82679 152122 82681
rect 151963 82678 152123 82679
rect 151963 82519 151963 82678
rect 152122 82519 152123 82678
rect 151963 82519 152123 82519
rect 151963 82516 152122 82519
rect 51 81961 156 81963
rect -1006 81861 -1003 81961
rect -903 81861 54 81961
rect 154 81861 156 81961
rect 51 81858 156 81861
rect 151963 81179 152122 81181
rect 151963 81178 152123 81179
rect 151963 81019 151963 81178
rect 152122 81019 152123 81178
rect 151963 81019 152123 81019
rect 151963 81016 152122 81019
rect 51 80461 156 80463
rect -1006 80361 -1003 80461
rect -903 80361 54 80461
rect 154 80361 156 80461
rect 51 80358 156 80361
rect 151963 79679 152122 79681
rect 151963 79678 152123 79679
rect 151963 79519 151963 79678
rect 152122 79519 152123 79678
rect 151963 79519 152123 79519
rect 151963 79516 152122 79519
rect 51 78961 156 78963
rect -1006 78861 -1003 78961
rect -903 78861 54 78961
rect 154 78861 156 78961
rect 51 78858 156 78861
rect 151963 78179 152122 78181
rect 151963 78178 152123 78179
rect 151963 78019 151963 78178
rect 152122 78019 152123 78178
rect 151963 78019 152123 78019
rect 151963 78016 152122 78019
rect 51 77461 156 77463
rect -1006 77361 -1003 77461
rect -903 77361 54 77461
rect 154 77361 156 77461
rect 51 77358 156 77361
rect 151963 76679 152122 76681
rect 151963 76678 152123 76679
rect 151963 76519 151963 76678
rect 152122 76519 152123 76678
rect 151963 76519 152123 76519
rect 151963 76516 152122 76519
rect 51 75961 156 75963
rect -1006 75861 -1003 75961
rect -903 75861 54 75961
rect 154 75861 156 75961
rect 51 75858 156 75861
rect 151963 75179 152122 75181
rect 151963 75178 152123 75179
rect 151963 75019 151963 75178
rect 152122 75019 152123 75178
rect 151963 75019 152123 75019
rect 151963 75016 152122 75019
rect 51 74461 156 74463
rect -1006 74361 -1003 74461
rect -903 74361 54 74461
rect 154 74361 156 74461
rect 51 74358 156 74361
rect 151963 73679 152122 73681
rect 151963 73678 152123 73679
rect 151963 73519 151963 73678
rect 152122 73519 152123 73678
rect 151963 73519 152123 73519
rect 151963 73516 152122 73519
rect 51 72961 156 72963
rect -1006 72861 -1003 72961
rect -903 72861 54 72961
rect 154 72861 156 72961
rect 51 72858 156 72861
rect 151963 72179 152122 72181
rect 151963 72178 152123 72179
rect 151963 72019 151963 72178
rect 152122 72019 152123 72178
rect 151963 72019 152123 72019
rect 151963 72016 152122 72019
rect 51 71461 156 71463
rect -1006 71361 -1003 71461
rect -903 71361 54 71461
rect 154 71361 156 71461
rect 51 71358 156 71361
rect 151963 70679 152122 70681
rect 151963 70678 152123 70679
rect 151963 70519 151963 70678
rect 152122 70519 152123 70678
rect 151963 70519 152123 70519
rect 151963 70516 152122 70519
rect 51 69961 156 69963
rect -1006 69861 -1003 69961
rect -903 69861 54 69961
rect 154 69861 156 69961
rect 51 69858 156 69861
rect 151963 69179 152122 69181
rect 151963 69178 152123 69179
rect 151963 69019 151963 69178
rect 152122 69019 152123 69178
rect 151963 69019 152123 69019
rect 151963 69016 152122 69019
rect 51 68461 156 68463
rect -1006 68361 -1003 68461
rect -903 68361 54 68461
rect 154 68361 156 68461
rect 51 68358 156 68361
rect 151963 67679 152122 67681
rect 151963 67678 152123 67679
rect 151963 67519 151963 67678
rect 152122 67519 152123 67678
rect 151963 67519 152123 67519
rect 151963 67516 152122 67519
rect 51 66961 156 66963
rect -1006 66861 -1003 66961
rect -903 66861 54 66961
rect 154 66861 156 66961
rect 51 66858 156 66861
rect 151963 66179 152122 66181
rect 151963 66178 152123 66179
rect 151963 66019 151963 66178
rect 152122 66019 152123 66178
rect 151963 66019 152123 66019
rect 151963 66016 152122 66019
rect 51 65461 156 65463
rect -1006 65361 -1003 65461
rect -903 65361 54 65461
rect 154 65361 156 65461
rect 51 65358 156 65361
rect 151963 64679 152122 64681
rect 151963 64678 152123 64679
rect 151963 64519 151963 64678
rect 152122 64519 152123 64678
rect 151963 64519 152123 64519
rect 151963 64516 152122 64519
rect 51 63961 156 63963
rect -1006 63861 -1003 63961
rect -903 63861 54 63961
rect 154 63861 156 63961
rect 51 63858 156 63861
rect 151963 63179 152122 63181
rect 151963 63178 152123 63179
rect 151963 63019 151963 63178
rect 152122 63019 152123 63178
rect 151963 63019 152123 63019
rect 151963 63016 152122 63019
rect 51 62461 156 62463
rect -1006 62361 -1003 62461
rect -903 62361 54 62461
rect 154 62361 156 62461
rect 51 62358 156 62361
rect 151963 61679 152122 61681
rect 151963 61678 152123 61679
rect 151963 61519 151963 61678
rect 152122 61519 152123 61678
rect 151963 61519 152123 61519
rect 151963 61516 152122 61519
rect 51 60961 156 60963
rect -1006 60861 -1003 60961
rect -903 60861 54 60961
rect 154 60861 156 60961
rect 51 60858 156 60861
rect 151963 60179 152122 60181
rect 151963 60178 152123 60179
rect 151963 60019 151963 60178
rect 152122 60019 152123 60178
rect 151963 60019 152123 60019
rect 151963 60016 152122 60019
rect 51 59461 156 59463
rect -1006 59361 -1003 59461
rect -903 59361 54 59461
rect 154 59361 156 59461
rect 51 59358 156 59361
rect 151963 58679 152122 58681
rect 151963 58678 152123 58679
rect 151963 58519 151963 58678
rect 152122 58519 152123 58678
rect 151963 58519 152123 58519
rect 151963 58516 152122 58519
rect 51 57961 156 57963
rect -1006 57861 -1003 57961
rect -903 57861 54 57961
rect 154 57861 156 57961
rect 51 57858 156 57861
rect 151963 57179 152122 57181
rect 151963 57178 152123 57179
rect 151963 57019 151963 57178
rect 152122 57019 152123 57178
rect 151963 57019 152123 57019
rect 151963 57016 152122 57019
rect 51 56461 156 56463
rect -1006 56361 -1003 56461
rect -903 56361 54 56461
rect 154 56361 156 56461
rect 51 56358 156 56361
rect 151963 55679 152122 55681
rect 151963 55678 152123 55679
rect 151963 55519 151963 55678
rect 152122 55519 152123 55678
rect 151963 55519 152123 55519
rect 151963 55516 152122 55519
rect 51 54961 156 54963
rect -1006 54861 -1003 54961
rect -903 54861 54 54961
rect 154 54861 156 54961
rect 51 54858 156 54861
rect 151963 54179 152122 54181
rect 151963 54178 152123 54179
rect 151963 54019 151963 54178
rect 152122 54019 152123 54178
rect 151963 54019 152123 54019
rect 151963 54016 152122 54019
rect 51 53461 156 53463
rect -1006 53361 -1003 53461
rect -903 53361 54 53461
rect 154 53361 156 53461
rect 51 53358 156 53361
rect 151963 52679 152122 52681
rect 151963 52678 152123 52679
rect 151963 52519 151963 52678
rect 152122 52519 152123 52678
rect 151963 52519 152123 52519
rect 151963 52516 152122 52519
rect 51 51961 156 51963
rect -1006 51861 -1003 51961
rect -903 51861 54 51961
rect 154 51861 156 51961
rect 51 51858 156 51861
rect 151963 51179 152122 51181
rect 151963 51178 152123 51179
rect 151963 51019 151963 51178
rect 152122 51019 152123 51178
rect 151963 51019 152123 51019
rect 151963 51016 152122 51019
rect 51 50461 156 50463
rect -1006 50361 -1003 50461
rect -903 50361 54 50461
rect 154 50361 156 50461
rect 51 50358 156 50361
rect 151963 49679 152122 49681
rect 151963 49678 152123 49679
rect 151963 49519 151963 49678
rect 152122 49519 152123 49678
rect 151963 49519 152123 49519
rect 151963 49516 152122 49519
rect 51 48961 156 48963
rect -1006 48861 -1003 48961
rect -903 48861 54 48961
rect 154 48861 156 48961
rect 51 48858 156 48861
rect 151963 48179 152122 48181
rect 151963 48178 152123 48179
rect 151963 48019 151963 48178
rect 152122 48019 152123 48178
rect 151963 48019 152123 48019
rect 151963 48016 152122 48019
rect 51 47461 156 47463
rect -1006 47361 -1003 47461
rect -903 47361 54 47461
rect 154 47361 156 47461
rect 51 47358 156 47361
rect 151963 46679 152122 46681
rect 151963 46678 152123 46679
rect 151963 46519 151963 46678
rect 152122 46519 152123 46678
rect 151963 46519 152123 46519
rect 151963 46516 152122 46519
rect 51 45961 156 45963
rect -1006 45861 -1003 45961
rect -903 45861 54 45961
rect 154 45861 156 45961
rect 51 45858 156 45861
rect 151963 45179 152122 45181
rect 151963 45178 152123 45179
rect 151963 45019 151963 45178
rect 152122 45019 152123 45178
rect 151963 45019 152123 45019
rect 151963 45016 152122 45019
rect 51 44461 156 44463
rect -1006 44361 -1003 44461
rect -903 44361 54 44461
rect 154 44361 156 44461
rect 51 44358 156 44361
rect 151963 43679 152122 43681
rect 151963 43678 152123 43679
rect 151963 43519 151963 43678
rect 152122 43519 152123 43678
rect 151963 43519 152123 43519
rect 151963 43516 152122 43519
rect 51 42961 156 42963
rect -1006 42861 -1003 42961
rect -903 42861 54 42961
rect 154 42861 156 42961
rect 51 42858 156 42861
rect 151963 42179 152122 42181
rect 151963 42178 152123 42179
rect 151963 42019 151963 42178
rect 152122 42019 152123 42178
rect 151963 42019 152123 42019
rect 151963 42016 152122 42019
rect 51 41461 156 41463
rect -1006 41361 -1003 41461
rect -903 41361 54 41461
rect 154 41361 156 41461
rect 51 41358 156 41361
rect 151963 40679 152122 40681
rect 151963 40678 152123 40679
rect 151963 40519 151963 40678
rect 152122 40519 152123 40678
rect 151963 40519 152123 40519
rect 151963 40516 152122 40519
rect 51 39961 156 39963
rect -1006 39861 -1003 39961
rect -903 39861 54 39961
rect 154 39861 156 39961
rect 51 39858 156 39861
rect 151963 39179 152122 39181
rect 151963 39178 152123 39179
rect 151963 39019 151963 39178
rect 152122 39019 152123 39178
rect 151963 39019 152123 39019
rect 151963 39016 152122 39019
rect 51 38461 156 38463
rect -1006 38361 -1003 38461
rect -903 38361 54 38461
rect 154 38361 156 38461
rect 51 38358 156 38361
rect 151963 37679 152122 37681
rect 151963 37678 152123 37679
rect 151963 37519 151963 37678
rect 152122 37519 152123 37678
rect 151963 37519 152123 37519
rect 151963 37516 152122 37519
rect 51 36961 156 36963
rect -1006 36861 -1003 36961
rect -903 36861 54 36961
rect 154 36861 156 36961
rect 51 36858 156 36861
rect 151963 36179 152122 36181
rect 151963 36178 152123 36179
rect 151963 36019 151963 36178
rect 152122 36019 152123 36178
rect 151963 36019 152123 36019
rect 151963 36016 152122 36019
rect 51 35461 156 35463
rect -1006 35361 -1003 35461
rect -903 35361 54 35461
rect 154 35361 156 35461
rect 51 35358 156 35361
rect 151963 34679 152122 34681
rect 151963 34678 152123 34679
rect 151963 34519 151963 34678
rect 152122 34519 152123 34678
rect 151963 34519 152123 34519
rect 151963 34516 152122 34519
rect 51 33961 156 33963
rect -1006 33861 -1003 33961
rect -903 33861 54 33961
rect 154 33861 156 33961
rect 51 33858 156 33861
rect 151963 33179 152122 33181
rect 151963 33178 152123 33179
rect 151963 33019 151963 33178
rect 152122 33019 152123 33178
rect 151963 33019 152123 33019
rect 151963 33016 152122 33019
rect 51 32461 156 32463
rect -1006 32361 -1003 32461
rect -903 32361 54 32461
rect 154 32361 156 32461
rect 51 32358 156 32361
rect 151963 31679 152122 31681
rect 151963 31678 152123 31679
rect 151963 31519 151963 31678
rect 152122 31519 152123 31678
rect 151963 31519 152123 31519
rect 151963 31516 152122 31519
rect 51 30961 156 30963
rect -1006 30861 -1003 30961
rect -903 30861 54 30961
rect 154 30861 156 30961
rect 51 30858 156 30861
rect 151963 30179 152122 30181
rect 151963 30178 152123 30179
rect 151963 30019 151963 30178
rect 152122 30019 152123 30178
rect 151963 30019 152123 30019
rect 151963 30016 152122 30019
rect 51 29461 156 29463
rect -1006 29361 -1003 29461
rect -903 29361 54 29461
rect 154 29361 156 29461
rect 51 29358 156 29361
rect 151963 28679 152122 28681
rect 151963 28678 152123 28679
rect 151963 28519 151963 28678
rect 152122 28519 152123 28678
rect 151963 28519 152123 28519
rect 151963 28516 152122 28519
rect 51 27961 156 27963
rect -1006 27861 -1003 27961
rect -903 27861 54 27961
rect 154 27861 156 27961
rect 51 27858 156 27861
rect 151963 27179 152122 27181
rect 151963 27178 152123 27179
rect 151963 27019 151963 27178
rect 152122 27019 152123 27178
rect 151963 27019 152123 27019
rect 151963 27016 152122 27019
rect 51 26461 156 26463
rect -1006 26361 -1003 26461
rect -903 26361 54 26461
rect 154 26361 156 26461
rect 51 26358 156 26361
rect 151963 25679 152122 25681
rect 151963 25678 152123 25679
rect 151963 25519 151963 25678
rect 152122 25519 152123 25678
rect 151963 25519 152123 25519
rect 151963 25516 152122 25519
rect 51 24961 156 24963
rect -1006 24861 -1003 24961
rect -903 24861 54 24961
rect 154 24861 156 24961
rect 51 24858 156 24861
rect 151963 24179 152122 24181
rect 151963 24178 152123 24179
rect 151963 24019 151963 24178
rect 152122 24019 152123 24178
rect 151963 24019 152123 24019
rect 151963 24016 152122 24019
rect 51 23461 156 23463
rect -1006 23361 -1003 23461
rect -903 23361 54 23461
rect 154 23361 156 23461
rect 51 23358 156 23361
rect 151963 22679 152122 22681
rect 151963 22678 152123 22679
rect 151963 22519 151963 22678
rect 152122 22519 152123 22678
rect 151963 22519 152123 22519
rect 151963 22516 152122 22519
rect 51 21961 156 21963
rect -1006 21861 -1003 21961
rect -903 21861 54 21961
rect 154 21861 156 21961
rect 51 21858 156 21861
rect 151963 21179 152122 21181
rect 151963 21178 152123 21179
rect 151963 21019 151963 21178
rect 152122 21019 152123 21178
rect 151963 21019 152123 21019
rect 151963 21016 152122 21019
rect 51 20461 156 20463
rect -1006 20361 -1003 20461
rect -903 20361 54 20461
rect 154 20361 156 20461
rect 51 20358 156 20361
rect 151963 19679 152122 19681
rect 151963 19678 152123 19679
rect 151963 19519 151963 19678
rect 152122 19519 152123 19678
rect 151963 19519 152123 19519
rect 151963 19516 152122 19519
rect 51 18961 156 18963
rect -1006 18861 -1003 18961
rect -903 18861 54 18961
rect 154 18861 156 18961
rect 51 18858 156 18861
rect 151963 18179 152122 18181
rect 151963 18178 152123 18179
rect 151963 18019 151963 18178
rect 152122 18019 152123 18178
rect 151963 18019 152123 18019
rect 151963 18016 152122 18019
rect 51 17461 156 17463
rect -1006 17361 -1003 17461
rect -903 17361 54 17461
rect 154 17361 156 17461
rect 51 17358 156 17361
rect 151963 16679 152122 16681
rect 151963 16678 152123 16679
rect 151963 16519 151963 16678
rect 152122 16519 152123 16678
rect 151963 16519 152123 16519
rect 151963 16516 152122 16519
rect 51 15961 156 15963
rect -1006 15861 -1003 15961
rect -903 15861 54 15961
rect 154 15861 156 15961
rect 51 15858 156 15861
rect 151963 15179 152122 15181
rect 151963 15178 152123 15179
rect 151963 15019 151963 15178
rect 152122 15019 152123 15178
rect 151963 15019 152123 15019
rect 151963 15016 152122 15019
rect 51 14461 156 14463
rect -1006 14361 -1003 14461
rect -903 14361 54 14461
rect 154 14361 156 14461
rect 51 14358 156 14361
rect 151963 13679 152122 13681
rect 151963 13678 152123 13679
rect 151963 13519 151963 13678
rect 152122 13519 152123 13678
rect 151963 13519 152123 13519
rect 151963 13516 152122 13519
rect 51 12961 156 12963
rect -1006 12861 -1003 12961
rect -903 12861 54 12961
rect 154 12861 156 12961
rect 51 12858 156 12861
rect 151963 12179 152122 12181
rect 151963 12178 152123 12179
rect 151963 12019 151963 12178
rect 152122 12019 152123 12178
rect 151963 12019 152123 12019
rect 151963 12016 152122 12019
rect 51 11461 156 11463
rect -1006 11361 -1003 11461
rect -903 11361 54 11461
rect 154 11361 156 11461
rect 51 11358 156 11361
rect 151963 10679 152122 10681
rect 151963 10678 152123 10679
rect 151963 10519 151963 10678
rect 152122 10519 152123 10678
rect 151963 10519 152123 10519
rect 151963 10516 152122 10519
rect 19164 9609 19274 9609
rect 9935 9597 10044 9599
rect 9934 9596 10044 9597
rect 9934 9487 9935 9596
rect 10044 9487 10044 9596
rect 14539 9531 14654 9533
rect 12972 9506 13081 9508
rect 9934 9487 10044 9487
rect 12971 9505 13081 9506
rect 9935 9484 10044 9487
rect 6901 9465 7010 9467
rect 6900 9464 7010 9465
rect 3741 9445 3851 9446
rect 2664 9392 2773 9395
rect 2664 9392 2774 9392
rect 1832 9379 1992 9380
rect 1829 9220 1832 9379
rect 1991 9220 1994 9379
rect 2664 9283 2664 9392
rect 2773 9283 2774 9392
rect 3738 9336 3741 9445
rect 3850 9336 3853 9445
rect 5356 9418 5465 9420
rect 5355 9417 5465 9418
rect 3741 9336 3851 9336
rect 5355 9308 5356 9417
rect 5465 9308 5465 9417
rect 6900 9355 6901 9464
rect 7010 9355 7010 9464
rect 8456 9408 8565 9411
rect 6900 9355 7010 9355
rect 8455 9408 8565 9408
rect 6901 9352 7010 9355
rect 5355 9308 5465 9308
rect 5356 9305 5465 9308
rect 8455 9299 8456 9408
rect 8565 9299 8565 9408
rect 12971 9396 12972 9505
rect 13081 9396 13081 9505
rect 14539 9421 14542 9531
rect 14652 9421 14654 9531
rect 17664 9527 17774 9528
rect 16164 9493 16273 9496
rect 14539 9418 14654 9421
rect 16164 9493 16274 9493
rect 12971 9396 13081 9396
rect 12972 9393 13081 9396
rect 16164 9384 16164 9493
rect 16273 9384 16274 9493
rect 17661 9418 17664 9527
rect 17773 9418 17776 9527
rect 19161 9500 19164 9609
rect 19273 9500 19276 9609
rect 28308 9581 28417 9584
rect 28307 9581 28417 9581
rect 23664 9565 23774 9565
rect 19164 9499 19274 9500
rect 22164 9461 22274 9462
rect 20664 9436 20774 9436
rect 17664 9418 17774 9418
rect 16164 9383 16274 9384
rect 16164 9381 16273 9383
rect 9044 9379 9204 9380
rect 16457 9379 16617 9380
rect 8455 9298 8565 9299
rect 8456 9296 8565 9298
rect 2664 9282 2774 9283
rect 2664 9280 2773 9282
rect 9041 9220 9044 9379
rect 9203 9220 9206 9379
rect 11449 9329 11558 9332
rect 11448 9329 11558 9329
rect 1832 9220 1992 9220
rect 9044 9220 9204 9220
rect 11448 9220 11449 9329
rect 11558 9220 11558 9329
rect 16454 9220 16457 9379
rect 16616 9220 16619 9379
rect 20661 9327 20664 9436
rect 20773 9327 20776 9436
rect 22161 9352 22164 9461
rect 22273 9352 22276 9461
rect 23661 9456 23664 9565
rect 23773 9456 23776 9565
rect 26769 9521 26878 9524
rect 26768 9521 26878 9521
rect 25258 9506 25367 9508
rect 25258 9505 25368 9506
rect 23664 9455 23774 9456
rect 25258 9396 25258 9505
rect 25367 9396 25368 9505
rect 26768 9412 26769 9521
rect 26878 9412 26878 9521
rect 28307 9472 28308 9581
rect 28417 9472 28417 9581
rect 87183 9567 87293 9568
rect 35964 9530 36073 9533
rect 35964 9530 36074 9530
rect 34164 9476 34385 9476
rect 28307 9471 28417 9472
rect 28308 9469 28417 9471
rect 32871 9441 32980 9443
rect 32871 9440 32981 9441
rect 29815 9433 29924 9436
rect 26768 9411 26878 9412
rect 29815 9433 29925 9433
rect 26769 9409 26878 9411
rect 25258 9396 25368 9396
rect 25258 9393 25367 9396
rect 22164 9352 22274 9352
rect 20664 9326 20774 9327
rect 29815 9324 29815 9433
rect 29924 9324 29925 9433
rect 31316 9395 31425 9398
rect 29815 9323 29925 9324
rect 31316 9395 31426 9395
rect 29815 9321 29924 9323
rect 31316 9286 31316 9395
rect 31425 9286 31426 9395
rect 32128 9379 32288 9380
rect 31316 9285 31426 9286
rect 31316 9283 31425 9285
rect 32125 9220 32128 9379
rect 32287 9220 32290 9379
rect 32871 9331 32871 9440
rect 32980 9331 32981 9440
rect 34161 9367 34164 9476
rect 34273 9474 34385 9476
rect 34273 9369 34277 9474
rect 34382 9369 34385 9474
rect 34273 9367 34385 9369
rect 34164 9366 34385 9367
rect 35964 9421 35964 9530
rect 36073 9421 36074 9530
rect 37539 9515 37648 9518
rect 54451 9516 54560 9519
rect 54450 9516 54560 9516
rect 32871 9331 32981 9331
rect 32871 9328 32980 9331
rect 35964 9260 36074 9421
rect 37539 9515 37649 9515
rect 37539 9406 37539 9515
rect 37648 9406 37649 9515
rect 40595 9452 40705 9453
rect 37539 9405 37649 9406
rect 37539 9403 37648 9405
rect 40592 9343 40595 9452
rect 40704 9343 40707 9452
rect 48226 9437 48336 9438
rect 45206 9418 45316 9419
rect 16457 9220 16617 9220
rect 32128 9220 32288 9220
rect 1164 9219 1274 9220
rect 11448 9219 11558 9220
rect 1161 9110 1164 9219
rect 1273 9110 1276 9219
rect 11449 9217 11558 9219
rect 35964 9155 35966 9260
rect 36071 9155 36074 9260
rect 40595 9248 40597 9343
rect 40702 9248 40705 9343
rect 45203 9309 45206 9418
rect 45315 9309 45318 9418
rect 46778 9396 46888 9397
rect 45206 9309 45316 9309
rect 46775 9287 46778 9396
rect 46887 9287 46890 9396
rect 48224 9328 48227 9437
rect 48336 9328 48339 9437
rect 54450 9407 54451 9516
rect 54560 9407 54560 9516
rect 78922 9499 79031 9501
rect 78921 9498 79031 9499
rect 57477 9492 57586 9495
rect 57476 9492 57586 9492
rect 55974 9468 56083 9470
rect 54450 9406 54560 9407
rect 55974 9467 56084 9468
rect 54451 9404 54560 9406
rect 52837 9377 52947 9378
rect 51356 9370 51465 9373
rect 51355 9370 51465 9370
rect 48226 9328 48336 9328
rect 46778 9287 46888 9287
rect 51355 9261 51356 9370
rect 51465 9261 51465 9370
rect 52835 9268 52838 9377
rect 52947 9268 52950 9377
rect 55974 9358 55974 9467
rect 56083 9358 56084 9467
rect 57476 9383 57477 9492
rect 57586 9383 57586 9492
rect 58984 9489 59093 9491
rect 57476 9382 57586 9383
rect 58984 9488 59094 9489
rect 57477 9380 57586 9382
rect 58984 9379 58984 9488
rect 59093 9379 59094 9488
rect 63621 9471 63730 9474
rect 63620 9471 63730 9471
rect 60575 9432 60684 9435
rect 58984 9379 59094 9379
rect 60575 9432 60685 9432
rect 58984 9376 59093 9379
rect 55974 9358 56084 9358
rect 55974 9355 56083 9358
rect 60575 9323 60575 9432
rect 60684 9323 60685 9432
rect 62056 9426 62171 9428
rect 60839 9379 60999 9380
rect 60575 9322 60685 9323
rect 60575 9320 60684 9322
rect 52837 9268 52947 9268
rect 51355 9260 51465 9261
rect 51356 9258 51465 9260
rect 49799 9251 49908 9253
rect 40595 9245 40705 9248
rect 49798 9250 49908 9251
rect 42137 9202 42246 9204
rect 42137 9201 42247 9202
rect 35964 9152 36074 9155
rect 39049 9153 39158 9156
rect 39049 9153 39159 9153
rect 1164 9110 1274 9110
rect 39049 9044 39049 9153
rect 39158 9044 39159 9153
rect 39049 9038 39159 9044
rect -3102 8973 -2997 8976
rect -3102 8971 -3099 8973
rect -2999 8971 -2997 8973
rect 39049 8933 39051 9038
rect 39156 8933 39159 9038
rect 39049 8931 39159 8933
rect 42137 9092 42137 9201
rect 42246 9092 42247 9201
rect 43668 9157 43777 9160
rect 42137 8990 42247 9092
rect 43667 9157 43777 9157
rect 43667 9048 43668 9157
rect 43777 9048 43777 9157
rect 49798 9141 49799 9250
rect 49908 9141 49908 9250
rect 60836 9220 60839 9379
rect 60998 9220 61001 9379
rect 62056 9316 62059 9426
rect 62169 9316 62171 9426
rect 63620 9362 63621 9471
rect 63730 9362 63730 9471
rect 66703 9433 66818 9436
rect 65125 9407 65234 9409
rect 63620 9361 63730 9362
rect 65125 9406 65235 9407
rect 63621 9359 63730 9361
rect 62056 9313 62171 9316
rect 65125 9297 65125 9406
rect 65234 9297 65235 9406
rect 66703 9323 66706 9433
rect 66816 9323 66818 9433
rect 77396 9429 77505 9432
rect 77396 9429 77506 9429
rect 72789 9422 72898 9424
rect 74377 9422 74486 9424
rect 72789 9421 72899 9422
rect 71300 9334 71409 9337
rect 66703 9321 66818 9323
rect 71299 9334 71409 9334
rect 69776 9300 69885 9303
rect 65125 9297 65235 9297
rect 69776 9300 69886 9300
rect 65125 9294 65234 9297
rect 60839 9220 60999 9220
rect 69776 9191 69776 9300
rect 69885 9191 69886 9300
rect 71299 9225 71300 9334
rect 71409 9225 71409 9334
rect 72789 9312 72789 9421
rect 72898 9312 72899 9421
rect 72789 9312 72899 9312
rect 74377 9421 74487 9422
rect 74377 9312 74377 9421
rect 74486 9312 74487 9421
rect 75886 9387 75995 9390
rect 74377 9312 74487 9312
rect 75886 9387 75996 9387
rect 72789 9309 72898 9312
rect 74377 9309 74486 9312
rect 75886 9278 75886 9387
rect 75995 9278 75996 9387
rect 77396 9320 77396 9429
rect 77505 9320 77506 9429
rect 78921 9389 78922 9498
rect 79031 9389 79031 9498
rect 87180 9458 87183 9567
rect 87292 9458 87295 9567
rect 152693 9550 152802 9552
rect 152692 9549 152802 9550
rect 145164 9478 145273 9480
rect 145164 9477 145274 9478
rect 114829 9469 114939 9470
rect 87183 9458 87293 9458
rect 88164 9406 88274 9406
rect 78921 9389 79031 9389
rect 78922 9386 79031 9389
rect 83774 9379 83934 9380
rect 80443 9379 80553 9379
rect 77396 9319 77506 9320
rect 77396 9317 77505 9319
rect 75886 9277 75996 9278
rect 75886 9275 75995 9277
rect 80440 9270 80443 9379
rect 80552 9270 80555 9379
rect 80443 9269 80553 9270
rect 81619 9229 81729 9230
rect 71299 9224 71409 9225
rect 71300 9222 71409 9224
rect 69776 9190 69886 9191
rect 69776 9188 69885 9190
rect 49798 9141 49908 9141
rect 49799 9138 49908 9141
rect 68233 9120 68343 9121
rect 81616 9120 81619 9229
rect 81728 9120 81731 9229
rect 83771 9220 83774 9379
rect 83933 9220 83936 9379
rect 88161 9297 88164 9406
rect 88273 9297 88276 9406
rect 90274 9379 90434 9380
rect 94774 9379 94934 9380
rect 99274 9379 99434 9380
rect 102274 9379 102434 9380
rect 105774 9379 105934 9380
rect 111774 9379 111934 9380
rect 88164 9296 88274 9297
rect 86541 9245 86650 9247
rect 86541 9244 86651 9245
rect 83774 9220 83934 9220
rect 86541 9135 86541 9244
rect 86650 9135 86651 9244
rect 90271 9220 90274 9379
rect 90433 9220 90436 9379
rect 94771 9220 94774 9379
rect 94933 9220 94936 9379
rect 99271 9220 99274 9379
rect 99433 9220 99436 9379
rect 102271 9220 102274 9379
rect 102433 9220 102436 9379
rect 103164 9228 103273 9230
rect 103164 9227 103274 9228
rect 90274 9220 90434 9220
rect 94774 9220 94934 9220
rect 99274 9220 99434 9220
rect 102274 9220 102434 9220
rect 86541 9135 86651 9135
rect 86541 9132 86650 9135
rect 43667 9047 43777 9048
rect 43668 9045 43777 9047
rect 68231 9011 68234 9120
rect 68343 9011 68346 9120
rect 81619 9120 81729 9120
rect 103164 9118 103164 9227
rect 103273 9118 103274 9227
rect 105771 9220 105774 9379
rect 105933 9220 105936 9379
rect 107664 9282 107773 9284
rect 107664 9281 107774 9282
rect 105774 9220 105934 9220
rect 107664 9172 107664 9281
rect 107773 9172 107774 9281
rect 111771 9220 111774 9379
rect 111933 9220 111936 9379
rect 114826 9360 114829 9469
rect 114938 9360 114941 9469
rect 116274 9379 116434 9380
rect 119274 9379 119434 9380
rect 125274 9379 125434 9380
rect 131974 9379 132134 9380
rect 134974 9379 135134 9380
rect 136474 9379 136634 9380
rect 137974 9379 138134 9380
rect 140974 9379 141134 9380
rect 142974 9379 143134 9380
rect 114829 9360 114939 9360
rect 116271 9220 116274 9379
rect 116433 9220 116436 9379
rect 116664 9345 116773 9347
rect 116664 9344 116774 9345
rect 116664 9235 116664 9344
rect 116773 9235 116774 9344
rect 116664 9235 116774 9235
rect 116664 9232 116773 9235
rect 119271 9220 119274 9379
rect 119433 9220 119436 9379
rect 121164 9285 121273 9288
rect 121164 9285 121274 9285
rect 120836 9267 120945 9270
rect 120836 9267 120946 9267
rect 111774 9220 111934 9220
rect 116274 9220 116434 9220
rect 119274 9220 119434 9220
rect 113597 9214 113707 9214
rect 107664 9172 107774 9172
rect 107664 9169 107773 9172
rect 103164 9118 103274 9118
rect 103164 9115 103273 9118
rect 113594 9105 113597 9214
rect 113706 9105 113709 9214
rect 120836 9158 120836 9267
rect 120945 9158 120946 9267
rect 121164 9176 121164 9285
rect 121273 9176 121274 9285
rect 125271 9220 125274 9379
rect 125433 9220 125436 9379
rect 127164 9350 127273 9353
rect 127164 9350 127274 9350
rect 126962 9254 127072 9255
rect 125274 9220 125434 9220
rect 121164 9175 121274 9176
rect 121164 9173 121273 9175
rect 120836 9157 120946 9158
rect 120836 9155 120945 9157
rect 117325 9151 117435 9152
rect 113597 9104 113707 9105
rect 82964 9087 83073 9090
rect 82964 9087 83074 9087
rect 68233 9011 68343 9011
rect 42137 8885 42139 8990
rect 42244 8885 42247 8990
rect 82964 8978 82964 9087
rect 83073 8978 83074 9087
rect 106578 9049 106687 9052
rect 106577 9049 106687 9049
rect 92664 9018 92773 9021
rect 82964 8977 83074 8978
rect 92664 9018 92774 9018
rect 82964 8975 83073 8977
rect 91236 8929 91346 8930
rect 42137 8882 42247 8885
rect -3102 8868 -2997 8871
rect 91234 8820 91237 8929
rect 91346 8820 91349 8929
rect 92664 8909 92664 9018
rect 92773 8909 92774 9018
rect 100458 8978 100567 8981
rect 100457 8978 100567 8978
rect 98396 8964 98506 8965
rect 92664 8908 92774 8909
rect 92664 8906 92773 8908
rect 98394 8855 98397 8964
rect 98506 8855 98509 8964
rect 100457 8869 100458 8978
rect 100567 8869 100567 8978
rect 106577 8940 106578 9049
rect 106687 8940 106687 9049
rect 117322 9042 117325 9151
rect 117434 9042 117437 9151
rect 126960 9145 126963 9254
rect 127072 9145 127075 9254
rect 127164 9241 127164 9350
rect 127273 9241 127274 9350
rect 127164 9240 127274 9241
rect 127164 9238 127273 9240
rect 131971 9220 131974 9379
rect 132133 9220 132136 9379
rect 134516 9280 134626 9280
rect 131974 9220 132134 9220
rect 134513 9171 134516 9280
rect 134625 9171 134628 9280
rect 134971 9220 134974 9379
rect 135133 9220 135136 9379
rect 136471 9220 136474 9379
rect 136633 9220 136636 9379
rect 137971 9220 137974 9379
rect 138133 9220 138136 9379
rect 139838 9349 139948 9349
rect 139835 9240 139838 9349
rect 139947 9240 139950 9349
rect 139838 9239 139948 9240
rect 140971 9220 140974 9379
rect 141133 9220 141136 9379
rect 142971 9220 142974 9379
rect 143133 9220 143136 9379
rect 145164 9368 145164 9477
rect 145273 9368 145274 9477
rect 152692 9440 152693 9549
rect 152802 9440 152802 9549
rect 152692 9440 152802 9440
rect 152693 9437 152802 9440
rect 146974 9379 147134 9380
rect 148474 9379 148634 9380
rect 149974 9379 150134 9380
rect 151474 9379 151634 9380
rect 145164 9368 145274 9368
rect 145164 9365 145273 9368
rect 146971 9220 146974 9379
rect 147133 9220 147136 9379
rect 148471 9220 148474 9379
rect 148633 9220 148636 9379
rect 149971 9220 149974 9379
rect 150133 9220 150136 9379
rect 151471 9220 151474 9379
rect 151633 9220 151636 9379
rect 134974 9220 135134 9220
rect 136474 9220 136634 9220
rect 137974 9220 138134 9220
rect 140974 9220 141134 9220
rect 142974 9220 143134 9220
rect 146974 9220 147134 9220
rect 148474 9220 148634 9220
rect 149974 9220 150134 9220
rect 151474 9220 151634 9220
rect 134516 9170 134626 9171
rect 126962 9145 127072 9145
rect 134664 9134 134773 9137
rect 134664 9134 134774 9134
rect 130522 9063 130631 9065
rect 130522 9062 130632 9063
rect 117325 9042 117435 9042
rect 120458 9008 120567 9010
rect 106577 8939 106687 8940
rect 120458 9007 120568 9008
rect 106578 8937 106687 8939
rect 120458 8898 120458 9007
rect 120567 8898 120568 9007
rect 130522 8953 130522 9062
rect 130631 8953 130632 9062
rect 134664 9025 134664 9134
rect 134773 9025 134774 9134
rect 146203 9113 146313 9114
rect 139439 9103 139549 9103
rect 134664 9024 134774 9025
rect 134664 9022 134773 9024
rect 139436 8994 139439 9103
rect 139548 8994 139551 9103
rect 142164 9069 142273 9071
rect 142164 9068 142274 9069
rect 139439 8993 139549 8994
rect 132935 8982 133044 8984
rect 130522 8953 130632 8953
rect 132935 8981 133045 8982
rect 130522 8950 130631 8953
rect 124833 8930 124943 8930
rect 120458 8898 120568 8898
rect 120458 8895 120567 8898
rect 103500 8876 103609 8878
rect 100457 8868 100567 8869
rect 103499 8875 103609 8876
rect 100458 8866 100567 8868
rect 98396 8855 98506 8855
rect 94164 8830 94273 8832
rect 94164 8829 94274 8830
rect 91236 8820 91346 8820
rect 94164 8720 94164 8829
rect 94273 8720 94274 8829
rect 103499 8766 103500 8875
rect 103609 8766 103609 8875
rect 110664 8856 110773 8858
rect 103499 8766 103609 8766
rect 110664 8855 110774 8856
rect 103500 8763 103609 8766
rect 110664 8746 110664 8855
rect 110773 8746 110774 8855
rect 124831 8821 124834 8930
rect 124943 8821 124946 8930
rect 132935 8872 132935 8981
rect 133044 8872 133045 8981
rect 142164 8959 142164 9068
rect 142273 8959 142274 9068
rect 146201 9004 146204 9113
rect 146313 9004 146316 9113
rect 146203 9004 146313 9004
rect 142164 8959 142274 8959
rect 142164 8956 142273 8959
rect 132935 8872 133045 8872
rect 132935 8869 133044 8872
rect 149629 8862 149738 8864
rect 149629 8861 149739 8862
rect 124833 8820 124943 8821
rect 138846 8791 138956 8791
rect 110664 8746 110774 8746
rect 110664 8743 110773 8746
rect 94164 8720 94274 8720
rect 94164 8717 94273 8720
rect 84432 8711 84541 8713
rect 84431 8710 84541 8711
rect 84431 8601 84432 8710
rect 84541 8601 84541 8710
rect 138844 8682 138847 8791
rect 138956 8682 138959 8791
rect 143465 8756 143574 8759
rect 143464 8756 143574 8756
rect 138846 8681 138956 8682
rect 143464 8647 143465 8756
rect 143574 8647 143574 8756
rect 149629 8752 149629 8861
rect 149738 8752 149739 8861
rect 149629 8752 149739 8752
rect 149629 8749 149738 8752
rect 143464 8646 143574 8647
rect 143465 8644 143574 8646
rect 106952 8635 107061 8637
rect 84431 8601 84541 8601
rect 106952 8634 107062 8635
rect 84432 8598 84541 8601
rect 92005 8576 92114 8579
rect 92005 8576 92115 8576
rect 92005 8467 92005 8576
rect 92114 8467 92115 8576
rect 106952 8525 106952 8634
rect 107061 8525 107062 8634
rect 130027 8623 130136 8626
rect 130026 8623 130136 8623
rect 110344 8614 110453 8617
rect 106952 8525 107062 8525
rect 110344 8614 110454 8614
rect 106952 8522 107061 8525
rect 96733 8510 96842 8512
rect 92005 8466 92115 8467
rect 96732 8509 96842 8510
rect 92005 8464 92114 8466
rect 96732 8400 96733 8509
rect 96842 8400 96842 8509
rect 110344 8505 110344 8614
rect 110453 8505 110454 8614
rect 124356 8539 124465 8541
rect 110344 8504 110454 8505
rect 124355 8538 124465 8539
rect 110344 8502 110453 8504
rect 101002 8447 101111 8450
rect 96732 8400 96842 8400
rect 101001 8447 101111 8447
rect 96733 8397 96842 8400
rect 101001 8338 101002 8447
rect 101111 8338 101111 8447
rect 124355 8429 124356 8538
rect 124465 8429 124465 8538
rect 130026 8514 130027 8623
rect 130136 8514 130136 8623
rect 150126 8553 150235 8555
rect 130026 8513 130136 8514
rect 150125 8552 150235 8553
rect 130027 8511 130136 8513
rect 150125 8443 150126 8552
rect 150235 8443 150235 8552
rect 150125 8443 150235 8443
rect 150126 8440 150235 8443
rect 124355 8429 124465 8429
rect 124356 8426 124465 8429
rect 101001 8337 101111 8338
rect 101002 8335 101111 8337
rect 151471 8208 151637 8210
rect 151471 8205 151473 8208
rect 151634 8205 151637 8208
rect 151471 8041 151637 8044
rect 9041 7856 9206 7858
rect 9041 7853 9044 7856
rect 9204 7853 9206 7856
rect 1829 7847 1994 7849
rect 1829 7844 1832 7847
rect 1992 7844 1994 7847
rect 51 7794 156 7796
rect 51 7791 54 7794
rect 154 7791 156 7794
rect 51 7688 156 7691
rect 60836 7855 61001 7857
rect 60836 7852 60839 7855
rect 60999 7852 61001 7855
rect 32125 7848 32290 7850
rect 9041 7690 9206 7693
rect 16454 7844 16619 7846
rect 16454 7841 16457 7844
rect 16617 7841 16619 7844
rect 1829 7681 1994 7684
rect 32125 7845 32128 7848
rect 32288 7845 32290 7848
rect 60836 7689 61001 7692
rect 83771 7856 83936 7858
rect 83771 7853 83774 7856
rect 83934 7853 83936 7856
rect 83771 7690 83936 7693
rect 90271 7856 90436 7858
rect 90271 7853 90274 7856
rect 90434 7853 90436 7856
rect 90271 7690 90436 7693
rect 94771 7856 94936 7858
rect 94771 7853 94774 7856
rect 94934 7853 94936 7856
rect 94771 7690 94936 7693
rect 99271 7856 99436 7858
rect 99271 7853 99274 7856
rect 99434 7853 99436 7856
rect 99271 7690 99436 7693
rect 102271 7856 102436 7858
rect 102271 7853 102274 7856
rect 102434 7853 102436 7856
rect 102271 7690 102436 7693
rect 105771 7856 105936 7858
rect 105771 7853 105774 7856
rect 105934 7853 105936 7856
rect 105771 7690 105936 7693
rect 111771 7856 111936 7858
rect 111771 7853 111774 7856
rect 111934 7853 111936 7856
rect 111771 7690 111936 7693
rect 116271 7856 116436 7858
rect 116271 7853 116274 7856
rect 116434 7853 116436 7856
rect 116271 7690 116436 7693
rect 119271 7856 119436 7858
rect 119271 7853 119274 7856
rect 119434 7853 119436 7856
rect 119271 7690 119436 7693
rect 125271 7856 125436 7858
rect 125271 7853 125274 7856
rect 125434 7853 125436 7856
rect 125271 7690 125436 7693
rect 131971 7856 132136 7858
rect 131971 7853 131974 7856
rect 132134 7853 132136 7856
rect 131971 7690 132136 7693
rect 134971 7856 135136 7858
rect 134971 7853 134974 7856
rect 135134 7853 135136 7856
rect 134971 7690 135136 7693
rect 136471 7856 136636 7858
rect 136471 7853 136474 7856
rect 136634 7853 136636 7856
rect 136471 7690 136636 7693
rect 137971 7856 138136 7858
rect 137971 7853 137974 7856
rect 138134 7853 138136 7856
rect 137971 7690 138136 7693
rect 140971 7856 141136 7858
rect 140971 7853 140974 7856
rect 141134 7853 141136 7856
rect 140971 7690 141136 7693
rect 142971 7856 143136 7858
rect 142971 7853 142974 7856
rect 143134 7853 143136 7856
rect 142971 7690 143136 7693
rect 146971 7856 147136 7858
rect 146971 7853 146974 7856
rect 147134 7853 147136 7856
rect 146971 7690 147136 7693
rect 148471 7856 148636 7858
rect 148471 7853 148474 7856
rect 148634 7853 148636 7856
rect 148471 7690 148636 7693
rect 149971 7856 150136 7858
rect 149971 7853 149974 7856
rect 150134 7853 150136 7856
rect 149971 7690 150136 7693
rect 151471 7856 151636 7858
rect 151471 7853 151474 7856
rect 151634 7853 151636 7856
rect 151471 7690 151636 7693
rect 32125 7682 32290 7685
rect 16454 7678 16619 7681
<< via3 >>
rect 151251 162266 151356 162269
rect 151251 162169 151254 162266
rect 151254 162169 151354 162266
rect 151354 162169 151356 162266
rect 151963 160676 152122 160678
rect 151963 160521 151965 160676
rect 151965 160521 152120 160676
rect 152120 160521 152122 160676
rect 151963 160519 152122 160521
rect -1003 159861 -903 159961
rect 151963 159176 152122 159178
rect 151963 159021 151965 159176
rect 151965 159021 152120 159176
rect 152120 159021 152122 159176
rect 151963 159019 152122 159021
rect -1003 158361 -903 158461
rect 151963 157676 152122 157678
rect 151963 157521 151965 157676
rect 151965 157521 152120 157676
rect 152120 157521 152122 157676
rect 151963 157519 152122 157521
rect -1003 156861 -903 156961
rect 151963 156176 152122 156178
rect 151963 156021 151965 156176
rect 151965 156021 152120 156176
rect 152120 156021 152122 156176
rect 151963 156019 152122 156021
rect -1003 155361 -903 155461
rect 151963 154676 152122 154678
rect 151963 154521 151965 154676
rect 151965 154521 152120 154676
rect 152120 154521 152122 154676
rect 151963 154519 152122 154521
rect -1003 153861 -903 153961
rect 151963 153176 152122 153178
rect 151963 153021 151965 153176
rect 151965 153021 152120 153176
rect 152120 153021 152122 153176
rect 151963 153019 152122 153021
rect -1003 152361 -903 152461
rect 151963 151676 152122 151678
rect 151963 151521 151965 151676
rect 151965 151521 152120 151676
rect 152120 151521 152122 151676
rect 151963 151519 152122 151521
rect -1003 150861 -903 150961
rect 151963 150176 152122 150178
rect 151963 150021 151965 150176
rect 151965 150021 152120 150176
rect 152120 150021 152122 150176
rect 151963 150019 152122 150021
rect -1003 149361 -903 149461
rect 151963 148676 152122 148678
rect 151963 148521 151965 148676
rect 151965 148521 152120 148676
rect 152120 148521 152122 148676
rect 151963 148519 152122 148521
rect -1003 147861 -903 147961
rect 151963 147176 152122 147178
rect 151963 147021 151965 147176
rect 151965 147021 152120 147176
rect 152120 147021 152122 147176
rect 151963 147019 152122 147021
rect -1003 146361 -903 146461
rect 151963 145676 152122 145678
rect 151963 145521 151965 145676
rect 151965 145521 152120 145676
rect 152120 145521 152122 145676
rect 151963 145519 152122 145521
rect -1003 144861 -903 144961
rect 151963 144176 152122 144178
rect 151963 144021 151965 144176
rect 151965 144021 152120 144176
rect 152120 144021 152122 144176
rect 151963 144019 152122 144021
rect -1003 143361 -903 143461
rect 151963 142676 152122 142678
rect 151963 142521 151965 142676
rect 151965 142521 152120 142676
rect 152120 142521 152122 142676
rect 151963 142519 152122 142521
rect -1003 141861 -903 141961
rect 151963 141176 152122 141178
rect 151963 141021 151965 141176
rect 151965 141021 152120 141176
rect 152120 141021 152122 141176
rect 151963 141019 152122 141021
rect -1003 140361 -903 140461
rect 151963 139676 152122 139678
rect 151963 139521 151965 139676
rect 151965 139521 152120 139676
rect 152120 139521 152122 139676
rect 151963 139519 152122 139521
rect -1003 138861 -903 138961
rect 151963 138176 152122 138178
rect 151963 138021 151965 138176
rect 151965 138021 152120 138176
rect 152120 138021 152122 138176
rect 151963 138019 152122 138021
rect -1003 137361 -903 137461
rect 151963 136676 152122 136678
rect 151963 136521 151965 136676
rect 151965 136521 152120 136676
rect 152120 136521 152122 136676
rect 151963 136519 152122 136521
rect -1003 135861 -903 135961
rect 151963 135176 152122 135178
rect 151963 135021 151965 135176
rect 151965 135021 152120 135176
rect 152120 135021 152122 135176
rect 151963 135019 152122 135021
rect -1003 134361 -903 134461
rect 151963 133676 152122 133678
rect 151963 133521 151965 133676
rect 151965 133521 152120 133676
rect 152120 133521 152122 133676
rect 151963 133519 152122 133521
rect -1003 132861 -903 132961
rect 151963 132176 152122 132178
rect 151963 132021 151965 132176
rect 151965 132021 152120 132176
rect 152120 132021 152122 132176
rect 151963 132019 152122 132021
rect -1003 131361 -903 131461
rect 151963 130676 152122 130678
rect 151963 130521 151965 130676
rect 151965 130521 152120 130676
rect 152120 130521 152122 130676
rect 151963 130519 152122 130521
rect -1003 129861 -903 129961
rect 151963 129176 152122 129178
rect 151963 129021 151965 129176
rect 151965 129021 152120 129176
rect 152120 129021 152122 129176
rect 151963 129019 152122 129021
rect -1003 128361 -903 128461
rect 151963 127676 152122 127678
rect 151963 127521 151965 127676
rect 151965 127521 152120 127676
rect 152120 127521 152122 127676
rect 151963 127519 152122 127521
rect -1003 126861 -903 126961
rect 151963 126176 152122 126178
rect 151963 126021 151965 126176
rect 151965 126021 152120 126176
rect 152120 126021 152122 126176
rect 151963 126019 152122 126021
rect -1003 125361 -903 125461
rect 151963 124676 152122 124678
rect 151963 124521 151965 124676
rect 151965 124521 152120 124676
rect 152120 124521 152122 124676
rect 151963 124519 152122 124521
rect -1003 123861 -903 123961
rect 151963 123176 152122 123178
rect 151963 123021 151965 123176
rect 151965 123021 152120 123176
rect 152120 123021 152122 123176
rect 151963 123019 152122 123021
rect -1003 122361 -903 122461
rect 151963 121676 152122 121678
rect 151963 121521 151965 121676
rect 151965 121521 152120 121676
rect 152120 121521 152122 121676
rect 151963 121519 152122 121521
rect -1003 120861 -903 120961
rect 151963 120176 152122 120178
rect 151963 120021 151965 120176
rect 151965 120021 152120 120176
rect 152120 120021 152122 120176
rect 151963 120019 152122 120021
rect -1003 119361 -903 119461
rect 151963 118676 152122 118678
rect 151963 118521 151965 118676
rect 151965 118521 152120 118676
rect 152120 118521 152122 118676
rect 151963 118519 152122 118521
rect -1003 117861 -903 117961
rect 151963 117176 152122 117178
rect 151963 117021 151965 117176
rect 151965 117021 152120 117176
rect 152120 117021 152122 117176
rect 151963 117019 152122 117021
rect -1003 116361 -903 116461
rect 151963 115676 152122 115678
rect 151963 115521 151965 115676
rect 151965 115521 152120 115676
rect 152120 115521 152122 115676
rect 151963 115519 152122 115521
rect -1003 114861 -903 114961
rect 151963 114176 152122 114178
rect 151963 114021 151965 114176
rect 151965 114021 152120 114176
rect 152120 114021 152122 114176
rect 151963 114019 152122 114021
rect -1003 113361 -903 113461
rect 151963 112676 152122 112678
rect 151963 112521 151965 112676
rect 151965 112521 152120 112676
rect 152120 112521 152122 112676
rect 151963 112519 152122 112521
rect -1003 111861 -903 111961
rect 151963 111176 152122 111178
rect 151963 111021 151965 111176
rect 151965 111021 152120 111176
rect 152120 111021 152122 111176
rect 151963 111019 152122 111021
rect -1003 110361 -903 110461
rect 151963 109676 152122 109678
rect 151963 109521 151965 109676
rect 151965 109521 152120 109676
rect 152120 109521 152122 109676
rect 151963 109519 152122 109521
rect -1003 108861 -903 108961
rect 151963 108176 152122 108178
rect 151963 108021 151965 108176
rect 151965 108021 152120 108176
rect 152120 108021 152122 108176
rect 151963 108019 152122 108021
rect -1003 107361 -903 107461
rect 151963 106676 152122 106678
rect 151963 106521 151965 106676
rect 151965 106521 152120 106676
rect 152120 106521 152122 106676
rect 151963 106519 152122 106521
rect -1003 105861 -903 105961
rect 151963 105176 152122 105178
rect 151963 105021 151965 105176
rect 151965 105021 152120 105176
rect 152120 105021 152122 105176
rect 151963 105019 152122 105021
rect -1003 104361 -903 104461
rect 151963 103676 152122 103678
rect 151963 103521 151965 103676
rect 151965 103521 152120 103676
rect 152120 103521 152122 103676
rect 151963 103519 152122 103521
rect -1003 102861 -903 102961
rect 151963 102176 152122 102178
rect 151963 102021 151965 102176
rect 151965 102021 152120 102176
rect 152120 102021 152122 102176
rect 151963 102019 152122 102021
rect -1003 101361 -903 101461
rect 151963 100676 152122 100678
rect 151963 100521 151965 100676
rect 151965 100521 152120 100676
rect 152120 100521 152122 100676
rect 151963 100519 152122 100521
rect -1003 99861 -903 99961
rect 151963 99176 152122 99178
rect 151963 99021 151965 99176
rect 151965 99021 152120 99176
rect 152120 99021 152122 99176
rect 151963 99019 152122 99021
rect -1003 98361 -903 98461
rect 151963 97676 152122 97678
rect 151963 97521 151965 97676
rect 151965 97521 152120 97676
rect 152120 97521 152122 97676
rect 151963 97519 152122 97521
rect -1003 96861 -903 96961
rect 151963 96176 152122 96178
rect 151963 96021 151965 96176
rect 151965 96021 152120 96176
rect 152120 96021 152122 96176
rect 151963 96019 152122 96021
rect -1003 95361 -903 95461
rect 151963 94676 152122 94678
rect 151963 94521 151965 94676
rect 151965 94521 152120 94676
rect 152120 94521 152122 94676
rect 151963 94519 152122 94521
rect -1003 93861 -903 93961
rect 151963 93176 152122 93178
rect 151963 93021 151965 93176
rect 151965 93021 152120 93176
rect 152120 93021 152122 93176
rect 151963 93019 152122 93021
rect -1003 92361 -903 92461
rect 151963 91676 152122 91678
rect 151963 91521 151965 91676
rect 151965 91521 152120 91676
rect 152120 91521 152122 91676
rect 151963 91519 152122 91521
rect -1003 90861 -903 90961
rect 151963 90176 152122 90178
rect 151963 90021 151965 90176
rect 151965 90021 152120 90176
rect 152120 90021 152122 90176
rect 151963 90019 152122 90021
rect -1003 89361 -903 89461
rect 151963 88676 152122 88678
rect 151963 88521 151965 88676
rect 151965 88521 152120 88676
rect 152120 88521 152122 88676
rect 151963 88519 152122 88521
rect -1003 87861 -903 87961
rect 151963 87176 152122 87178
rect 151963 87021 151965 87176
rect 151965 87021 152120 87176
rect 152120 87021 152122 87176
rect 151963 87019 152122 87021
rect -1003 86361 -903 86461
rect 151963 85676 152122 85678
rect 151963 85521 151965 85676
rect 151965 85521 152120 85676
rect 152120 85521 152122 85676
rect 151963 85519 152122 85521
rect -1003 84861 -903 84961
rect 151963 84176 152122 84178
rect 151963 84021 151965 84176
rect 151965 84021 152120 84176
rect 152120 84021 152122 84176
rect 151963 84019 152122 84021
rect -1003 83361 -903 83461
rect 151963 82676 152122 82678
rect 151963 82521 151965 82676
rect 151965 82521 152120 82676
rect 152120 82521 152122 82676
rect 151963 82519 152122 82521
rect -1003 81861 -903 81961
rect 151963 81176 152122 81178
rect 151963 81021 151965 81176
rect 151965 81021 152120 81176
rect 152120 81021 152122 81176
rect 151963 81019 152122 81021
rect -1003 80361 -903 80461
rect 151963 79676 152122 79678
rect 151963 79521 151965 79676
rect 151965 79521 152120 79676
rect 152120 79521 152122 79676
rect 151963 79519 152122 79521
rect -1003 78861 -903 78961
rect 151963 78176 152122 78178
rect 151963 78021 151965 78176
rect 151965 78021 152120 78176
rect 152120 78021 152122 78176
rect 151963 78019 152122 78021
rect -1003 77361 -903 77461
rect 151963 76676 152122 76678
rect 151963 76521 151965 76676
rect 151965 76521 152120 76676
rect 152120 76521 152122 76676
rect 151963 76519 152122 76521
rect -1003 75861 -903 75961
rect 151963 75176 152122 75178
rect 151963 75021 151965 75176
rect 151965 75021 152120 75176
rect 152120 75021 152122 75176
rect 151963 75019 152122 75021
rect -1003 74361 -903 74461
rect 151963 73676 152122 73678
rect 151963 73521 151965 73676
rect 151965 73521 152120 73676
rect 152120 73521 152122 73676
rect 151963 73519 152122 73521
rect -1003 72861 -903 72961
rect 151963 72176 152122 72178
rect 151963 72021 151965 72176
rect 151965 72021 152120 72176
rect 152120 72021 152122 72176
rect 151963 72019 152122 72021
rect -1003 71361 -903 71461
rect 151963 70676 152122 70678
rect 151963 70521 151965 70676
rect 151965 70521 152120 70676
rect 152120 70521 152122 70676
rect 151963 70519 152122 70521
rect -1003 69861 -903 69961
rect 151963 69176 152122 69178
rect 151963 69021 151965 69176
rect 151965 69021 152120 69176
rect 152120 69021 152122 69176
rect 151963 69019 152122 69021
rect -1003 68361 -903 68461
rect 151963 67676 152122 67678
rect 151963 67521 151965 67676
rect 151965 67521 152120 67676
rect 152120 67521 152122 67676
rect 151963 67519 152122 67521
rect -1003 66861 -903 66961
rect 151963 66176 152122 66178
rect 151963 66021 151965 66176
rect 151965 66021 152120 66176
rect 152120 66021 152122 66176
rect 151963 66019 152122 66021
rect -1003 65361 -903 65461
rect 151963 64676 152122 64678
rect 151963 64521 151965 64676
rect 151965 64521 152120 64676
rect 152120 64521 152122 64676
rect 151963 64519 152122 64521
rect -1003 63861 -903 63961
rect 151963 63176 152122 63178
rect 151963 63021 151965 63176
rect 151965 63021 152120 63176
rect 152120 63021 152122 63176
rect 151963 63019 152122 63021
rect -1003 62361 -903 62461
rect 151963 61676 152122 61678
rect 151963 61521 151965 61676
rect 151965 61521 152120 61676
rect 152120 61521 152122 61676
rect 151963 61519 152122 61521
rect -1003 60861 -903 60961
rect 151963 60176 152122 60178
rect 151963 60021 151965 60176
rect 151965 60021 152120 60176
rect 152120 60021 152122 60176
rect 151963 60019 152122 60021
rect -1003 59361 -903 59461
rect 151963 58676 152122 58678
rect 151963 58521 151965 58676
rect 151965 58521 152120 58676
rect 152120 58521 152122 58676
rect 151963 58519 152122 58521
rect -1003 57861 -903 57961
rect 151963 57176 152122 57178
rect 151963 57021 151965 57176
rect 151965 57021 152120 57176
rect 152120 57021 152122 57176
rect 151963 57019 152122 57021
rect -1003 56361 -903 56461
rect 151963 55676 152122 55678
rect 151963 55521 151965 55676
rect 151965 55521 152120 55676
rect 152120 55521 152122 55676
rect 151963 55519 152122 55521
rect -1003 54861 -903 54961
rect 151963 54176 152122 54178
rect 151963 54021 151965 54176
rect 151965 54021 152120 54176
rect 152120 54021 152122 54176
rect 151963 54019 152122 54021
rect -1003 53361 -903 53461
rect 151963 52676 152122 52678
rect 151963 52521 151965 52676
rect 151965 52521 152120 52676
rect 152120 52521 152122 52676
rect 151963 52519 152122 52521
rect -1003 51861 -903 51961
rect 151963 51176 152122 51178
rect 151963 51021 151965 51176
rect 151965 51021 152120 51176
rect 152120 51021 152122 51176
rect 151963 51019 152122 51021
rect -1003 50361 -903 50461
rect 151963 49676 152122 49678
rect 151963 49521 151965 49676
rect 151965 49521 152120 49676
rect 152120 49521 152122 49676
rect 151963 49519 152122 49521
rect -1003 48861 -903 48961
rect 151963 48176 152122 48178
rect 151963 48021 151965 48176
rect 151965 48021 152120 48176
rect 152120 48021 152122 48176
rect 151963 48019 152122 48021
rect -1003 47361 -903 47461
rect 151963 46676 152122 46678
rect 151963 46521 151965 46676
rect 151965 46521 152120 46676
rect 152120 46521 152122 46676
rect 151963 46519 152122 46521
rect -1003 45861 -903 45961
rect 151963 45176 152122 45178
rect 151963 45021 151965 45176
rect 151965 45021 152120 45176
rect 152120 45021 152122 45176
rect 151963 45019 152122 45021
rect -1003 44361 -903 44461
rect 151963 43676 152122 43678
rect 151963 43521 151965 43676
rect 151965 43521 152120 43676
rect 152120 43521 152122 43676
rect 151963 43519 152122 43521
rect -1003 42861 -903 42961
rect 151963 42176 152122 42178
rect 151963 42021 151965 42176
rect 151965 42021 152120 42176
rect 152120 42021 152122 42176
rect 151963 42019 152122 42021
rect -1003 41361 -903 41461
rect 151963 40676 152122 40678
rect 151963 40521 151965 40676
rect 151965 40521 152120 40676
rect 152120 40521 152122 40676
rect 151963 40519 152122 40521
rect -1003 39861 -903 39961
rect 151963 39176 152122 39178
rect 151963 39021 151965 39176
rect 151965 39021 152120 39176
rect 152120 39021 152122 39176
rect 151963 39019 152122 39021
rect -1003 38361 -903 38461
rect 151963 37676 152122 37678
rect 151963 37521 151965 37676
rect 151965 37521 152120 37676
rect 152120 37521 152122 37676
rect 151963 37519 152122 37521
rect -1003 36861 -903 36961
rect 151963 36176 152122 36178
rect 151963 36021 151965 36176
rect 151965 36021 152120 36176
rect 152120 36021 152122 36176
rect 151963 36019 152122 36021
rect -1003 35361 -903 35461
rect 151963 34676 152122 34678
rect 151963 34521 151965 34676
rect 151965 34521 152120 34676
rect 152120 34521 152122 34676
rect 151963 34519 152122 34521
rect -1003 33861 -903 33961
rect 151963 33176 152122 33178
rect 151963 33021 151965 33176
rect 151965 33021 152120 33176
rect 152120 33021 152122 33176
rect 151963 33019 152122 33021
rect -1003 32361 -903 32461
rect 151963 31676 152122 31678
rect 151963 31521 151965 31676
rect 151965 31521 152120 31676
rect 152120 31521 152122 31676
rect 151963 31519 152122 31521
rect -1003 30861 -903 30961
rect 151963 30176 152122 30178
rect 151963 30021 151965 30176
rect 151965 30021 152120 30176
rect 152120 30021 152122 30176
rect 151963 30019 152122 30021
rect -1003 29361 -903 29461
rect 151963 28676 152122 28678
rect 151963 28521 151965 28676
rect 151965 28521 152120 28676
rect 152120 28521 152122 28676
rect 151963 28519 152122 28521
rect -1003 27861 -903 27961
rect 151963 27176 152122 27178
rect 151963 27021 151965 27176
rect 151965 27021 152120 27176
rect 152120 27021 152122 27176
rect 151963 27019 152122 27021
rect -1003 26361 -903 26461
rect 151963 25676 152122 25678
rect 151963 25521 151965 25676
rect 151965 25521 152120 25676
rect 152120 25521 152122 25676
rect 151963 25519 152122 25521
rect -1003 24861 -903 24961
rect 151963 24176 152122 24178
rect 151963 24021 151965 24176
rect 151965 24021 152120 24176
rect 152120 24021 152122 24176
rect 151963 24019 152122 24021
rect -1003 23361 -903 23461
rect 151963 22676 152122 22678
rect 151963 22521 151965 22676
rect 151965 22521 152120 22676
rect 152120 22521 152122 22676
rect 151963 22519 152122 22521
rect -1003 21861 -903 21961
rect 151963 21176 152122 21178
rect 151963 21021 151965 21176
rect 151965 21021 152120 21176
rect 152120 21021 152122 21176
rect 151963 21019 152122 21021
rect -1003 20361 -903 20461
rect 151963 19676 152122 19678
rect 151963 19521 151965 19676
rect 151965 19521 152120 19676
rect 152120 19521 152122 19676
rect 151963 19519 152122 19521
rect -1003 18861 -903 18961
rect 151963 18176 152122 18178
rect 151963 18021 151965 18176
rect 151965 18021 152120 18176
rect 152120 18021 152122 18176
rect 151963 18019 152122 18021
rect -1003 17361 -903 17461
rect 151963 16676 152122 16678
rect 151963 16521 151965 16676
rect 151965 16521 152120 16676
rect 152120 16521 152122 16676
rect 151963 16519 152122 16521
rect -1003 15861 -903 15961
rect 151963 15176 152122 15178
rect 151963 15021 151965 15176
rect 151965 15021 152120 15176
rect 152120 15021 152122 15176
rect 151963 15019 152122 15021
rect -1003 14361 -903 14461
rect 151963 13676 152122 13678
rect 151963 13521 151965 13676
rect 151965 13521 152120 13676
rect 152120 13521 152122 13676
rect 151963 13519 152122 13521
rect -1003 12861 -903 12961
rect 151963 12176 152122 12178
rect 151963 12021 151965 12176
rect 151965 12021 152120 12176
rect 152120 12021 152122 12176
rect 151963 12019 152122 12021
rect -1003 11361 -903 11461
rect 151963 10676 152122 10678
rect 151963 10521 151965 10676
rect 151965 10521 152120 10676
rect 152120 10521 152122 10676
rect 151963 10519 152122 10521
rect 9935 9594 10044 9596
rect 9935 9489 9937 9594
rect 9937 9489 10042 9594
rect 10042 9489 10044 9594
rect 9935 9487 10044 9489
rect 1832 9377 1991 9379
rect 1832 9222 1834 9377
rect 1834 9222 1989 9377
rect 1989 9222 1991 9377
rect 1832 9220 1991 9222
rect 2664 9390 2773 9392
rect 2664 9285 2666 9390
rect 2666 9285 2771 9390
rect 2771 9285 2773 9390
rect 2664 9283 2773 9285
rect 3741 9443 3850 9445
rect 3741 9338 3743 9443
rect 3743 9338 3848 9443
rect 3848 9338 3850 9443
rect 3741 9336 3850 9338
rect 5356 9415 5465 9417
rect 5356 9310 5358 9415
rect 5358 9310 5463 9415
rect 5463 9310 5465 9415
rect 5356 9308 5465 9310
rect 6901 9462 7010 9464
rect 6901 9357 6903 9462
rect 6903 9357 7008 9462
rect 7008 9357 7010 9462
rect 6901 9355 7010 9357
rect 8456 9406 8565 9408
rect 8456 9301 8458 9406
rect 8458 9301 8563 9406
rect 8563 9301 8565 9406
rect 8456 9299 8565 9301
rect 12972 9503 13081 9505
rect 12972 9398 12974 9503
rect 12974 9398 13079 9503
rect 13079 9398 13081 9503
rect 12972 9396 13081 9398
rect 14542 9421 14651 9530
rect 16164 9491 16273 9493
rect 16164 9386 16166 9491
rect 16166 9386 16271 9491
rect 16271 9386 16273 9491
rect 16164 9384 16273 9386
rect 17664 9525 17773 9527
rect 17664 9420 17666 9525
rect 17666 9420 17771 9525
rect 17771 9420 17773 9525
rect 17664 9418 17773 9420
rect 19164 9607 19273 9609
rect 19164 9502 19166 9607
rect 19166 9502 19271 9607
rect 19271 9502 19273 9607
rect 19164 9500 19273 9502
rect 9044 9377 9203 9379
rect 9044 9222 9046 9377
rect 9046 9222 9201 9377
rect 9201 9222 9203 9377
rect 9044 9220 9203 9222
rect 11449 9327 11558 9329
rect 11449 9222 11451 9327
rect 11451 9222 11556 9327
rect 11556 9222 11558 9327
rect 11449 9220 11558 9222
rect 16457 9377 16616 9379
rect 16457 9222 16459 9377
rect 16459 9222 16614 9377
rect 16614 9222 16616 9377
rect 16457 9220 16616 9222
rect 20664 9434 20773 9436
rect 20664 9329 20666 9434
rect 20666 9329 20771 9434
rect 20771 9329 20773 9434
rect 20664 9327 20773 9329
rect 22164 9459 22273 9461
rect 22164 9354 22166 9459
rect 22166 9354 22271 9459
rect 22271 9354 22273 9459
rect 22164 9352 22273 9354
rect 23664 9563 23773 9565
rect 23664 9458 23666 9563
rect 23666 9458 23771 9563
rect 23771 9458 23773 9563
rect 23664 9456 23773 9458
rect 25258 9503 25367 9505
rect 25258 9398 25260 9503
rect 25260 9398 25365 9503
rect 25365 9398 25367 9503
rect 25258 9396 25367 9398
rect 26769 9519 26878 9521
rect 26769 9414 26771 9519
rect 26771 9414 26876 9519
rect 26876 9414 26878 9519
rect 26769 9412 26878 9414
rect 28308 9579 28417 9581
rect 28308 9474 28310 9579
rect 28310 9474 28415 9579
rect 28415 9474 28417 9579
rect 28308 9472 28417 9474
rect 29815 9431 29924 9433
rect 29815 9326 29817 9431
rect 29817 9326 29922 9431
rect 29922 9326 29924 9431
rect 29815 9324 29924 9326
rect 31316 9393 31425 9395
rect 31316 9288 31318 9393
rect 31318 9288 31423 9393
rect 31423 9288 31425 9393
rect 31316 9286 31425 9288
rect 32128 9377 32287 9379
rect 32128 9222 32130 9377
rect 32130 9222 32285 9377
rect 32285 9222 32287 9377
rect 32128 9220 32287 9222
rect 32871 9438 32980 9440
rect 32871 9333 32873 9438
rect 32873 9333 32978 9438
rect 32978 9333 32980 9438
rect 32871 9331 32980 9333
rect 34164 9367 34273 9476
rect 35964 9421 36073 9530
rect 37539 9513 37648 9515
rect 37539 9408 37541 9513
rect 37541 9408 37646 9513
rect 37646 9408 37648 9513
rect 37539 9406 37648 9408
rect 40595 9353 40704 9452
rect 40595 9343 40597 9353
rect 40597 9343 40702 9353
rect 40702 9343 40704 9353
rect 1164 9217 1273 9219
rect 1164 9112 1166 9217
rect 1166 9112 1271 9217
rect 1271 9112 1273 9217
rect 1164 9110 1273 9112
rect 45206 9416 45315 9418
rect 45206 9311 45208 9416
rect 45208 9311 45313 9416
rect 45313 9311 45315 9416
rect 45206 9309 45315 9311
rect 46778 9394 46887 9396
rect 46778 9289 46780 9394
rect 46780 9289 46885 9394
rect 46885 9289 46887 9394
rect 46778 9287 46887 9289
rect 48227 9435 48336 9437
rect 48227 9330 48229 9435
rect 48229 9330 48334 9435
rect 48334 9330 48336 9435
rect 48227 9328 48336 9330
rect 54451 9514 54560 9516
rect 54451 9409 54453 9514
rect 54453 9409 54558 9514
rect 54558 9409 54560 9514
rect 54451 9407 54560 9409
rect 51356 9368 51465 9370
rect 51356 9263 51358 9368
rect 51358 9263 51463 9368
rect 51463 9263 51465 9368
rect 51356 9261 51465 9263
rect 52838 9375 52947 9377
rect 52838 9270 52840 9375
rect 52840 9270 52945 9375
rect 52945 9270 52947 9375
rect 52838 9268 52947 9270
rect 55974 9465 56083 9467
rect 55974 9360 55976 9465
rect 55976 9360 56081 9465
rect 56081 9360 56083 9465
rect 55974 9358 56083 9360
rect 57477 9490 57586 9492
rect 57477 9385 57479 9490
rect 57479 9385 57584 9490
rect 57584 9385 57586 9490
rect 57477 9383 57586 9385
rect 58984 9486 59093 9488
rect 58984 9381 58986 9486
rect 58986 9381 59091 9486
rect 59091 9381 59093 9486
rect 58984 9379 59093 9381
rect 60575 9430 60684 9432
rect 60575 9325 60577 9430
rect 60577 9325 60682 9430
rect 60682 9325 60684 9430
rect 60575 9323 60684 9325
rect 39049 9044 39158 9153
rect -3102 8873 -3099 8971
rect -3099 8873 -2999 8971
rect -2999 8873 -2997 8971
rect 42137 9092 42246 9201
rect 43668 9155 43777 9157
rect 43668 9050 43670 9155
rect 43670 9050 43775 9155
rect 43775 9050 43777 9155
rect 43668 9048 43777 9050
rect 49799 9248 49908 9250
rect 49799 9143 49801 9248
rect 49801 9143 49906 9248
rect 49906 9143 49908 9248
rect 49799 9141 49908 9143
rect 60839 9377 60998 9379
rect 60839 9222 60841 9377
rect 60841 9222 60996 9377
rect 60996 9222 60998 9377
rect 60839 9220 60998 9222
rect 62059 9316 62168 9425
rect 63621 9469 63730 9471
rect 63621 9364 63623 9469
rect 63623 9364 63728 9469
rect 63728 9364 63730 9469
rect 63621 9362 63730 9364
rect 65125 9404 65234 9406
rect 65125 9299 65127 9404
rect 65127 9299 65232 9404
rect 65232 9299 65234 9404
rect 65125 9297 65234 9299
rect 66706 9324 66815 9433
rect 69776 9298 69885 9300
rect 69776 9193 69778 9298
rect 69778 9193 69883 9298
rect 69883 9193 69885 9298
rect 69776 9191 69885 9193
rect 71300 9332 71409 9334
rect 71300 9227 71302 9332
rect 71302 9227 71407 9332
rect 71407 9227 71409 9332
rect 71300 9225 71409 9227
rect 72789 9419 72898 9421
rect 72789 9314 72791 9419
rect 72791 9314 72896 9419
rect 72896 9314 72898 9419
rect 72789 9312 72898 9314
rect 74377 9419 74486 9421
rect 74377 9314 74379 9419
rect 74379 9314 74484 9419
rect 74484 9314 74486 9419
rect 74377 9312 74486 9314
rect 75886 9385 75995 9387
rect 75886 9280 75888 9385
rect 75888 9280 75993 9385
rect 75993 9280 75995 9385
rect 75886 9278 75995 9280
rect 77396 9427 77505 9429
rect 77396 9322 77398 9427
rect 77398 9322 77503 9427
rect 77503 9322 77505 9427
rect 77396 9320 77505 9322
rect 78922 9496 79031 9498
rect 78922 9391 78924 9496
rect 78924 9391 79029 9496
rect 79029 9391 79031 9496
rect 78922 9389 79031 9391
rect 87183 9565 87292 9567
rect 87183 9460 87185 9565
rect 87185 9460 87290 9565
rect 87290 9460 87292 9565
rect 87183 9458 87292 9460
rect 80443 9377 80552 9379
rect 80443 9272 80445 9377
rect 80445 9272 80550 9377
rect 80550 9272 80552 9377
rect 80443 9270 80552 9272
rect 81619 9227 81728 9229
rect 81619 9122 81621 9227
rect 81621 9122 81726 9227
rect 81726 9122 81728 9227
rect 81619 9120 81728 9122
rect 83774 9377 83933 9379
rect 83774 9222 83776 9377
rect 83776 9222 83931 9377
rect 83931 9222 83933 9377
rect 83774 9220 83933 9222
rect 88164 9404 88273 9406
rect 88164 9299 88166 9404
rect 88166 9299 88271 9404
rect 88271 9299 88273 9404
rect 88164 9297 88273 9299
rect 86541 9242 86650 9244
rect 86541 9137 86543 9242
rect 86543 9137 86648 9242
rect 86648 9137 86650 9242
rect 86541 9135 86650 9137
rect 90274 9377 90433 9379
rect 90274 9222 90276 9377
rect 90276 9222 90431 9377
rect 90431 9222 90433 9377
rect 90274 9220 90433 9222
rect 94774 9377 94933 9379
rect 94774 9222 94776 9377
rect 94776 9222 94931 9377
rect 94931 9222 94933 9377
rect 94774 9220 94933 9222
rect 99274 9377 99433 9379
rect 99274 9222 99276 9377
rect 99276 9222 99431 9377
rect 99431 9222 99433 9377
rect 99274 9220 99433 9222
rect 102274 9377 102433 9379
rect 102274 9222 102276 9377
rect 102276 9222 102431 9377
rect 102431 9222 102433 9377
rect 102274 9220 102433 9222
rect 68234 9118 68343 9120
rect 68234 9013 68236 9118
rect 68236 9013 68341 9118
rect 68341 9013 68343 9118
rect 68234 9011 68343 9013
rect 103164 9225 103273 9227
rect 103164 9120 103166 9225
rect 103166 9120 103271 9225
rect 103271 9120 103273 9225
rect 103164 9118 103273 9120
rect 105774 9377 105933 9379
rect 105774 9222 105776 9377
rect 105776 9222 105931 9377
rect 105931 9222 105933 9377
rect 105774 9220 105933 9222
rect 107664 9279 107773 9281
rect 107664 9174 107666 9279
rect 107666 9174 107771 9279
rect 107771 9174 107773 9279
rect 107664 9172 107773 9174
rect 111774 9377 111933 9379
rect 111774 9222 111776 9377
rect 111776 9222 111931 9377
rect 111931 9222 111933 9377
rect 111774 9220 111933 9222
rect 114829 9467 114938 9469
rect 114829 9362 114831 9467
rect 114831 9362 114936 9467
rect 114936 9362 114938 9467
rect 114829 9360 114938 9362
rect 116274 9377 116433 9379
rect 116274 9222 116276 9377
rect 116276 9222 116431 9377
rect 116431 9222 116433 9377
rect 116274 9220 116433 9222
rect 116664 9342 116773 9344
rect 116664 9237 116666 9342
rect 116666 9237 116771 9342
rect 116771 9237 116773 9342
rect 116664 9235 116773 9237
rect 119274 9377 119433 9379
rect 119274 9222 119276 9377
rect 119276 9222 119431 9377
rect 119431 9222 119433 9377
rect 119274 9220 119433 9222
rect 113597 9212 113706 9214
rect 113597 9107 113599 9212
rect 113599 9107 113704 9212
rect 113704 9107 113706 9212
rect 113597 9105 113706 9107
rect 120836 9265 120945 9267
rect 120836 9160 120838 9265
rect 120838 9160 120943 9265
rect 120943 9160 120945 9265
rect 120836 9158 120945 9160
rect 121164 9283 121273 9285
rect 121164 9178 121166 9283
rect 121166 9178 121271 9283
rect 121271 9178 121273 9283
rect 121164 9176 121273 9178
rect 125274 9377 125433 9379
rect 125274 9222 125276 9377
rect 125276 9222 125431 9377
rect 125431 9222 125433 9377
rect 125274 9220 125433 9222
rect 82964 9085 83073 9087
rect 82964 8980 82966 9085
rect 82966 8980 83071 9085
rect 83071 8980 83073 9085
rect 82964 8978 83073 8980
rect -3102 8871 -2997 8873
rect 91237 8927 91346 8929
rect 91237 8822 91239 8927
rect 91239 8822 91344 8927
rect 91344 8822 91346 8927
rect 91237 8820 91346 8822
rect 92664 9016 92773 9018
rect 92664 8911 92666 9016
rect 92666 8911 92771 9016
rect 92771 8911 92773 9016
rect 92664 8909 92773 8911
rect 98397 8962 98506 8964
rect 98397 8857 98399 8962
rect 98399 8857 98504 8962
rect 98504 8857 98506 8962
rect 98397 8855 98506 8857
rect 100458 8976 100567 8978
rect 100458 8871 100460 8976
rect 100460 8871 100565 8976
rect 100565 8871 100567 8976
rect 100458 8869 100567 8871
rect 106578 9047 106687 9049
rect 106578 8942 106580 9047
rect 106580 8942 106685 9047
rect 106685 8942 106687 9047
rect 106578 8940 106687 8942
rect 117325 9149 117434 9151
rect 117325 9044 117327 9149
rect 117327 9044 117432 9149
rect 117432 9044 117434 9149
rect 117325 9042 117434 9044
rect 126963 9252 127072 9254
rect 126963 9147 126965 9252
rect 126965 9147 127070 9252
rect 127070 9147 127072 9252
rect 126963 9145 127072 9147
rect 127164 9348 127273 9350
rect 127164 9243 127166 9348
rect 127166 9243 127271 9348
rect 127271 9243 127273 9348
rect 127164 9241 127273 9243
rect 131974 9377 132133 9379
rect 131974 9222 131976 9377
rect 131976 9222 132131 9377
rect 132131 9222 132133 9377
rect 131974 9220 132133 9222
rect 134516 9278 134625 9280
rect 134516 9173 134518 9278
rect 134518 9173 134623 9278
rect 134623 9173 134625 9278
rect 134516 9171 134625 9173
rect 134974 9377 135133 9379
rect 134974 9222 134976 9377
rect 134976 9222 135131 9377
rect 135131 9222 135133 9377
rect 134974 9220 135133 9222
rect 136474 9377 136633 9379
rect 136474 9222 136476 9377
rect 136476 9222 136631 9377
rect 136631 9222 136633 9377
rect 136474 9220 136633 9222
rect 137974 9377 138133 9379
rect 137974 9222 137976 9377
rect 137976 9222 138131 9377
rect 138131 9222 138133 9377
rect 137974 9220 138133 9222
rect 139838 9347 139947 9349
rect 139838 9242 139840 9347
rect 139840 9242 139945 9347
rect 139945 9242 139947 9347
rect 139838 9240 139947 9242
rect 140974 9377 141133 9379
rect 140974 9222 140976 9377
rect 140976 9222 141131 9377
rect 141131 9222 141133 9377
rect 140974 9220 141133 9222
rect 142974 9377 143133 9379
rect 142974 9222 142976 9377
rect 142976 9222 143131 9377
rect 143131 9222 143133 9377
rect 142974 9220 143133 9222
rect 145164 9475 145273 9477
rect 145164 9370 145166 9475
rect 145166 9370 145271 9475
rect 145271 9370 145273 9475
rect 145164 9368 145273 9370
rect 152693 9547 152802 9549
rect 152693 9442 152695 9547
rect 152695 9442 152800 9547
rect 152800 9442 152802 9547
rect 152693 9440 152802 9442
rect 146974 9377 147133 9379
rect 146974 9222 146976 9377
rect 146976 9222 147131 9377
rect 147131 9222 147133 9377
rect 146974 9220 147133 9222
rect 148474 9377 148633 9379
rect 148474 9222 148476 9377
rect 148476 9222 148631 9377
rect 148631 9222 148633 9377
rect 148474 9220 148633 9222
rect 149974 9377 150133 9379
rect 149974 9222 149976 9377
rect 149976 9222 150131 9377
rect 150131 9222 150133 9377
rect 149974 9220 150133 9222
rect 151474 9377 151633 9379
rect 151474 9222 151476 9377
rect 151476 9222 151631 9377
rect 151631 9222 151633 9377
rect 151474 9220 151633 9222
rect 120458 9005 120567 9007
rect 120458 8900 120460 9005
rect 120460 8900 120565 9005
rect 120565 8900 120567 9005
rect 120458 8898 120567 8900
rect 130522 9060 130631 9062
rect 130522 8955 130524 9060
rect 130524 8955 130629 9060
rect 130629 8955 130631 9060
rect 130522 8953 130631 8955
rect 134664 9132 134773 9134
rect 134664 9027 134666 9132
rect 134666 9027 134771 9132
rect 134771 9027 134773 9132
rect 134664 9025 134773 9027
rect 139439 9101 139548 9103
rect 139439 8996 139441 9101
rect 139441 8996 139546 9101
rect 139546 8996 139548 9101
rect 139439 8994 139548 8996
rect 94164 8827 94273 8829
rect 94164 8722 94166 8827
rect 94166 8722 94271 8827
rect 94271 8722 94273 8827
rect 94164 8720 94273 8722
rect 103500 8873 103609 8875
rect 103500 8768 103502 8873
rect 103502 8768 103607 8873
rect 103607 8768 103609 8873
rect 103500 8766 103609 8768
rect 110664 8853 110773 8855
rect 110664 8748 110666 8853
rect 110666 8748 110771 8853
rect 110771 8748 110773 8853
rect 110664 8746 110773 8748
rect 124834 8928 124943 8930
rect 124834 8823 124836 8928
rect 124836 8823 124941 8928
rect 124941 8823 124943 8928
rect 124834 8821 124943 8823
rect 132935 8979 133044 8981
rect 132935 8874 132937 8979
rect 132937 8874 133042 8979
rect 133042 8874 133044 8979
rect 132935 8872 133044 8874
rect 142164 9066 142273 9068
rect 142164 8961 142166 9066
rect 142166 8961 142271 9066
rect 142271 8961 142273 9066
rect 142164 8959 142273 8961
rect 146204 9111 146313 9113
rect 146204 9006 146206 9111
rect 146206 9006 146311 9111
rect 146311 9006 146313 9111
rect 146204 9004 146313 9006
rect 84432 8708 84541 8710
rect 84432 8603 84434 8708
rect 84434 8603 84539 8708
rect 84539 8603 84541 8708
rect 84432 8601 84541 8603
rect 138847 8789 138956 8791
rect 138847 8684 138849 8789
rect 138849 8684 138954 8789
rect 138954 8684 138956 8789
rect 138847 8682 138956 8684
rect 143465 8754 143574 8756
rect 143465 8649 143467 8754
rect 143467 8649 143572 8754
rect 143572 8649 143574 8754
rect 143465 8647 143574 8649
rect 149629 8859 149738 8861
rect 149629 8754 149631 8859
rect 149631 8754 149736 8859
rect 149736 8754 149738 8859
rect 149629 8752 149738 8754
rect 92005 8574 92114 8576
rect 92005 8469 92007 8574
rect 92007 8469 92112 8574
rect 92112 8469 92114 8574
rect 92005 8467 92114 8469
rect 106952 8632 107061 8634
rect 106952 8527 106954 8632
rect 106954 8527 107059 8632
rect 107059 8527 107061 8632
rect 106952 8525 107061 8527
rect 96733 8507 96842 8509
rect 96733 8402 96735 8507
rect 96735 8402 96840 8507
rect 96840 8402 96842 8507
rect 96733 8400 96842 8402
rect 110344 8612 110453 8614
rect 110344 8507 110346 8612
rect 110346 8507 110451 8612
rect 110451 8507 110453 8612
rect 110344 8505 110453 8507
rect 101002 8445 101111 8447
rect 101002 8340 101004 8445
rect 101004 8340 101109 8445
rect 101109 8340 101111 8445
rect 101002 8338 101111 8340
rect 124356 8536 124465 8538
rect 124356 8431 124358 8536
rect 124358 8431 124463 8536
rect 124463 8431 124465 8536
rect 124356 8429 124465 8431
rect 130027 8621 130136 8623
rect 130027 8516 130029 8621
rect 130029 8516 130134 8621
rect 130134 8516 130136 8621
rect 130027 8514 130136 8516
rect 150126 8550 150235 8552
rect 150126 8445 150128 8550
rect 150128 8445 150233 8550
rect 150233 8445 150235 8550
rect 150126 8443 150235 8445
rect 151471 8047 151473 8205
rect 151473 8047 151634 8205
rect 151634 8047 151637 8205
rect 151471 8044 151637 8047
rect 51 7694 54 7791
rect 54 7694 154 7791
rect 154 7694 156 7791
rect 51 7691 156 7694
rect 1829 7687 1832 7844
rect 1832 7687 1992 7844
rect 1992 7687 1994 7844
rect 9041 7696 9044 7853
rect 9044 7696 9204 7853
rect 9204 7696 9206 7853
rect 9041 7693 9206 7696
rect 1829 7684 1994 7687
rect 16454 7684 16457 7841
rect 16457 7684 16617 7841
rect 16617 7684 16619 7841
rect 16454 7681 16619 7684
rect 32125 7688 32128 7845
rect 32128 7688 32288 7845
rect 32288 7688 32290 7845
rect 60836 7695 60839 7852
rect 60839 7695 60999 7852
rect 60999 7695 61001 7852
rect 60836 7692 61001 7695
rect 83771 7696 83774 7853
rect 83774 7696 83934 7853
rect 83934 7696 83936 7853
rect 83771 7693 83936 7696
rect 90271 7696 90274 7853
rect 90274 7696 90434 7853
rect 90434 7696 90436 7853
rect 90271 7693 90436 7696
rect 94771 7696 94774 7853
rect 94774 7696 94934 7853
rect 94934 7696 94936 7853
rect 94771 7693 94936 7696
rect 99271 7696 99274 7853
rect 99274 7696 99434 7853
rect 99434 7696 99436 7853
rect 99271 7693 99436 7696
rect 102271 7696 102274 7853
rect 102274 7696 102434 7853
rect 102434 7696 102436 7853
rect 102271 7693 102436 7696
rect 105771 7696 105774 7853
rect 105774 7696 105934 7853
rect 105934 7696 105936 7853
rect 105771 7693 105936 7696
rect 111771 7696 111774 7853
rect 111774 7696 111934 7853
rect 111934 7696 111936 7853
rect 111771 7693 111936 7696
rect 116271 7696 116274 7853
rect 116274 7696 116434 7853
rect 116434 7696 116436 7853
rect 116271 7693 116436 7696
rect 119271 7696 119274 7853
rect 119274 7696 119434 7853
rect 119434 7696 119436 7853
rect 119271 7693 119436 7696
rect 125271 7696 125274 7853
rect 125274 7696 125434 7853
rect 125434 7696 125436 7853
rect 125271 7693 125436 7696
rect 131971 7696 131974 7853
rect 131974 7696 132134 7853
rect 132134 7696 132136 7853
rect 131971 7693 132136 7696
rect 134971 7696 134974 7853
rect 134974 7696 135134 7853
rect 135134 7696 135136 7853
rect 134971 7693 135136 7696
rect 136471 7696 136474 7853
rect 136474 7696 136634 7853
rect 136634 7696 136636 7853
rect 136471 7693 136636 7696
rect 137971 7696 137974 7853
rect 137974 7696 138134 7853
rect 138134 7696 138136 7853
rect 137971 7693 138136 7696
rect 140971 7696 140974 7853
rect 140974 7696 141134 7853
rect 141134 7696 141136 7853
rect 140971 7693 141136 7696
rect 142971 7696 142974 7853
rect 142974 7696 143134 7853
rect 143134 7696 143136 7853
rect 142971 7693 143136 7696
rect 146971 7696 146974 7853
rect 146974 7696 147134 7853
rect 147134 7696 147136 7853
rect 146971 7693 147136 7696
rect 148471 7696 148474 7853
rect 148474 7696 148634 7853
rect 148634 7696 148636 7853
rect 148471 7693 148636 7696
rect 149971 7696 149974 7853
rect 149974 7696 150134 7853
rect 150134 7696 150136 7853
rect 149971 7693 150136 7696
rect 151471 7696 151474 7853
rect 151474 7696 151634 7853
rect 151634 7696 151636 7853
rect 151471 7693 151636 7696
rect 32125 7685 32290 7688
<< metal4 >>
rect -3798 162933 -381 162988
rect -2601 161026 -603 161038
rect -2601 160890 -751 161026
rect -615 160890 -603 161026
rect -2601 160880 -603 160890
rect -2601 160878 -763 160880
rect -436 160464 -381 162933
rect 151963 160678 152123 160679
rect 151963 160519 151963 160678
rect 152122 160519 152123 160678
rect 151963 160519 152123 160519
rect -2987 159900 -1881 160060
rect -1003 159961 -902 159961
rect -1337 159861 -1003 159961
rect -903 159861 -902 159961
rect -1003 159860 -902 159861
rect -2601 159526 -603 159538
rect -2601 159390 -751 159526
rect -615 159390 -603 159526
rect -2601 159380 -603 159390
rect -2601 159378 -763 159380
rect 151963 159178 152123 159179
rect 151963 159019 151963 159178
rect 152122 159019 152123 159178
rect 151963 159019 152123 159019
rect -2987 158400 -1881 158560
rect -1003 158461 -902 158461
rect -1337 158361 -1003 158461
rect -903 158361 -902 158461
rect -1003 158360 -902 158361
rect -2601 158026 -603 158038
rect -2601 157890 -751 158026
rect -615 157890 -603 158026
rect -2601 157880 -603 157890
rect -2601 157878 -763 157880
rect 151963 157678 152123 157679
rect 151963 157519 151963 157678
rect 152122 157519 152123 157678
rect 151963 157519 152123 157519
rect -2987 156900 -1881 157060
rect -1003 156961 -902 156961
rect -1337 156861 -1003 156961
rect -903 156861 -902 156961
rect -1003 156860 -902 156861
rect -2601 156526 -603 156538
rect -2601 156390 -751 156526
rect -615 156390 -603 156526
rect -2601 156380 -603 156390
rect -2601 156378 -763 156380
rect 151963 156178 152123 156179
rect 151963 156019 151963 156178
rect 152122 156019 152123 156178
rect 151963 156019 152123 156019
rect -2987 155400 -1881 155560
rect -1003 155461 -902 155461
rect -1337 155361 -1003 155461
rect -903 155361 -902 155461
rect -1003 155360 -902 155361
rect -2601 155026 -603 155038
rect -2601 154890 -751 155026
rect -615 154890 -603 155026
rect -2601 154880 -603 154890
rect -2601 154878 -763 154880
rect 151963 154678 152123 154679
rect 151963 154519 151963 154678
rect 152122 154519 152123 154678
rect 151963 154519 152123 154519
rect -2987 153900 -1881 154060
rect -1003 153961 -902 153961
rect -1337 153861 -1003 153961
rect -903 153861 -902 153961
rect -1003 153860 -902 153861
rect -2601 153526 -603 153538
rect -2601 153390 -751 153526
rect -615 153390 -603 153526
rect -2601 153380 -603 153390
rect -2601 153378 -763 153380
rect 151963 153178 152123 153179
rect 151963 153019 151963 153178
rect 152122 153019 152123 153178
rect 151963 153019 152123 153019
rect -2987 152400 -1881 152560
rect -1003 152461 -902 152461
rect -1337 152361 -1003 152461
rect -903 152361 -902 152461
rect -1003 152360 -902 152361
rect -2601 152026 -603 152038
rect -2601 151890 -751 152026
rect -615 151890 -603 152026
rect -2601 151880 -603 151890
rect -2601 151878 -763 151880
rect 151963 151678 152123 151679
rect 151963 151519 151963 151678
rect 152122 151519 152123 151678
rect 151963 151519 152123 151519
rect -2987 150900 -1881 151060
rect -1003 150961 -902 150961
rect -1337 150861 -1003 150961
rect -903 150861 -902 150961
rect -1003 150860 -902 150861
rect -2601 150526 -603 150538
rect -2601 150390 -751 150526
rect -615 150390 -603 150526
rect -2601 150380 -603 150390
rect -2601 150378 -763 150380
rect 151963 150178 152123 150179
rect 151963 150019 151963 150178
rect 152122 150019 152123 150178
rect 151963 150019 152123 150019
rect -2987 149400 -1881 149560
rect -1003 149461 -902 149461
rect -1337 149361 -1003 149461
rect -903 149361 -902 149461
rect -1003 149360 -902 149361
rect -2601 149026 -603 149038
rect -2601 148890 -751 149026
rect -615 148890 -603 149026
rect -2601 148880 -603 148890
rect -2601 148878 -763 148880
rect 151963 148678 152123 148679
rect 151963 148519 151963 148678
rect 152122 148519 152123 148678
rect 151963 148519 152123 148519
rect -2987 147900 -1881 148060
rect -1003 147961 -902 147961
rect -1337 147861 -1003 147961
rect -903 147861 -902 147961
rect -1003 147860 -902 147861
rect -2601 147526 -603 147538
rect -2601 147390 -751 147526
rect -615 147390 -603 147526
rect -2601 147380 -603 147390
rect -2601 147378 -763 147380
rect 151963 147178 152123 147179
rect 151963 147019 151963 147178
rect 152122 147019 152123 147178
rect 151963 147019 152123 147019
rect -2987 146400 -1881 146560
rect -1003 146461 -902 146461
rect -1337 146361 -1003 146461
rect -903 146361 -902 146461
rect -1003 146360 -902 146361
rect -2601 146026 -603 146038
rect -2601 145890 -751 146026
rect -615 145890 -603 146026
rect -2601 145880 -603 145890
rect -2601 145878 -763 145880
rect 151963 145678 152123 145679
rect 151963 145519 151963 145678
rect 152122 145519 152123 145678
rect 151963 145519 152123 145519
rect -2987 144900 -1881 145060
rect -1003 144961 -902 144961
rect -1337 144861 -1003 144961
rect -903 144861 -902 144961
rect -1003 144860 -902 144861
rect -2601 144526 -603 144538
rect -2601 144390 -751 144526
rect -615 144390 -603 144526
rect -2601 144380 -603 144390
rect -2601 144378 -763 144380
rect 151963 144178 152123 144179
rect 151963 144019 151963 144178
rect 152122 144019 152123 144178
rect 151963 144019 152123 144019
rect -2987 143400 -1881 143560
rect -1003 143461 -902 143461
rect -1337 143361 -1003 143461
rect -903 143361 -902 143461
rect -1003 143360 -902 143361
rect -2601 143026 -603 143038
rect -2601 142890 -751 143026
rect -615 142890 -603 143026
rect -2601 142880 -603 142890
rect -2601 142878 -763 142880
rect 151963 142678 152123 142679
rect 151963 142519 151963 142678
rect 152122 142519 152123 142678
rect 151963 142519 152123 142519
rect -2987 141900 -1881 142060
rect -1003 141961 -902 141961
rect -1337 141861 -1003 141961
rect -903 141861 -902 141961
rect -1003 141860 -902 141861
rect -2601 141526 -603 141538
rect -2601 141390 -751 141526
rect -615 141390 -603 141526
rect -2601 141380 -603 141390
rect -2601 141378 -763 141380
rect 151963 141178 152123 141179
rect 151963 141019 151963 141178
rect 152122 141019 152123 141178
rect 151963 141019 152123 141019
rect -2987 140400 -1881 140560
rect -1003 140461 -902 140461
rect -1337 140361 -1003 140461
rect -903 140361 -902 140461
rect -1003 140360 -902 140361
rect -2601 140026 -603 140038
rect -2601 139890 -751 140026
rect -615 139890 -603 140026
rect -2601 139880 -603 139890
rect -2601 139878 -763 139880
rect 151963 139678 152123 139679
rect 151963 139519 151963 139678
rect 152122 139519 152123 139678
rect 151963 139519 152123 139519
rect -2987 138900 -1881 139060
rect -1003 138961 -902 138961
rect -1337 138861 -1003 138961
rect -903 138861 -902 138961
rect -1003 138860 -902 138861
rect -2601 138526 -603 138538
rect -2601 138390 -751 138526
rect -615 138390 -603 138526
rect -2601 138380 -603 138390
rect -2601 138378 -763 138380
rect 151963 138178 152123 138179
rect 151963 138019 151963 138178
rect 152122 138019 152123 138178
rect 151963 138019 152123 138019
rect -2987 137400 -1881 137560
rect -1003 137461 -902 137461
rect -1337 137361 -1003 137461
rect -903 137361 -902 137461
rect -1003 137360 -902 137361
rect -2601 137026 -603 137038
rect -2601 136890 -751 137026
rect -615 136890 -603 137026
rect -2601 136880 -603 136890
rect -2601 136878 -763 136880
rect 151963 136678 152123 136679
rect 151963 136519 151963 136678
rect 152122 136519 152123 136678
rect 151963 136519 152123 136519
rect -2987 135900 -1881 136060
rect -1003 135961 -902 135961
rect -1337 135861 -1003 135961
rect -903 135861 -902 135961
rect -1003 135860 -902 135861
rect -2601 135526 -603 135538
rect -2601 135390 -751 135526
rect -615 135390 -603 135526
rect -2601 135380 -603 135390
rect -2601 135378 -763 135380
rect 151963 135178 152123 135179
rect 151963 135019 151963 135178
rect 152122 135019 152123 135178
rect 151963 135019 152123 135019
rect -2987 134400 -1881 134560
rect -1003 134461 -902 134461
rect -1337 134361 -1003 134461
rect -903 134361 -902 134461
rect -1003 134360 -902 134361
rect -2601 134026 -603 134038
rect -2601 133890 -751 134026
rect -615 133890 -603 134026
rect -2601 133880 -603 133890
rect -2601 133878 -763 133880
rect 151963 133678 152123 133679
rect 151963 133519 151963 133678
rect 152122 133519 152123 133678
rect 151963 133519 152123 133519
rect -2987 132900 -1881 133060
rect -1003 132961 -902 132961
rect -1337 132861 -1003 132961
rect -903 132861 -902 132961
rect -1003 132860 -902 132861
rect -2601 132526 -603 132538
rect -2601 132390 -751 132526
rect -615 132390 -603 132526
rect -2601 132380 -603 132390
rect -2601 132378 -763 132380
rect 151963 132178 152123 132179
rect 151963 132019 151963 132178
rect 152122 132019 152123 132178
rect 151963 132019 152123 132019
rect -2987 131400 -1881 131560
rect -1003 131461 -902 131461
rect -1337 131361 -1003 131461
rect -903 131361 -902 131461
rect -1003 131360 -902 131361
rect -2601 131026 -603 131038
rect -2601 130890 -751 131026
rect -615 130890 -603 131026
rect -2601 130880 -603 130890
rect -2601 130878 -763 130880
rect 151963 130678 152123 130679
rect 151963 130519 151963 130678
rect 152122 130519 152123 130678
rect 151963 130519 152123 130519
rect -2987 129900 -1881 130060
rect -1003 129961 -902 129961
rect -1337 129861 -1003 129961
rect -903 129861 -902 129961
rect -1003 129860 -902 129861
rect -2601 129526 -603 129538
rect -2601 129390 -751 129526
rect -615 129390 -603 129526
rect -2601 129380 -603 129390
rect -2601 129378 -763 129380
rect 151963 129178 152123 129179
rect 151963 129019 151963 129178
rect 152122 129019 152123 129178
rect 151963 129019 152123 129019
rect -2987 128400 -1881 128560
rect -1003 128461 -902 128461
rect -1337 128361 -1003 128461
rect -903 128361 -902 128461
rect -1003 128360 -902 128361
rect -2601 128026 -603 128038
rect -2601 127890 -751 128026
rect -615 127890 -603 128026
rect -2601 127880 -603 127890
rect -2601 127878 -763 127880
rect 151963 127678 152123 127679
rect 151963 127519 151963 127678
rect 152122 127519 152123 127678
rect 151963 127519 152123 127519
rect -2987 126900 -1881 127060
rect -1003 126961 -902 126961
rect -1337 126861 -1003 126961
rect -903 126861 -902 126961
rect -1003 126860 -902 126861
rect -2601 126526 -603 126538
rect -2601 126390 -751 126526
rect -615 126390 -603 126526
rect -2601 126380 -603 126390
rect -2601 126378 -763 126380
rect 151963 126178 152123 126179
rect 151963 126019 151963 126178
rect 152122 126019 152123 126178
rect 151963 126019 152123 126019
rect -2987 125400 -1881 125560
rect -1003 125461 -902 125461
rect -1337 125361 -1003 125461
rect -903 125361 -902 125461
rect -1003 125360 -902 125361
rect -2601 125026 -603 125038
rect -2601 124890 -751 125026
rect -615 124890 -603 125026
rect -2601 124880 -603 124890
rect -2601 124878 -763 124880
rect 151963 124678 152123 124679
rect 151963 124519 151963 124678
rect 152122 124519 152123 124678
rect 151963 124519 152123 124519
rect -2987 123900 -1881 124060
rect -1003 123961 -902 123961
rect -1337 123861 -1003 123961
rect -903 123861 -902 123961
rect -1003 123860 -902 123861
rect 151963 123178 152123 123179
rect 151963 123019 151963 123178
rect 152122 123019 152123 123178
rect 151963 123019 152123 123019
rect -2987 122400 -1881 122560
rect -1003 122461 -902 122461
rect -1337 122361 -1003 122461
rect -903 122361 -902 122461
rect -1003 122360 -902 122361
rect -2601 122026 -603 122038
rect -2601 121890 -751 122026
rect -615 121890 -603 122026
rect -2601 121880 -603 121890
rect -2601 121878 -763 121880
rect 151963 121678 152123 121679
rect 151963 121519 151963 121678
rect 152122 121519 152123 121678
rect 151963 121519 152123 121519
rect -2987 120900 -1881 121060
rect -1003 120961 -902 120961
rect -1337 120861 -1003 120961
rect -903 120861 -902 120961
rect -1003 120860 -902 120861
rect -2601 120526 -603 120538
rect -2601 120390 -751 120526
rect -615 120390 -603 120526
rect -2601 120380 -603 120390
rect -2601 120378 -763 120380
rect 151963 120178 152123 120179
rect 151963 120019 151963 120178
rect 152122 120019 152123 120178
rect 151963 120019 152123 120019
rect -2987 119400 -1881 119560
rect -1003 119461 -902 119461
rect -1337 119361 -1003 119461
rect -903 119361 -902 119461
rect -1003 119360 -902 119361
rect -2601 119026 -603 119038
rect -2601 118890 -751 119026
rect -615 118890 -603 119026
rect -2601 118880 -603 118890
rect -2601 118878 -763 118880
rect 151963 118678 152123 118679
rect 151963 118519 151963 118678
rect 152122 118519 152123 118678
rect 151963 118519 152123 118519
rect -2987 117900 -1881 118060
rect -1003 117961 -902 117961
rect -1337 117861 -1003 117961
rect -903 117861 -902 117961
rect -1003 117860 -902 117861
rect -2601 117526 -603 117538
rect -2601 117390 -751 117526
rect -615 117390 -603 117526
rect -2601 117380 -603 117390
rect -2601 117378 -763 117380
rect 151963 117178 152123 117179
rect 151963 117019 151963 117178
rect 152122 117019 152123 117178
rect 151963 117019 152123 117019
rect -2987 116400 -1881 116560
rect -1003 116461 -902 116461
rect -1337 116361 -1003 116461
rect -903 116361 -902 116461
rect -1003 116360 -902 116361
rect -2601 116026 -603 116038
rect -2601 115890 -751 116026
rect -615 115890 -603 116026
rect -2601 115880 -603 115890
rect -2601 115878 -763 115880
rect 151963 115678 152123 115679
rect 151963 115519 151963 115678
rect 152122 115519 152123 115678
rect 151963 115519 152123 115519
rect -2987 114900 -1881 115060
rect -1003 114961 -902 114961
rect -1337 114861 -1003 114961
rect -903 114861 -902 114961
rect -1003 114860 -902 114861
rect -2601 114526 -603 114538
rect -2601 114390 -751 114526
rect -615 114390 -603 114526
rect -2601 114380 -603 114390
rect -2601 114378 -763 114380
rect 151963 114178 152123 114179
rect 151963 114019 151963 114178
rect 152122 114019 152123 114178
rect 151963 114019 152123 114019
rect -2987 113400 -1881 113560
rect -1003 113461 -902 113461
rect -1337 113361 -1003 113461
rect -903 113361 -902 113461
rect -1003 113360 -902 113361
rect -2601 113026 -603 113038
rect -2601 112890 -751 113026
rect -615 112890 -603 113026
rect -2601 112880 -603 112890
rect -2601 112878 -763 112880
rect 151963 112678 152123 112679
rect 151963 112519 151963 112678
rect 152122 112519 152123 112678
rect 151963 112519 152123 112519
rect -2987 111900 -1881 112060
rect -1003 111961 -902 111961
rect -1337 111861 -1003 111961
rect -903 111861 -902 111961
rect -1003 111860 -902 111861
rect -2601 111526 -603 111538
rect -2601 111390 -751 111526
rect -615 111390 -603 111526
rect -2601 111380 -603 111390
rect -2601 111378 -763 111380
rect 151963 111178 152123 111179
rect 151963 111019 151963 111178
rect 152122 111019 152123 111178
rect 151963 111019 152123 111019
rect -2987 110400 -1881 110560
rect -1003 110461 -902 110461
rect -1337 110361 -1003 110461
rect -903 110361 -902 110461
rect -1003 110360 -902 110361
rect -2601 110026 -603 110038
rect -2601 109890 -751 110026
rect -615 109890 -603 110026
rect -2601 109880 -603 109890
rect -2601 109878 -763 109880
rect 151963 109678 152123 109679
rect 151963 109519 151963 109678
rect 152122 109519 152123 109678
rect 151963 109519 152123 109519
rect -2987 108900 -1881 109060
rect -1003 108961 -902 108961
rect -1337 108861 -1003 108961
rect -903 108861 -902 108961
rect -1003 108860 -902 108861
rect -2601 108526 -603 108538
rect -2601 108390 -751 108526
rect -615 108390 -603 108526
rect -2601 108380 -603 108390
rect -2601 108378 -763 108380
rect 151963 108178 152123 108179
rect 151963 108019 151963 108178
rect 152122 108019 152123 108178
rect 151963 108019 152123 108019
rect -2987 107400 -1881 107560
rect -1003 107461 -902 107461
rect -1337 107361 -1003 107461
rect -903 107361 -902 107461
rect -1003 107360 -902 107361
rect -2601 107026 -603 107038
rect -2601 106890 -751 107026
rect -615 106890 -603 107026
rect -2601 106880 -603 106890
rect -2601 106878 -763 106880
rect 151963 106678 152123 106679
rect 151963 106519 151963 106678
rect 152122 106519 152123 106678
rect 151963 106519 152123 106519
rect -2987 105900 -1881 106060
rect -1003 105961 -902 105961
rect -1337 105861 -1003 105961
rect -903 105861 -902 105961
rect -1003 105860 -902 105861
rect -2601 105526 -603 105538
rect -2601 105390 -751 105526
rect -615 105390 -603 105526
rect -2601 105380 -603 105390
rect -2601 105378 -763 105380
rect 151963 105178 152123 105179
rect 151963 105019 151963 105178
rect 152122 105019 152123 105178
rect 151963 105019 152123 105019
rect -1003 104461 -902 104461
rect -1337 104361 -1003 104461
rect -903 104361 -902 104461
rect -1003 104360 -902 104361
rect -2601 104026 -603 104038
rect -2601 103890 -751 104026
rect -615 103890 -603 104026
rect -2601 103880 -603 103890
rect -2601 103878 -763 103880
rect 151963 103678 152123 103679
rect 151963 103519 151963 103678
rect 152122 103519 152123 103678
rect 151963 103519 152123 103519
rect -2987 102900 -1881 103060
rect -1003 102961 -902 102961
rect -1337 102861 -1003 102961
rect -903 102861 -902 102961
rect -1003 102860 -902 102861
rect -2601 102526 -603 102538
rect -2601 102390 -751 102526
rect -615 102390 -603 102526
rect -2601 102380 -603 102390
rect -2601 102378 -763 102380
rect 151963 102178 152123 102179
rect 151963 102019 151963 102178
rect 152122 102019 152123 102178
rect 151963 102019 152123 102019
rect -2987 101400 -1881 101560
rect -1003 101461 -902 101461
rect -1337 101361 -1003 101461
rect -903 101361 -902 101461
rect -1003 101360 -902 101361
rect -2601 101026 -603 101038
rect -2601 100890 -751 101026
rect -615 100890 -603 101026
rect -2601 100880 -603 100890
rect -2601 100878 -763 100880
rect 151963 100678 152123 100679
rect 151963 100519 151963 100678
rect 152122 100519 152123 100678
rect 151963 100519 152123 100519
rect -2987 99900 -1881 100060
rect -1003 99961 -902 99961
rect -1337 99861 -1003 99961
rect -903 99861 -902 99961
rect -1003 99860 -902 99861
rect -2601 99526 -603 99538
rect -2601 99390 -751 99526
rect -615 99390 -603 99526
rect -2601 99380 -603 99390
rect -2601 99378 -763 99380
rect 151963 99178 152123 99179
rect 151963 99019 151963 99178
rect 152122 99019 152123 99178
rect 151963 99019 152123 99019
rect -2987 98400 -1881 98560
rect -1003 98461 -902 98461
rect -1337 98361 -1003 98461
rect -903 98361 -902 98461
rect -1003 98360 -902 98361
rect -2601 98026 -603 98038
rect -2601 97890 -751 98026
rect -615 97890 -603 98026
rect -2601 97880 -603 97890
rect -2601 97878 -763 97880
rect 151963 97678 152123 97679
rect 151963 97519 151963 97678
rect 152122 97519 152123 97678
rect 151963 97519 152123 97519
rect -2987 96900 -1881 97060
rect -1003 96961 -902 96961
rect -1337 96861 -1003 96961
rect -903 96861 -902 96961
rect -1003 96860 -902 96861
rect -2601 96526 -603 96538
rect -2601 96390 -751 96526
rect -615 96390 -603 96526
rect -2601 96380 -603 96390
rect -2601 96378 -763 96380
rect 151963 96178 152123 96179
rect 151963 96019 151963 96178
rect 152122 96019 152123 96178
rect 151963 96019 152123 96019
rect -2987 95400 -1881 95560
rect -1003 95461 -902 95461
rect -1337 95361 -1003 95461
rect -903 95361 -902 95461
rect -1003 95360 -902 95361
rect -2601 95026 -603 95038
rect -2601 94890 -751 95026
rect -615 94890 -603 95026
rect -2601 94880 -603 94890
rect -2601 94878 -763 94880
rect 151963 94678 152123 94679
rect 151963 94519 151963 94678
rect 152122 94519 152123 94678
rect 151963 94519 152123 94519
rect -2987 93900 -1881 94060
rect -1003 93961 -902 93961
rect -1337 93861 -1003 93961
rect -903 93861 -902 93961
rect -1003 93860 -902 93861
rect -2601 93526 -603 93538
rect -2601 93390 -751 93526
rect -615 93390 -603 93526
rect -2601 93380 -603 93390
rect -2601 93378 -763 93380
rect 151963 93178 152123 93179
rect 151963 93019 151963 93178
rect 152122 93019 152123 93178
rect 151963 93019 152123 93019
rect -2987 92400 -1881 92560
rect -1003 92461 -902 92461
rect -1337 92361 -1003 92461
rect -903 92361 -902 92461
rect -1003 92360 -902 92361
rect -2601 92026 -603 92038
rect -2601 91890 -751 92026
rect -615 91890 -603 92026
rect -2601 91880 -603 91890
rect -2601 91878 -763 91880
rect 151963 91678 152123 91679
rect 151963 91519 151963 91678
rect 152122 91519 152123 91678
rect 151963 91519 152123 91519
rect -2987 90900 -1881 91060
rect -1003 90961 -902 90961
rect -1337 90861 -1003 90961
rect -903 90861 -902 90961
rect -1003 90860 -902 90861
rect -2601 90526 -603 90538
rect -2601 90390 -751 90526
rect -615 90390 -603 90526
rect -2601 90380 -603 90390
rect -2601 90378 -763 90380
rect 151963 90178 152123 90179
rect 151963 90019 151963 90178
rect 152122 90019 152123 90178
rect 151963 90019 152123 90019
rect -2987 89400 -1881 89560
rect -1003 89461 -902 89461
rect -1337 89361 -1003 89461
rect -903 89361 -902 89461
rect -1003 89360 -902 89361
rect -2601 89026 -603 89038
rect -2601 88890 -751 89026
rect -615 88890 -603 89026
rect -2601 88880 -603 88890
rect -2601 88878 -763 88880
rect 151963 88678 152123 88679
rect 151963 88519 151963 88678
rect 152122 88519 152123 88678
rect 151963 88519 152123 88519
rect -2987 87900 -1881 88060
rect -1003 87961 -902 87961
rect -1337 87861 -1003 87961
rect -903 87861 -902 87961
rect -1003 87860 -902 87861
rect -2601 87526 -603 87538
rect -2601 87390 -751 87526
rect -615 87390 -603 87526
rect -2601 87380 -603 87390
rect -2601 87378 -763 87380
rect 151963 87178 152123 87179
rect 151963 87019 151963 87178
rect 152122 87019 152123 87178
rect 151963 87019 152123 87019
rect -2987 86400 -1881 86560
rect -1003 86461 -902 86461
rect -1337 86361 -1003 86461
rect -903 86361 -902 86461
rect -1003 86360 -902 86361
rect -2601 86026 -603 86038
rect -2601 85890 -751 86026
rect -615 85890 -603 86026
rect -2601 85880 -603 85890
rect -2601 85878 -763 85880
rect 151963 85678 152123 85679
rect 151963 85519 151963 85678
rect 152122 85519 152123 85678
rect 151963 85519 152123 85519
rect -2987 84900 -1881 85060
rect -1003 84961 -902 84961
rect -1337 84861 -1003 84961
rect -903 84861 -902 84961
rect -1003 84860 -902 84861
rect -2601 84526 -603 84538
rect -2601 84390 -751 84526
rect -615 84390 -603 84526
rect -2601 84380 -603 84390
rect -2601 84378 -763 84380
rect 151963 84178 152123 84179
rect 151963 84019 151963 84178
rect 152122 84019 152123 84178
rect 151963 84019 152123 84019
rect -2987 83400 -1881 83560
rect -1003 83461 -902 83461
rect -1337 83361 -1003 83461
rect -903 83361 -902 83461
rect -1003 83360 -902 83361
rect -2601 83026 -603 83038
rect -2601 82890 -751 83026
rect -615 82890 -603 83026
rect -2601 82880 -603 82890
rect -2601 82878 -763 82880
rect 151963 82678 152123 82679
rect 151963 82519 151963 82678
rect 152122 82519 152123 82678
rect 151963 82519 152123 82519
rect -2987 81900 -1881 82060
rect -1003 81961 -902 81961
rect -1337 81861 -1003 81961
rect -903 81861 -902 81961
rect -1003 81860 -902 81861
rect -2601 81526 -603 81538
rect -2601 81390 -751 81526
rect -615 81390 -603 81526
rect -2601 81380 -603 81390
rect -2601 81378 -763 81380
rect 151963 81178 152123 81179
rect 151963 81019 151963 81178
rect 152122 81019 152123 81178
rect 151963 81019 152123 81019
rect -2987 80400 -1881 80560
rect -1003 80461 -902 80461
rect -1337 80361 -1003 80461
rect -903 80361 -902 80461
rect -1003 80360 -902 80361
rect -2601 80026 -603 80038
rect -2601 79890 -751 80026
rect -615 79890 -603 80026
rect -2601 79880 -603 79890
rect -2601 79878 -763 79880
rect 151963 79678 152123 79679
rect 151963 79519 151963 79678
rect 152122 79519 152123 79678
rect 151963 79519 152123 79519
rect -2987 78900 -1881 79060
rect -1003 78961 -902 78961
rect -1337 78861 -1003 78961
rect -903 78861 -902 78961
rect -1003 78860 -902 78861
rect -2601 78526 -603 78538
rect -2601 78390 -751 78526
rect -615 78390 -603 78526
rect -2601 78380 -603 78390
rect -2601 78378 -763 78380
rect 151963 78178 152123 78179
rect 151963 78019 151963 78178
rect 152122 78019 152123 78178
rect 151963 78019 152123 78019
rect -2987 77400 -1881 77560
rect -1003 77461 -902 77461
rect -1337 77361 -1003 77461
rect -903 77361 -902 77461
rect -1003 77360 -902 77361
rect -2601 77026 -603 77038
rect -2601 76890 -751 77026
rect -615 76890 -603 77026
rect -2601 76880 -603 76890
rect -2601 76878 -763 76880
rect 151963 76678 152123 76679
rect 151963 76519 151963 76678
rect 152122 76519 152123 76678
rect 151963 76519 152123 76519
rect -2987 75900 -1881 76060
rect -1003 75961 -902 75961
rect -1337 75861 -1003 75961
rect -903 75861 -902 75961
rect -1003 75860 -902 75861
rect -2601 75526 -603 75538
rect -2601 75390 -751 75526
rect -615 75390 -603 75526
rect -2601 75380 -603 75390
rect -2601 75378 -763 75380
rect 151963 75178 152123 75179
rect 151963 75019 151963 75178
rect 152122 75019 152123 75178
rect 151963 75019 152123 75019
rect -2987 74400 -1881 74560
rect -1003 74461 -902 74461
rect -1337 74361 -1003 74461
rect -903 74361 -902 74461
rect -1003 74360 -902 74361
rect -2601 74026 -603 74038
rect -2601 73890 -751 74026
rect -615 73890 -603 74026
rect -2601 73880 -603 73890
rect -2601 73878 -763 73880
rect 151963 73678 152123 73679
rect 151963 73519 151963 73678
rect 152122 73519 152123 73678
rect 151963 73519 152123 73519
rect -2987 72900 -1881 73060
rect -1003 72961 -902 72961
rect -1337 72861 -1003 72961
rect -903 72861 -902 72961
rect -1003 72860 -902 72861
rect -2601 72526 -603 72538
rect -2601 72390 -751 72526
rect -615 72390 -603 72526
rect -2601 72380 -603 72390
rect -2601 72378 -763 72380
rect 151963 72178 152123 72179
rect 151963 72019 151963 72178
rect 152122 72019 152123 72178
rect 151963 72019 152123 72019
rect -2987 71400 -1881 71560
rect -1003 71461 -902 71461
rect -1337 71361 -1003 71461
rect -903 71361 -902 71461
rect -1003 71360 -902 71361
rect -2601 71026 -603 71038
rect -2601 70890 -751 71026
rect -615 70890 -603 71026
rect -2601 70880 -603 70890
rect -2601 70878 -763 70880
rect 151963 70678 152123 70679
rect 151963 70519 151963 70678
rect 152122 70519 152123 70678
rect 151963 70519 152123 70519
rect -2987 69900 -1881 70060
rect -1003 69961 -902 69961
rect -1337 69861 -1003 69961
rect -903 69861 -902 69961
rect -1003 69860 -902 69861
rect -2601 69526 -603 69538
rect -2601 69390 -751 69526
rect -615 69390 -603 69526
rect -2601 69380 -603 69390
rect -2601 69378 -763 69380
rect 151963 69178 152123 69179
rect 151963 69019 151963 69178
rect 152122 69019 152123 69178
rect 151963 69019 152123 69019
rect -2987 68400 -1881 68560
rect -1003 68461 -902 68461
rect -1337 68361 -1003 68461
rect -903 68361 -902 68461
rect -1003 68360 -902 68361
rect -2601 68026 -603 68038
rect -2601 67890 -751 68026
rect -615 67890 -603 68026
rect -2601 67880 -603 67890
rect -2601 67878 -763 67880
rect 151963 67678 152123 67679
rect 151963 67519 151963 67678
rect 152122 67519 152123 67678
rect 151963 67519 152123 67519
rect -2987 66900 -1881 67060
rect -1003 66961 -902 66961
rect -1337 66861 -1003 66961
rect -903 66861 -902 66961
rect -1003 66860 -902 66861
rect -2601 66526 -603 66538
rect -2601 66390 -751 66526
rect -615 66390 -603 66526
rect -2601 66380 -603 66390
rect -2601 66378 -763 66380
rect 151963 66178 152123 66179
rect 151963 66019 151963 66178
rect 152122 66019 152123 66178
rect 151963 66019 152123 66019
rect -2987 65400 -1881 65560
rect -1003 65461 -902 65461
rect -1337 65361 -1003 65461
rect -903 65361 -902 65461
rect -1003 65360 -902 65361
rect -2601 65026 -603 65038
rect -2601 64890 -751 65026
rect -615 64890 -603 65026
rect -2601 64880 -603 64890
rect -2601 64878 -763 64880
rect 151963 64678 152123 64679
rect 151963 64519 151963 64678
rect 152122 64519 152123 64678
rect 151963 64519 152123 64519
rect -2987 63900 -1881 64060
rect -1003 63961 -902 63961
rect -1337 63861 -1003 63961
rect -903 63861 -902 63961
rect -1003 63860 -902 63861
rect -2601 63526 -603 63538
rect -2601 63390 -751 63526
rect -615 63390 -603 63526
rect -2601 63380 -603 63390
rect -2601 63378 -763 63380
rect 151963 63178 152123 63179
rect 151963 63019 151963 63178
rect 152122 63019 152123 63178
rect 151963 63019 152123 63019
rect -2987 62400 -1881 62560
rect -1003 62461 -902 62461
rect -1337 62361 -1003 62461
rect -903 62361 -902 62461
rect -1003 62360 -902 62361
rect -2601 62026 -603 62038
rect -2601 61890 -751 62026
rect -615 61890 -603 62026
rect -2601 61880 -603 61890
rect -2601 61878 -763 61880
rect 151963 61678 152123 61679
rect 151963 61519 151963 61678
rect 152122 61519 152123 61678
rect 151963 61519 152123 61519
rect -2987 60900 -1881 61060
rect -1003 60961 -902 60961
rect -1337 60861 -1003 60961
rect -903 60861 -902 60961
rect -1003 60860 -902 60861
rect -2601 60526 -603 60538
rect -2601 60390 -751 60526
rect -615 60390 -603 60526
rect -2601 60380 -603 60390
rect -2601 60378 -763 60380
rect 151963 60178 152123 60179
rect 151963 60019 151963 60178
rect 152122 60019 152123 60178
rect 151963 60019 152123 60019
rect -2987 59400 -1881 59560
rect -1003 59461 -902 59461
rect -1337 59361 -1003 59461
rect -903 59361 -902 59461
rect -1003 59360 -902 59361
rect -2601 59026 -603 59038
rect -2601 58890 -751 59026
rect -615 58890 -603 59026
rect -2601 58880 -603 58890
rect -2601 58878 -763 58880
rect 151963 58678 152123 58679
rect 151963 58519 151963 58678
rect 152122 58519 152123 58678
rect 151963 58519 152123 58519
rect -2987 57900 -1881 58060
rect -1003 57961 -902 57961
rect -1337 57861 -1003 57961
rect -903 57861 -902 57961
rect -1003 57860 -902 57861
rect -2601 57526 -603 57538
rect -2601 57390 -751 57526
rect -615 57390 -603 57526
rect -2601 57380 -603 57390
rect -2601 57378 -763 57380
rect 151963 57178 152123 57179
rect 151963 57019 151963 57178
rect 152122 57019 152123 57178
rect 151963 57019 152123 57019
rect -2987 56400 -1881 56560
rect -1003 56461 -902 56461
rect -1337 56361 -1003 56461
rect -903 56361 -902 56461
rect -1003 56360 -902 56361
rect -2601 56026 -603 56038
rect -2601 55890 -751 56026
rect -615 55890 -603 56026
rect -2601 55880 -603 55890
rect -2601 55878 -763 55880
rect 151963 55678 152123 55679
rect 151963 55519 151963 55678
rect 152122 55519 152123 55678
rect 151963 55519 152123 55519
rect -2987 54900 -1881 55060
rect -1003 54961 -902 54961
rect -1337 54861 -1003 54961
rect -903 54861 -902 54961
rect -1003 54860 -902 54861
rect -2601 54526 -603 54538
rect -2601 54390 -751 54526
rect -615 54390 -603 54526
rect -2601 54380 -603 54390
rect -2601 54378 -763 54380
rect 151963 54178 152123 54179
rect 151963 54019 151963 54178
rect 152122 54019 152123 54178
rect 151963 54019 152123 54019
rect -2987 53400 -1881 53560
rect -1003 53461 -902 53461
rect -1337 53361 -1003 53461
rect -903 53361 -902 53461
rect -1003 53360 -902 53361
rect -2601 53026 -603 53038
rect -2601 52890 -751 53026
rect -615 52890 -603 53026
rect -2601 52880 -603 52890
rect -2601 52878 -763 52880
rect 151963 52678 152123 52679
rect 151963 52519 151963 52678
rect 152122 52519 152123 52678
rect 151963 52519 152123 52519
rect -2987 51900 -1881 52060
rect -1003 51961 -902 51961
rect -1337 51861 -1003 51961
rect -903 51861 -902 51961
rect -1003 51860 -902 51861
rect -2601 51526 -603 51538
rect -2601 51390 -751 51526
rect -615 51390 -603 51526
rect -2601 51380 -603 51390
rect -2601 51378 -763 51380
rect 151963 51178 152123 51179
rect 151963 51019 151963 51178
rect 152122 51019 152123 51178
rect 151963 51019 152123 51019
rect -2987 50400 -1881 50560
rect -1003 50461 -902 50461
rect -1337 50361 -1003 50461
rect -903 50361 -902 50461
rect -1003 50360 -902 50361
rect -2601 50026 -603 50038
rect -2601 49890 -751 50026
rect -615 49890 -603 50026
rect -2601 49880 -603 49890
rect -2601 49878 -763 49880
rect 151963 49678 152123 49679
rect 151963 49519 151963 49678
rect 152122 49519 152123 49678
rect 151963 49519 152123 49519
rect -2987 48900 -1881 49060
rect -1003 48961 -902 48961
rect -1337 48861 -1003 48961
rect -903 48861 -902 48961
rect -1003 48860 -902 48861
rect -2601 48526 -603 48538
rect -2601 48390 -751 48526
rect -615 48390 -603 48526
rect -2601 48380 -603 48390
rect -2601 48378 -763 48380
rect 151963 48178 152123 48179
rect 151963 48019 151963 48178
rect 152122 48019 152123 48178
rect 151963 48019 152123 48019
rect -2987 47400 -1881 47560
rect -1003 47461 -902 47461
rect -1337 47361 -1003 47461
rect -903 47361 -902 47461
rect -1003 47360 -902 47361
rect 151963 46678 152123 46679
rect 151963 46519 151963 46678
rect 152122 46519 152123 46678
rect 151963 46519 152123 46519
rect -2987 45900 -1881 46060
rect -1003 45961 -902 45961
rect -1337 45861 -1003 45961
rect -903 45861 -902 45961
rect -1003 45860 -902 45861
rect -2601 45526 -603 45538
rect -2601 45390 -751 45526
rect -615 45390 -603 45526
rect -2601 45380 -603 45390
rect -2601 45378 -763 45380
rect 151963 45178 152123 45179
rect 151963 45019 151963 45178
rect 152122 45019 152123 45178
rect 151963 45019 152123 45019
rect -2987 44400 -1881 44560
rect -1003 44461 -902 44461
rect -1337 44361 -1003 44461
rect -903 44361 -902 44461
rect -1003 44360 -902 44361
rect -2601 44026 -603 44038
rect -2601 43890 -751 44026
rect -615 43890 -603 44026
rect -2601 43880 -603 43890
rect -2601 43878 -763 43880
rect 151963 43678 152123 43679
rect 151963 43519 151963 43678
rect 152122 43519 152123 43678
rect 151963 43519 152123 43519
rect -2987 42900 -1881 43060
rect -1003 42961 -902 42961
rect -1337 42861 -1003 42961
rect -903 42861 -902 42961
rect -1003 42860 -902 42861
rect -2601 42526 -603 42538
rect -2601 42390 -751 42526
rect -615 42390 -603 42526
rect -2601 42380 -603 42390
rect -2601 42378 -763 42380
rect 151963 42178 152123 42179
rect 151963 42019 151963 42178
rect 152122 42019 152123 42178
rect 151963 42019 152123 42019
rect -2987 41400 -1881 41560
rect -1003 41461 -902 41461
rect -1337 41361 -1003 41461
rect -903 41361 -902 41461
rect -1003 41360 -902 41361
rect -2601 41026 -603 41038
rect -2601 40890 -751 41026
rect -615 40890 -603 41026
rect -2601 40880 -603 40890
rect -2601 40878 -763 40880
rect 151963 40678 152123 40679
rect 151963 40519 151963 40678
rect 152122 40519 152123 40678
rect 151963 40519 152123 40519
rect -2987 39900 -1881 40060
rect -1003 39961 -902 39961
rect -1337 39861 -1003 39961
rect -903 39861 -902 39961
rect -1003 39860 -902 39861
rect -2601 39526 -603 39538
rect -2601 39390 -751 39526
rect -615 39390 -603 39526
rect -2601 39380 -603 39390
rect -2601 39378 -763 39380
rect 151963 39178 152123 39179
rect 151963 39019 151963 39178
rect 152122 39019 152123 39178
rect 151963 39019 152123 39019
rect -2987 38400 -1881 38560
rect -1003 38461 -902 38461
rect -1337 38361 -1003 38461
rect -903 38361 -902 38461
rect -1003 38360 -902 38361
rect -2601 38026 -603 38038
rect -2601 37890 -751 38026
rect -615 37890 -603 38026
rect -2601 37880 -603 37890
rect -2601 37878 -763 37880
rect 151963 37678 152123 37679
rect 151963 37519 151963 37678
rect 152122 37519 152123 37678
rect 151963 37519 152123 37519
rect -2987 36900 -1881 37060
rect -1003 36961 -902 36961
rect -1337 36861 -1003 36961
rect -903 36861 -902 36961
rect -1003 36860 -902 36861
rect -2601 36526 -603 36538
rect -2601 36390 -751 36526
rect -615 36390 -603 36526
rect -2601 36380 -603 36390
rect -2601 36378 -763 36380
rect 151963 36178 152123 36179
rect 151963 36019 151963 36178
rect 152122 36019 152123 36178
rect 151963 36019 152123 36019
rect -2987 35400 -1881 35560
rect -1003 35461 -902 35461
rect -1337 35361 -1003 35461
rect -903 35361 -902 35461
rect -1003 35360 -902 35361
rect -2601 35026 -603 35038
rect -2601 34890 -751 35026
rect -615 34890 -603 35026
rect -2601 34880 -603 34890
rect -2601 34878 -763 34880
rect 151963 34678 152123 34679
rect 151963 34519 151963 34678
rect 152122 34519 152123 34678
rect 151963 34519 152123 34519
rect -2987 33900 -1881 34060
rect -1003 33961 -902 33961
rect -1337 33861 -1003 33961
rect -903 33861 -902 33961
rect -1003 33860 -902 33861
rect -2601 33526 -603 33538
rect -2601 33390 -751 33526
rect -615 33390 -603 33526
rect -2601 33380 -603 33390
rect -2601 33378 -763 33380
rect 151963 33178 152123 33179
rect 151963 33019 151963 33178
rect 152122 33019 152123 33178
rect 151963 33019 152123 33019
rect -2987 32400 -1881 32560
rect -1003 32461 -902 32461
rect -1337 32361 -1003 32461
rect -903 32361 -902 32461
rect -1003 32360 -902 32361
rect -2601 32026 -603 32038
rect -2601 31890 -751 32026
rect -615 31890 -603 32026
rect -2601 31880 -603 31890
rect -2601 31878 -763 31880
rect 151963 31678 152123 31679
rect 151963 31519 151963 31678
rect 152122 31519 152123 31678
rect 151963 31519 152123 31519
rect -2987 30900 -1881 31060
rect -1003 30961 -902 30961
rect -1337 30861 -1003 30961
rect -903 30861 -902 30961
rect -1003 30860 -902 30861
rect -2601 30526 -603 30538
rect -2601 30390 -751 30526
rect -615 30390 -603 30526
rect -2601 30380 -603 30390
rect -2601 30378 -763 30380
rect 151963 30178 152123 30179
rect 151963 30019 151963 30178
rect 152122 30019 152123 30178
rect 151963 30019 152123 30019
rect -2987 29400 -1881 29560
rect -1003 29461 -902 29461
rect -1337 29361 -1003 29461
rect -903 29361 -902 29461
rect -1003 29360 -902 29361
rect -2601 29026 -603 29038
rect -2601 28890 -751 29026
rect -615 28890 -603 29026
rect -2601 28880 -603 28890
rect -2601 28878 -763 28880
rect 151963 28678 152123 28679
rect 151963 28519 151963 28678
rect 152122 28519 152123 28678
rect 151963 28519 152123 28519
rect -1003 27961 -902 27961
rect -1337 27861 -1003 27961
rect -903 27861 -902 27961
rect -1003 27860 -902 27861
rect -2601 27526 -603 27538
rect -2601 27390 -751 27526
rect -615 27390 -603 27526
rect -2601 27380 -603 27390
rect -2601 27378 -763 27380
rect 151963 27178 152123 27179
rect 151963 27019 151963 27178
rect 152122 27019 152123 27178
rect 151963 27019 152123 27019
rect -2987 26400 -1881 26560
rect -1003 26461 -902 26461
rect -1337 26361 -1003 26461
rect -903 26361 -902 26461
rect -1003 26360 -902 26361
rect -2601 26026 -603 26038
rect -2601 25890 -751 26026
rect -615 25890 -603 26026
rect -2601 25880 -603 25890
rect -2601 25878 -763 25880
rect 151963 25678 152123 25679
rect 151963 25519 151963 25678
rect 152122 25519 152123 25678
rect 151963 25519 152123 25519
rect -2987 24900 -1881 25060
rect -1003 24961 -902 24961
rect -1337 24861 -1003 24961
rect -903 24861 -902 24961
rect -1003 24860 -902 24861
rect -2601 24526 -603 24538
rect -2601 24390 -751 24526
rect -615 24390 -603 24526
rect -2601 24380 -603 24390
rect -2601 24378 -763 24380
rect 151963 24178 152123 24179
rect 151963 24019 151963 24178
rect 152122 24019 152123 24178
rect 151963 24019 152123 24019
rect -2987 23400 -1881 23560
rect -1003 23461 -902 23461
rect -1337 23361 -1003 23461
rect -903 23361 -902 23461
rect -1003 23360 -902 23361
rect -2601 23026 -603 23038
rect -2601 22890 -751 23026
rect -615 22890 -603 23026
rect -2601 22880 -603 22890
rect -2601 22878 -763 22880
rect 151963 22678 152123 22679
rect 151963 22519 151963 22678
rect 152122 22519 152123 22678
rect 151963 22519 152123 22519
rect -2987 21900 -1881 22060
rect -1003 21961 -902 21961
rect -1337 21861 -1003 21961
rect -903 21861 -902 21961
rect -1003 21860 -902 21861
rect -2601 21526 -603 21538
rect -2601 21390 -751 21526
rect -615 21390 -603 21526
rect -2601 21380 -603 21390
rect -2601 21378 -763 21380
rect 151963 21178 152123 21179
rect 151963 21019 151963 21178
rect 152122 21019 152123 21178
rect 151963 21019 152123 21019
rect -2987 20400 -1881 20560
rect -1003 20461 -902 20461
rect -1337 20361 -1003 20461
rect -903 20361 -902 20461
rect -1003 20360 -902 20361
rect -2601 20026 -603 20038
rect -2601 19890 -751 20026
rect -615 19890 -603 20026
rect -2601 19880 -603 19890
rect -2601 19878 -763 19880
rect 151963 19678 152123 19679
rect 151963 19519 151963 19678
rect 152122 19519 152123 19678
rect 151963 19519 152123 19519
rect -2987 18900 -1881 19060
rect -1003 18961 -902 18961
rect -1337 18861 -1003 18961
rect -903 18861 -902 18961
rect -1003 18860 -902 18861
rect -2601 18526 -603 18538
rect -2601 18390 -751 18526
rect -615 18390 -603 18526
rect -2601 18380 -603 18390
rect -2601 18378 -763 18380
rect 151963 18178 152123 18179
rect 151963 18019 151963 18178
rect 152122 18019 152123 18178
rect 151963 18019 152123 18019
rect -2987 17400 -1881 17560
rect -1003 17461 -902 17461
rect -1337 17361 -1003 17461
rect -903 17361 -902 17461
rect -1003 17360 -902 17361
rect -2601 17026 -603 17038
rect -2601 16890 -751 17026
rect -615 16890 -603 17026
rect -2601 16880 -603 16890
rect -2601 16878 -763 16880
rect 151963 16678 152123 16679
rect 151963 16519 151963 16678
rect 152122 16519 152123 16678
rect 151963 16519 152123 16519
rect -2987 15900 -1881 16060
rect -1003 15961 -902 15961
rect -1337 15861 -1003 15961
rect -903 15861 -902 15961
rect -1003 15860 -902 15861
rect -2601 15526 -603 15538
rect -2601 15390 -751 15526
rect -615 15390 -603 15526
rect -2601 15380 -603 15390
rect -2601 15378 -763 15380
rect 151963 15178 152123 15179
rect 151963 15019 151963 15178
rect 152122 15019 152123 15178
rect 151963 15019 152123 15019
rect -2987 14400 -1881 14560
rect -1003 14461 -902 14461
rect -1337 14361 -1003 14461
rect -903 14361 -902 14461
rect -1003 14360 -902 14361
rect -2601 14026 -603 14038
rect -2601 13890 -751 14026
rect -615 13890 -603 14026
rect -2601 13880 -603 13890
rect -2601 13878 -763 13880
rect 151963 13678 152123 13679
rect 151963 13519 151963 13678
rect 152122 13519 152123 13678
rect 151963 13519 152123 13519
rect -2987 12900 -1881 13060
rect -1003 12961 -902 12961
rect -1337 12861 -1003 12961
rect -903 12861 -902 12961
rect -1003 12860 -902 12861
rect -2601 12526 -603 12538
rect -2601 12390 -751 12526
rect -615 12390 -603 12526
rect -2601 12380 -603 12390
rect -2601 12378 -763 12380
rect 151963 12178 152123 12179
rect 151963 12019 151963 12178
rect 152122 12019 152123 12178
rect 151963 12019 152123 12019
rect -2987 11400 -1881 11560
rect -1003 11461 -902 11461
rect -1337 11361 -1003 11461
rect -903 11361 -902 11461
rect -1003 11360 -902 11361
rect -2601 11026 -603 11038
rect -2601 10890 -751 11026
rect -615 10890 -603 11026
rect -2601 10880 -603 10890
rect -2601 10878 -763 10880
rect 151963 10678 152123 10679
rect 151963 10519 151963 10678
rect 152122 10519 152123 10678
rect 151963 10519 152123 10519
rect -2987 9900 -1881 10060
rect -2601 9526 -603 9538
rect -2601 9390 -751 9526
rect -615 9390 -603 9526
rect -2601 9380 -603 9390
rect -390 9397 869 9452
rect -2601 9378 -763 9380
rect -3047 8971 -2996 8971
rect -2997 8871 -2996 8971
rect -3047 8870 -2996 8871
rect -390 8398 -335 9397
rect 1164 9233 1274 9749
rect 2664 9405 2774 9803
rect 3735 9446 3860 9455
rect 4164 9446 4274 9827
rect 3735 9445 4274 9446
rect 2658 9392 2783 9405
rect 1832 9379 1992 9380
rect 1158 9219 1283 9233
rect 1832 9220 1832 9379
rect 1991 9220 1992 9379
rect 2658 9283 2664 9392
rect 2773 9283 2783 9392
rect 3735 9336 3741 9445
rect 3850 9336 4274 9445
rect 3735 9336 4274 9336
rect 5346 9418 5471 9429
rect 5664 9418 5774 9839
rect 5346 9417 5774 9418
rect 3735 9326 3860 9336
rect 5346 9308 5356 9417
rect 5465 9308 5774 9417
rect 6895 9465 7020 9475
rect 7164 9465 7274 9839
rect 6895 9464 7274 9465
rect 6895 9355 6901 9464
rect 7010 9355 7274 9464
rect 6895 9355 7274 9355
rect 8450 9408 8575 9412
rect 8664 9408 8774 9836
rect 9925 9597 10050 9601
rect 10164 9597 10274 9839
rect 9925 9596 10274 9597
rect 9925 9487 9935 9596
rect 10044 9487 10274 9596
rect 9925 9487 10274 9487
rect 9925 9472 10050 9487
rect 8450 9408 8774 9408
rect 6895 9346 7020 9355
rect 5346 9308 5774 9308
rect 5346 9300 5471 9308
rect 8450 9299 8456 9408
rect 8565 9299 8774 9408
rect 8450 9298 8774 9299
rect 9044 9379 9204 9380
rect 8450 9283 8575 9298
rect 2658 9276 2783 9283
rect 1832 9220 1992 9220
rect 9044 9220 9044 9379
rect 9203 9220 9204 9379
rect 9044 9220 9204 9220
rect 11436 9329 11594 9336
rect 11664 9329 11774 9839
rect 12954 9506 13113 9514
rect 13164 9506 13274 9839
rect 14664 9531 14774 9839
rect 12954 9505 13274 9506
rect 12954 9396 12972 9505
rect 13081 9396 13274 9505
rect 14542 9530 14774 9531
rect 14542 9421 14542 9530
rect 14651 9421 14774 9530
rect 14542 9421 14774 9421
rect 16164 9493 16274 9839
rect 17664 9533 17774 9798
rect 19164 9613 19274 9817
rect 19156 9609 19281 9613
rect 12954 9396 13274 9396
rect 12954 9381 13113 9396
rect 16164 9384 16164 9493
rect 16273 9384 16274 9493
rect 17649 9527 17792 9533
rect 17649 9418 17664 9527
rect 17773 9418 17792 9527
rect 19156 9500 19164 9609
rect 19273 9500 19281 9609
rect 19156 9484 19281 9500
rect 20664 9446 20774 9839
rect 22164 9468 22274 9836
rect 23664 9572 23774 9839
rect 23659 9565 23784 9572
rect 22160 9461 22285 9468
rect 17649 9414 17792 9418
rect 20659 9436 20784 9446
rect 16164 9383 16274 9384
rect 11436 9329 11774 9329
rect 11436 9220 11449 9329
rect 11558 9220 11774 9329
rect 16457 9379 16617 9380
rect 17664 9379 17774 9414
rect 16457 9220 16457 9379
rect 16616 9220 16617 9379
rect 20659 9327 20664 9436
rect 20773 9327 20784 9436
rect 22160 9352 22164 9461
rect 22273 9352 22285 9461
rect 23659 9456 23664 9565
rect 23773 9456 23784 9565
rect 23659 9443 23784 9456
rect 25164 9511 25274 9827
rect 26664 9532 26774 9839
rect 28164 9581 28274 9833
rect 28164 9581 28417 9581
rect 26664 9521 26885 9532
rect 25164 9505 25375 9511
rect 25164 9396 25258 9505
rect 25367 9396 25375 9505
rect 26664 9412 26769 9521
rect 26878 9412 26885 9521
rect 28164 9472 28308 9581
rect 28417 9472 28417 9581
rect 28164 9471 28417 9472
rect 26664 9411 26885 9412
rect 26760 9403 26885 9411
rect 29664 9433 29774 9839
rect 29664 9433 29925 9433
rect 25164 9396 25375 9396
rect 25250 9382 25375 9396
rect 22160 9339 22285 9352
rect 20659 9317 20784 9327
rect 29664 9324 29815 9433
rect 29924 9324 29925 9433
rect 29664 9323 29925 9324
rect 31164 9395 31274 9839
rect 32664 9441 32774 9822
rect 34164 9476 34274 9819
rect 32664 9440 32981 9441
rect 31164 9395 31426 9395
rect 31164 9286 31316 9395
rect 31425 9286 31426 9395
rect 31164 9285 31426 9286
rect 32128 9379 32288 9380
rect 16457 9220 16617 9220
rect 32128 9220 32128 9379
rect 32287 9220 32288 9379
rect 32664 9331 32871 9440
rect 32980 9331 32981 9440
rect 34164 9367 34164 9476
rect 34273 9367 34274 9476
rect 35664 9530 35774 9815
rect 35664 9530 36074 9530
rect 35664 9421 35964 9530
rect 36073 9421 36074 9530
rect 35664 9420 36074 9421
rect 37164 9515 37274 9838
rect 37164 9515 37649 9515
rect 37164 9406 37539 9515
rect 37648 9406 37649 9515
rect 37164 9405 37649 9406
rect 34164 9366 34274 9367
rect 32664 9331 32981 9331
rect 32128 9220 32288 9220
rect 1158 9110 1164 9219
rect 1273 9110 1283 9219
rect 11436 9219 11774 9220
rect 11436 9203 11594 9219
rect 1158 9104 1283 9110
rect 38664 9153 38774 9839
rect 40164 9453 40274 9838
rect 40164 9452 40705 9453
rect 40164 9343 40595 9452
rect 40704 9343 40705 9452
rect 40164 9343 40705 9343
rect 41664 9202 41774 9831
rect 41664 9201 42247 9202
rect 38664 9153 39159 9153
rect 38664 9044 39049 9153
rect 39158 9044 39159 9153
rect 41664 9092 42137 9201
rect 42246 9092 42247 9201
rect 41664 9092 42247 9092
rect 43164 9157 43274 9839
rect 44664 9419 44774 9816
rect 44664 9418 45316 9419
rect 44664 9309 45206 9418
rect 45315 9309 45316 9418
rect 44664 9309 45316 9309
rect 46164 9397 46274 9812
rect 47664 9438 47774 9816
rect 47664 9437 48336 9438
rect 46164 9396 46888 9397
rect 46164 9287 46778 9396
rect 46887 9287 46888 9396
rect 47664 9328 48227 9437
rect 48336 9328 48336 9437
rect 47664 9328 48336 9328
rect 46164 9287 46888 9287
rect 49164 9251 49274 9819
rect 50664 9370 50774 9805
rect 52164 9378 52274 9816
rect 53664 9516 53774 9812
rect 53664 9516 54560 9516
rect 53664 9407 54451 9516
rect 54560 9407 54560 9516
rect 53664 9406 54560 9407
rect 55164 9468 55274 9823
rect 56664 9492 56774 9829
rect 56664 9492 57586 9492
rect 55164 9467 56084 9468
rect 52164 9377 52947 9378
rect 50664 9370 51465 9370
rect 50664 9261 51356 9370
rect 51465 9261 51465 9370
rect 52164 9268 52838 9377
rect 52947 9268 52947 9377
rect 55164 9358 55974 9467
rect 56083 9358 56084 9467
rect 56664 9383 57477 9492
rect 57586 9383 57586 9492
rect 56664 9382 57586 9383
rect 58164 9489 58274 9806
rect 58164 9488 59094 9489
rect 58164 9379 58984 9488
rect 59093 9379 59094 9488
rect 58164 9379 59094 9379
rect 59664 9432 59774 9839
rect 59664 9432 60685 9432
rect 55164 9358 56084 9358
rect 59664 9323 60575 9432
rect 60684 9323 60685 9432
rect 61164 9426 61274 9829
rect 62664 9471 62774 9839
rect 62664 9471 63730 9471
rect 61164 9425 62169 9426
rect 59664 9322 60685 9323
rect 60839 9379 60999 9380
rect 52164 9268 52947 9268
rect 50664 9260 51465 9261
rect 49164 9250 49908 9251
rect 43164 9157 43777 9157
rect 43164 9048 43668 9157
rect 43777 9048 43777 9157
rect 49164 9141 49799 9250
rect 49908 9141 49908 9250
rect 60839 9220 60839 9379
rect 60998 9220 60999 9379
rect 61164 9316 62059 9425
rect 62168 9316 62169 9425
rect 62664 9362 63621 9471
rect 63730 9362 63730 9471
rect 62664 9361 63730 9362
rect 64164 9407 64274 9822
rect 65664 9433 65774 9837
rect 65664 9433 66816 9433
rect 64164 9406 65235 9407
rect 61164 9316 62169 9316
rect 64164 9297 65125 9406
rect 65234 9297 65235 9406
rect 65664 9324 66706 9433
rect 66815 9324 66816 9433
rect 65664 9323 66816 9324
rect 64164 9297 65235 9297
rect 60839 9220 60999 9220
rect 49164 9141 49908 9141
rect 43164 9047 43777 9048
rect 67164 9121 67274 9829
rect 68664 9300 68774 9807
rect 70164 9334 70274 9839
rect 71664 9422 71774 9837
rect 73164 9422 73274 9833
rect 71664 9421 72899 9422
rect 70164 9334 71409 9334
rect 68664 9300 69886 9300
rect 68664 9191 69776 9300
rect 69885 9191 69886 9300
rect 70164 9225 71300 9334
rect 71409 9225 71409 9334
rect 71664 9312 72789 9421
rect 72898 9312 72899 9421
rect 71664 9312 72899 9312
rect 73164 9421 74487 9422
rect 73164 9312 74377 9421
rect 74486 9312 74487 9421
rect 73164 9312 74487 9312
rect 74664 9387 74774 9829
rect 76164 9429 76274 9829
rect 77664 9499 77774 9829
rect 77664 9498 79031 9499
rect 76164 9429 77506 9429
rect 74664 9387 75996 9387
rect 74664 9278 75886 9387
rect 75995 9278 75996 9387
rect 76164 9320 77396 9429
rect 77505 9320 77506 9429
rect 77664 9389 78922 9498
rect 79031 9389 79031 9498
rect 77664 9389 79031 9389
rect 76164 9319 77506 9320
rect 79164 9379 79274 9839
rect 80664 9445 80774 9833
rect 82164 9514 82274 9833
rect 83664 9568 83774 9829
rect 79164 9379 80576 9379
rect 74664 9277 75996 9278
rect 79164 9270 80443 9379
rect 80552 9270 80576 9379
rect 80664 9335 81778 9445
rect 82164 9404 83074 9514
rect 83664 9458 84541 9568
rect 79164 9269 80576 9270
rect 70164 9224 71409 9225
rect 81619 9229 81729 9335
rect 68664 9190 69886 9191
rect 67164 9120 68343 9121
rect 38664 9043 39159 9044
rect 67164 9011 68234 9120
rect 68343 9011 68343 9120
rect 81619 9120 81619 9229
rect 81728 9120 81729 9229
rect 81619 9120 81729 9120
rect 67164 9011 68343 9011
rect 82964 9087 83074 9404
rect 83774 9379 83934 9380
rect 83774 9220 83774 9379
rect 83933 9220 83934 9379
rect 83774 9220 83934 9220
rect 82964 8978 82964 9087
rect 83073 8978 83074 9087
rect 82964 8977 83074 8978
rect 84431 8710 84541 9458
rect 85164 9245 85274 9821
rect 86664 9568 86774 9839
rect 86664 9567 87293 9568
rect 86664 9458 87183 9567
rect 87292 9458 87293 9567
rect 86664 9458 87293 9458
rect 88164 9406 88274 9814
rect 88164 9297 88164 9406
rect 88273 9297 88274 9406
rect 88164 9296 88274 9297
rect 85164 9244 86651 9245
rect 85164 9135 86541 9244
rect 86650 9135 86651 9244
rect 85164 9135 86651 9135
rect 89664 8930 89774 9839
rect 91164 9391 91274 9829
rect 90274 9379 90434 9380
rect 90274 9220 90274 9379
rect 90433 9220 90434 9379
rect 91164 9281 92115 9391
rect 90274 9220 90434 9220
rect 89664 8929 91346 8930
rect 89664 8820 91237 8929
rect 91346 8820 91346 8929
rect 89664 8820 91346 8820
rect 84431 8601 84432 8710
rect 84541 8601 84541 8710
rect 84431 8601 84541 8601
rect 92005 8576 92115 9281
rect 92664 9018 92774 9839
rect 92664 8909 92664 9018
rect 92773 8909 92774 9018
rect 92664 8908 92774 8909
rect 94164 8829 94274 9829
rect 94774 9379 94934 9380
rect 94774 9220 94774 9379
rect 94933 9220 94934 9379
rect 94774 9220 94934 9220
rect 95664 9313 95774 9817
rect 95664 9203 96842 9313
rect 94164 8720 94164 8829
rect 94273 8720 94274 8829
rect 94164 8720 94274 8720
rect 92005 8467 92005 8576
rect 92114 8467 92115 8576
rect 92005 8466 92115 8467
rect 96732 8509 96842 9203
rect 97164 8965 97274 9812
rect 98664 8978 98774 9830
rect 100164 9402 100274 9812
rect 99274 9379 99434 9380
rect 99274 9220 99274 9379
rect 99433 9220 99434 9379
rect 100164 9292 101111 9402
rect 99274 9220 99434 9220
rect 98664 8978 100567 8978
rect 97164 8964 98506 8965
rect 97164 8855 98397 8964
rect 98506 8855 98506 8964
rect 98664 8869 100458 8978
rect 100567 8869 100567 8978
rect 98664 8868 100567 8869
rect 97164 8855 98506 8855
rect 96732 8400 96733 8509
rect 96842 8400 96842 8509
rect 96732 8400 96842 8400
rect 101001 8447 101111 9292
rect 101664 8876 101774 9835
rect 102274 9379 102434 9380
rect 102274 9220 102274 9379
rect 102433 9220 102434 9379
rect 102274 9220 102434 9220
rect 103164 9227 103274 9839
rect 103164 9118 103164 9227
rect 103273 9118 103274 9227
rect 103164 9118 103274 9118
rect 104664 9049 104774 9826
rect 106164 9442 106274 9817
rect 105774 9379 105934 9380
rect 105774 9220 105774 9379
rect 105933 9220 105934 9379
rect 106164 9332 107062 9442
rect 105774 9220 105934 9220
rect 104664 9049 106687 9049
rect 104664 8940 106578 9049
rect 106687 8940 106687 9049
rect 104664 8939 106687 8940
rect 101664 8875 103609 8876
rect 101664 8766 103500 8875
rect 103609 8766 103609 8875
rect 101664 8766 103609 8766
rect 106952 8634 107062 9332
rect 107664 9281 107774 9833
rect 109164 9447 109274 9839
rect 109164 9337 110454 9447
rect 107664 9172 107664 9281
rect 107773 9172 107774 9281
rect 107664 9172 107774 9172
rect 106952 8525 106952 8634
rect 107061 8525 107062 8634
rect 106952 8525 107062 8525
rect 110344 8614 110454 9337
rect 110664 8855 110774 9833
rect 111774 9379 111934 9380
rect 111774 9220 111774 9379
rect 111933 9220 111934 9379
rect 111774 9220 111934 9220
rect 112164 9214 112274 9828
rect 113664 9470 113774 9837
rect 113664 9469 114939 9470
rect 113664 9360 114829 9469
rect 114938 9360 114939 9469
rect 113664 9360 114939 9360
rect 112164 9214 113707 9214
rect 112164 9105 113597 9214
rect 113706 9105 113707 9214
rect 112164 9104 113707 9105
rect 115164 9152 115274 9824
rect 116274 9379 116434 9380
rect 116274 9220 116274 9379
rect 116433 9220 116434 9379
rect 116664 9344 116774 9839
rect 116664 9235 116664 9344
rect 116773 9235 116774 9344
rect 116664 9235 116774 9235
rect 116274 9220 116434 9220
rect 115164 9151 117435 9152
rect 115164 9042 117325 9151
rect 117434 9042 117435 9151
rect 115164 9042 117435 9042
rect 118164 9008 118274 9749
rect 119274 9379 119434 9380
rect 119274 9220 119274 9379
rect 119433 9220 119434 9379
rect 119274 9220 119434 9220
rect 119664 9267 119774 9805
rect 121164 9285 121274 9839
rect 119664 9267 120946 9267
rect 119664 9158 120836 9267
rect 120945 9158 120946 9267
rect 121164 9176 121164 9285
rect 121273 9176 121274 9285
rect 122664 9299 122774 9839
rect 124164 9545 124274 9827
rect 124164 9435 124943 9545
rect 122664 9189 124465 9299
rect 121164 9175 121274 9176
rect 119664 9157 120946 9158
rect 118164 9007 120568 9008
rect 118164 8898 120458 9007
rect 120567 8898 120568 9007
rect 118164 8898 120568 8898
rect 110664 8746 110664 8855
rect 110773 8746 110774 8855
rect 110664 8746 110774 8746
rect 110344 8505 110344 8614
rect 110453 8505 110454 8614
rect 110344 8504 110454 8505
rect 124355 8538 124465 9189
rect 124833 8930 124943 9435
rect 125274 9379 125434 9380
rect 125274 9220 125274 9379
rect 125433 9220 125434 9379
rect 125274 9220 125434 9220
rect 125664 9255 125774 9839
rect 127164 9350 127274 9839
rect 125664 9254 127072 9255
rect 125664 9145 126963 9254
rect 127072 9145 127072 9254
rect 127164 9241 127164 9350
rect 127273 9241 127274 9350
rect 127164 9240 127274 9241
rect 128664 9288 128774 9835
rect 130164 9558 130274 9839
rect 130164 9448 130632 9558
rect 128664 9178 130136 9288
rect 125664 9145 127072 9145
rect 124833 8821 124834 8930
rect 124943 8821 124943 8930
rect 124833 8820 124943 8821
rect -2167 8343 -335 8398
rect -2167 6988 -2112 8343
rect 101001 8338 101002 8447
rect 101111 8338 101111 8447
rect 124355 8429 124356 8538
rect 124465 8429 124465 8538
rect 130026 8623 130136 9178
rect 130522 9062 130632 9448
rect 130522 8953 130522 9062
rect 130631 8953 130632 9062
rect 130522 8953 130632 8953
rect 131664 8982 131774 9839
rect 131974 9379 132134 9380
rect 131974 9220 131974 9379
rect 132133 9220 132134 9379
rect 131974 9220 132134 9220
rect 133164 9280 133274 9810
rect 133164 9280 134626 9280
rect 133164 9171 134516 9280
rect 134625 9171 134626 9280
rect 133164 9170 134626 9171
rect 134664 9134 134774 9797
rect 134974 9379 135134 9380
rect 134974 9220 134974 9379
rect 135133 9220 135134 9379
rect 134974 9220 135134 9220
rect 134664 9025 134664 9134
rect 134773 9025 134774 9134
rect 134664 9024 134774 9025
rect 131664 8981 133073 8982
rect 131664 8872 132935 8981
rect 133044 8872 133073 8981
rect 131664 8872 133073 8872
rect 136164 8791 136274 9824
rect 136474 9379 136634 9380
rect 136474 9220 136474 9379
rect 136633 9220 136634 9379
rect 136474 9220 136634 9220
rect 137664 9103 137774 9824
rect 137974 9379 138134 9380
rect 137974 9220 137974 9379
rect 138133 9220 138134 9379
rect 139164 9349 139274 9835
rect 139164 9349 139948 9349
rect 139164 9240 139838 9349
rect 139947 9240 139948 9349
rect 139164 9239 139948 9240
rect 137974 9220 138134 9220
rect 137664 9103 139549 9103
rect 137664 8994 139439 9103
rect 139548 8994 139549 9103
rect 137664 8993 139549 8994
rect 136164 8791 138956 8791
rect 136164 8682 138847 8791
rect 138956 8682 138956 8791
rect 136164 8681 138956 8682
rect 140664 8756 140774 9839
rect 140974 9379 141134 9380
rect 140974 9220 140974 9379
rect 141133 9220 141134 9379
rect 140974 9220 141134 9220
rect 142164 9068 142274 9839
rect 142974 9379 143134 9380
rect 142974 9220 142974 9379
rect 143133 9220 143134 9379
rect 142974 9220 143134 9220
rect 142164 8959 142164 9068
rect 142273 8959 142274 9068
rect 143664 9114 143774 9835
rect 145164 9477 145274 9839
rect 145164 9368 145164 9477
rect 145273 9368 145274 9477
rect 145164 9368 145274 9368
rect 143664 9113 146313 9114
rect 143664 9004 146204 9113
rect 146313 9004 146313 9113
rect 143664 9004 146313 9004
rect 142164 8959 142274 8959
rect 146664 8862 146774 9821
rect 146974 9379 147134 9380
rect 146974 9220 146974 9379
rect 147133 9220 147134 9379
rect 146974 9220 147134 9220
rect 148164 9164 148274 9827
rect 149664 9550 149774 9839
rect 149664 9549 152802 9550
rect 149664 9440 152693 9549
rect 152802 9440 152802 9549
rect 149664 9440 152802 9440
rect 148474 9379 148634 9380
rect 148474 9220 148474 9379
rect 148633 9220 148634 9379
rect 148474 9220 148634 9220
rect 149974 9379 150134 9380
rect 149974 9220 149974 9379
rect 150133 9220 150134 9379
rect 149974 9220 150134 9220
rect 151474 9379 151634 9380
rect 151474 9220 151474 9379
rect 151633 9220 151634 9379
rect 151474 9220 151634 9220
rect 148164 9054 150235 9164
rect 146664 8861 149739 8862
rect 140664 8756 143574 8756
rect 140664 8647 143465 8756
rect 143574 8647 143574 8756
rect 146664 8752 149629 8861
rect 149738 8752 149739 8861
rect 146664 8752 149739 8752
rect 140664 8646 143574 8647
rect 130026 8514 130027 8623
rect 130136 8514 130136 8623
rect 130026 8513 130136 8514
rect 150125 8552 150235 9054
rect 150125 8443 150126 8552
rect 150235 8443 150235 8552
rect 150125 8443 150235 8443
rect 151933 8632 152093 8644
rect 151933 8496 151945 8632
rect 152081 8496 152093 8632
rect 124355 8429 124465 8429
rect 101001 8337 101111 8338
rect 151470 8205 151637 8206
rect 151470 8205 151471 8205
rect 151637 8205 151637 8205
rect 9041 7853 9207 7854
rect 9041 7853 9041 7853
rect 9206 7853 9207 7853
rect 83771 7853 83937 7854
rect 83771 7853 83771 7853
rect 83936 7853 83937 7853
rect 1829 7844 1995 7845
rect 1829 7844 1829 7844
rect 1994 7844 1995 7844
rect 60836 7852 61002 7853
rect 60836 7852 60836 7852
rect 61001 7852 61002 7852
rect 32125 7845 32291 7846
rect 32125 7845 32125 7845
rect 32290 7845 32291 7845
rect 16454 7841 16620 7842
rect 16454 7841 16454 7841
rect 16619 7841 16620 7841
rect 90271 7853 90437 7854
rect 90271 7853 90271 7853
rect 90436 7853 90437 7853
rect 94771 7853 94937 7854
rect 94771 7853 94771 7853
rect 94936 7853 94937 7853
rect 99271 7853 99437 7854
rect 99271 7853 99271 7853
rect 99436 7853 99437 7853
rect 102271 7853 102437 7854
rect 102271 7853 102271 7853
rect 102436 7853 102437 7853
rect 105771 7853 105937 7854
rect 105771 7853 105771 7853
rect 105936 7853 105937 7853
rect 111771 7853 111937 7854
rect 111771 7853 111771 7853
rect 111936 7853 111937 7853
rect 116271 7853 116437 7854
rect 116271 7853 116271 7853
rect 116436 7853 116437 7853
rect 119271 7853 119437 7854
rect 119271 7853 119271 7853
rect 119436 7853 119437 7853
rect 125271 7853 125437 7854
rect 125271 7853 125271 7853
rect 125436 7853 125437 7853
rect 131971 7853 132137 7854
rect 131971 7853 131971 7853
rect 132136 7853 132137 7853
rect 134971 7853 135137 7854
rect 134971 7853 134971 7853
rect 135136 7853 135137 7853
rect 136471 7853 136637 7854
rect 136471 7853 136471 7853
rect 136636 7853 136637 7853
rect 137971 7853 138137 7854
rect 137971 7853 137971 7853
rect 138136 7853 138137 7853
rect 140971 7853 141137 7854
rect 140971 7853 140971 7853
rect 141136 7853 141137 7853
rect 142971 7853 143137 7854
rect 142971 7853 142971 7853
rect 143136 7853 143137 7853
rect 146971 7853 147137 7854
rect 146971 7853 146971 7853
rect 147136 7853 147137 7853
rect 148471 7853 148637 7854
rect 148471 7853 148471 7853
rect 148636 7853 148637 7853
rect 149971 7853 150137 7854
rect 149971 7853 149971 7853
rect 150136 7853 150137 7853
rect 151471 7853 151637 7854
rect 151471 7853 151471 7853
rect 151636 7853 151637 7853
rect 151933 7846 152093 8496
rect 151841 7698 151933 7834
<< via4 >>
rect -2761 160878 -2601 161038
rect -751 160890 -615 161026
rect 151224 162269 151384 162299
rect 151224 162169 151251 162269
rect 151251 162169 151356 162269
rect 151356 162169 151384 162269
rect 151224 162139 151384 162169
rect 151975 160531 152111 160667
rect -3147 159900 -2987 160060
rect -1881 159900 -1721 160060
rect -1497 159831 -1337 159991
rect -2761 159378 -2601 159538
rect -751 159390 -615 159526
rect 151975 159031 152111 159167
rect -3147 158400 -2987 158560
rect -1881 158400 -1721 158560
rect -1497 158331 -1337 158491
rect -2761 157878 -2601 158038
rect -751 157890 -615 158026
rect 151975 157531 152111 157667
rect -3147 156900 -2987 157060
rect -1881 156900 -1721 157060
rect -1497 156831 -1337 156991
rect -2761 156378 -2601 156538
rect -751 156390 -615 156526
rect 151975 156031 152111 156167
rect -3147 155400 -2987 155560
rect -1881 155400 -1721 155560
rect -1497 155331 -1337 155491
rect -2761 154878 -2601 155038
rect -751 154890 -615 155026
rect 151975 154531 152111 154667
rect -3147 153900 -2987 154060
rect -1881 153900 -1721 154060
rect -1497 153831 -1337 153991
rect -2761 153378 -2601 153538
rect -751 153390 -615 153526
rect 151975 153031 152111 153167
rect -3147 152400 -2987 152560
rect -1881 152400 -1721 152560
rect -1497 152331 -1337 152491
rect -2761 151878 -2601 152038
rect -751 151890 -615 152026
rect 151975 151531 152111 151667
rect -3147 150900 -2987 151060
rect -1881 150900 -1721 151060
rect -1497 150831 -1337 150991
rect -2761 150378 -2601 150538
rect -751 150390 -615 150526
rect 151975 150031 152111 150167
rect -3147 149400 -2987 149560
rect -1881 149400 -1721 149560
rect -1497 149331 -1337 149491
rect -2761 148878 -2601 149038
rect -751 148890 -615 149026
rect 151975 148531 152111 148667
rect -3147 147900 -2987 148060
rect -1881 147900 -1721 148060
rect -1497 147831 -1337 147991
rect -2761 147378 -2601 147538
rect -751 147390 -615 147526
rect 151975 147031 152111 147167
rect -3147 146400 -2987 146560
rect -1881 146400 -1721 146560
rect -1497 146331 -1337 146491
rect -2761 145878 -2601 146038
rect -751 145890 -615 146026
rect 151975 145531 152111 145667
rect -3147 144900 -2987 145060
rect -1881 144900 -1721 145060
rect -1497 144831 -1337 144991
rect -2761 144378 -2601 144538
rect -751 144390 -615 144526
rect 151975 144031 152111 144167
rect -3147 143400 -2987 143560
rect -1881 143400 -1721 143560
rect -1497 143331 -1337 143491
rect -2761 142878 -2601 143038
rect -751 142890 -615 143026
rect 151975 142531 152111 142667
rect -3147 141900 -2987 142060
rect -1881 141900 -1721 142060
rect -1497 141831 -1337 141991
rect -2761 141378 -2601 141538
rect -751 141390 -615 141526
rect 151975 141031 152111 141167
rect -3147 140400 -2987 140560
rect -1881 140400 -1721 140560
rect -1497 140331 -1337 140491
rect -2761 139878 -2601 140038
rect -751 139890 -615 140026
rect 151975 139531 152111 139667
rect -3147 138900 -2987 139060
rect -1881 138900 -1721 139060
rect -1497 138831 -1337 138991
rect -2761 138378 -2601 138538
rect -751 138390 -615 138526
rect 151975 138031 152111 138167
rect -3147 137400 -2987 137560
rect -1881 137400 -1721 137560
rect -1497 137331 -1337 137491
rect -2761 136878 -2601 137038
rect -751 136890 -615 137026
rect 151975 136531 152111 136667
rect -3147 135900 -2987 136060
rect -1881 135900 -1721 136060
rect -1497 135831 -1337 135991
rect -2761 135378 -2601 135538
rect -751 135390 -615 135526
rect 151975 135031 152111 135167
rect -3147 134400 -2987 134560
rect -1881 134400 -1721 134560
rect -1497 134331 -1337 134491
rect -2761 133878 -2601 134038
rect -751 133890 -615 134026
rect 151975 133531 152111 133667
rect -3147 132900 -2987 133060
rect -1881 132900 -1721 133060
rect -1497 132831 -1337 132991
rect -2761 132378 -2601 132538
rect -751 132390 -615 132526
rect 151975 132031 152111 132167
rect -3147 131400 -2987 131560
rect -1881 131400 -1721 131560
rect -1497 131331 -1337 131491
rect -2761 130878 -2601 131038
rect -751 130890 -615 131026
rect 151975 130531 152111 130667
rect -3147 129900 -2987 130060
rect -1881 129900 -1721 130060
rect -1497 129831 -1337 129991
rect -2761 129378 -2601 129538
rect -751 129390 -615 129526
rect 151975 129031 152111 129167
rect -3147 128400 -2987 128560
rect -1881 128400 -1721 128560
rect -1497 128331 -1337 128491
rect -2761 127878 -2601 128038
rect -751 127890 -615 128026
rect 151975 127531 152111 127667
rect -3147 126900 -2987 127060
rect -1881 126900 -1721 127060
rect -1497 126831 -1337 126991
rect -2761 126378 -2601 126538
rect -751 126390 -615 126526
rect 151975 126031 152111 126167
rect -3147 125400 -2987 125560
rect -1881 125400 -1721 125560
rect -1497 125331 -1337 125491
rect -2761 124878 -2601 125038
rect -751 124890 -615 125026
rect 151975 124531 152111 124667
rect -3147 123900 -2987 124060
rect -1881 123900 -1721 124060
rect -1497 123831 -1337 123991
rect 151975 123031 152111 123167
rect -3147 122400 -2987 122560
rect -1881 122400 -1721 122560
rect -1497 122331 -1337 122491
rect -2761 121878 -2601 122038
rect -751 121890 -615 122026
rect 151975 121531 152111 121667
rect -3147 120900 -2987 121060
rect -1881 120900 -1721 121060
rect -1497 120831 -1337 120991
rect -2761 120378 -2601 120538
rect -751 120390 -615 120526
rect 151975 120031 152111 120167
rect -3147 119400 -2987 119560
rect -1881 119400 -1721 119560
rect -1497 119331 -1337 119491
rect -2761 118878 -2601 119038
rect -751 118890 -615 119026
rect 151975 118531 152111 118667
rect -3147 117900 -2987 118060
rect -1881 117900 -1721 118060
rect -1497 117831 -1337 117991
rect -2761 117378 -2601 117538
rect -751 117390 -615 117526
rect 151975 117031 152111 117167
rect -3147 116400 -2987 116560
rect -1881 116400 -1721 116560
rect -1497 116331 -1337 116491
rect -2761 115878 -2601 116038
rect -751 115890 -615 116026
rect 151975 115531 152111 115667
rect -3147 114900 -2987 115060
rect -1881 114900 -1721 115060
rect -1497 114831 -1337 114991
rect -2761 114378 -2601 114538
rect -751 114390 -615 114526
rect 151975 114031 152111 114167
rect -3147 113400 -2987 113560
rect -1881 113400 -1721 113560
rect -1497 113331 -1337 113491
rect -2761 112878 -2601 113038
rect -751 112890 -615 113026
rect 151975 112531 152111 112667
rect -3147 111900 -2987 112060
rect -1881 111900 -1721 112060
rect -1497 111831 -1337 111991
rect -2761 111378 -2601 111538
rect -751 111390 -615 111526
rect 151975 111031 152111 111167
rect -3147 110400 -2987 110560
rect -1881 110400 -1721 110560
rect -1497 110331 -1337 110491
rect -2761 109878 -2601 110038
rect -751 109890 -615 110026
rect 151975 109531 152111 109667
rect -3147 108900 -2987 109060
rect -1881 108900 -1721 109060
rect -1497 108831 -1337 108991
rect -2761 108378 -2601 108538
rect -751 108390 -615 108526
rect 151975 108031 152111 108167
rect -3147 107400 -2987 107560
rect -1881 107400 -1721 107560
rect -1497 107331 -1337 107491
rect -2761 106878 -2601 107038
rect -751 106890 -615 107026
rect 151975 106531 152111 106667
rect -3147 105900 -2987 106060
rect -1881 105900 -1721 106060
rect -1497 105831 -1337 105991
rect -2761 105378 -2601 105538
rect -751 105390 -615 105526
rect 151975 105031 152111 105167
rect -1497 104331 -1337 104491
rect -2761 103878 -2601 104038
rect -751 103890 -615 104026
rect 151975 103531 152111 103667
rect -3147 102900 -2987 103060
rect -1881 102900 -1721 103060
rect -1497 102831 -1337 102991
rect -2761 102378 -2601 102538
rect -751 102390 -615 102526
rect 151975 102031 152111 102167
rect -3147 101400 -2987 101560
rect -1881 101400 -1721 101560
rect -1497 101331 -1337 101491
rect -2761 100878 -2601 101038
rect -751 100890 -615 101026
rect 151975 100531 152111 100667
rect -3147 99900 -2987 100060
rect -1881 99900 -1721 100060
rect -1497 99831 -1337 99991
rect -2761 99378 -2601 99538
rect -751 99390 -615 99526
rect 151975 99031 152111 99167
rect -3147 98400 -2987 98560
rect -1881 98400 -1721 98560
rect -1497 98331 -1337 98491
rect -2761 97878 -2601 98038
rect -751 97890 -615 98026
rect 151975 97531 152111 97667
rect -3147 96900 -2987 97060
rect -1881 96900 -1721 97060
rect -1497 96831 -1337 96991
rect -2761 96378 -2601 96538
rect -751 96390 -615 96526
rect 151975 96031 152111 96167
rect -3147 95400 -2987 95560
rect -1881 95400 -1721 95560
rect -1497 95331 -1337 95491
rect -2761 94878 -2601 95038
rect -751 94890 -615 95026
rect 151975 94531 152111 94667
rect -3147 93900 -2987 94060
rect -1881 93900 -1721 94060
rect -1497 93831 -1337 93991
rect -2761 93378 -2601 93538
rect -751 93390 -615 93526
rect 151975 93031 152111 93167
rect -3147 92400 -2987 92560
rect -1881 92400 -1721 92560
rect -1497 92331 -1337 92491
rect -2761 91878 -2601 92038
rect -751 91890 -615 92026
rect 151975 91531 152111 91667
rect -3147 90900 -2987 91060
rect -1881 90900 -1721 91060
rect -1497 90831 -1337 90991
rect -2761 90378 -2601 90538
rect -751 90390 -615 90526
rect 151975 90031 152111 90167
rect -3147 89400 -2987 89560
rect -1881 89400 -1721 89560
rect -1497 89331 -1337 89491
rect -2761 88878 -2601 89038
rect -751 88890 -615 89026
rect 151975 88531 152111 88667
rect -3147 87900 -2987 88060
rect -1881 87900 -1721 88060
rect -1497 87831 -1337 87991
rect -2761 87378 -2601 87538
rect -751 87390 -615 87526
rect 151975 87031 152111 87167
rect -3147 86400 -2987 86560
rect -1881 86400 -1721 86560
rect -1497 86331 -1337 86491
rect -2761 85878 -2601 86038
rect -751 85890 -615 86026
rect 151975 85531 152111 85667
rect -3147 84900 -2987 85060
rect -1881 84900 -1721 85060
rect -1497 84831 -1337 84991
rect -2761 84378 -2601 84538
rect -751 84390 -615 84526
rect 151975 84031 152111 84167
rect -3147 83400 -2987 83560
rect -1881 83400 -1721 83560
rect -1497 83331 -1337 83491
rect -2761 82878 -2601 83038
rect -751 82890 -615 83026
rect 151975 82531 152111 82667
rect -3147 81900 -2987 82060
rect -1881 81900 -1721 82060
rect -1497 81831 -1337 81991
rect -2761 81378 -2601 81538
rect -751 81390 -615 81526
rect 151975 81031 152111 81167
rect -3147 80400 -2987 80560
rect -1881 80400 -1721 80560
rect -1497 80331 -1337 80491
rect -2761 79878 -2601 80038
rect -751 79890 -615 80026
rect 151975 79531 152111 79667
rect -3147 78900 -2987 79060
rect -1881 78900 -1721 79060
rect -1497 78831 -1337 78991
rect -2761 78378 -2601 78538
rect -751 78390 -615 78526
rect 151975 78031 152111 78167
rect -3147 77400 -2987 77560
rect -1881 77400 -1721 77560
rect -1497 77331 -1337 77491
rect -2761 76878 -2601 77038
rect -751 76890 -615 77026
rect 151975 76531 152111 76667
rect -3147 75900 -2987 76060
rect -1881 75900 -1721 76060
rect -1497 75831 -1337 75991
rect -2761 75378 -2601 75538
rect -751 75390 -615 75526
rect 151975 75031 152111 75167
rect -3147 74400 -2987 74560
rect -1881 74400 -1721 74560
rect -1497 74331 -1337 74491
rect -2761 73878 -2601 74038
rect -751 73890 -615 74026
rect 151975 73531 152111 73667
rect -3147 72900 -2987 73060
rect -1881 72900 -1721 73060
rect -1497 72831 -1337 72991
rect -2761 72378 -2601 72538
rect -751 72390 -615 72526
rect 151975 72031 152111 72167
rect -3147 71400 -2987 71560
rect -1881 71400 -1721 71560
rect -1497 71331 -1337 71491
rect -2761 70878 -2601 71038
rect -751 70890 -615 71026
rect 151975 70531 152111 70667
rect -3147 69900 -2987 70060
rect -1881 69900 -1721 70060
rect -1497 69831 -1337 69991
rect -2761 69378 -2601 69538
rect -751 69390 -615 69526
rect 151975 69031 152111 69167
rect -3147 68400 -2987 68560
rect -1881 68400 -1721 68560
rect -1497 68331 -1337 68491
rect -2761 67878 -2601 68038
rect -751 67890 -615 68026
rect 151975 67531 152111 67667
rect -3147 66900 -2987 67060
rect -1881 66900 -1721 67060
rect -1497 66831 -1337 66991
rect -2761 66378 -2601 66538
rect -751 66390 -615 66526
rect 151975 66031 152111 66167
rect -3147 65400 -2987 65560
rect -1881 65400 -1721 65560
rect -1497 65331 -1337 65491
rect -2761 64878 -2601 65038
rect -751 64890 -615 65026
rect 151975 64531 152111 64667
rect -3147 63900 -2987 64060
rect -1881 63900 -1721 64060
rect -1497 63831 -1337 63991
rect -2761 63378 -2601 63538
rect -751 63390 -615 63526
rect 151975 63031 152111 63167
rect -3147 62400 -2987 62560
rect -1881 62400 -1721 62560
rect -1497 62331 -1337 62491
rect -2761 61878 -2601 62038
rect -751 61890 -615 62026
rect 151975 61531 152111 61667
rect -3147 60900 -2987 61060
rect -1881 60900 -1721 61060
rect -1497 60831 -1337 60991
rect -2761 60378 -2601 60538
rect -751 60390 -615 60526
rect 151975 60031 152111 60167
rect -3147 59400 -2987 59560
rect -1881 59400 -1721 59560
rect -1497 59331 -1337 59491
rect -2761 58878 -2601 59038
rect -751 58890 -615 59026
rect 151975 58531 152111 58667
rect -3147 57900 -2987 58060
rect -1881 57900 -1721 58060
rect -1497 57831 -1337 57991
rect -2761 57378 -2601 57538
rect -751 57390 -615 57526
rect 151975 57031 152111 57167
rect -3147 56400 -2987 56560
rect -1881 56400 -1721 56560
rect -1497 56331 -1337 56491
rect -2761 55878 -2601 56038
rect -751 55890 -615 56026
rect 151975 55531 152111 55667
rect -3147 54900 -2987 55060
rect -1881 54900 -1721 55060
rect -1497 54831 -1337 54991
rect -2761 54378 -2601 54538
rect -751 54390 -615 54526
rect 151975 54031 152111 54167
rect -3147 53400 -2987 53560
rect -1881 53400 -1721 53560
rect -1497 53331 -1337 53491
rect -2761 52878 -2601 53038
rect -751 52890 -615 53026
rect 151975 52531 152111 52667
rect -3147 51900 -2987 52060
rect -1881 51900 -1721 52060
rect -1497 51831 -1337 51991
rect -2761 51378 -2601 51538
rect -751 51390 -615 51526
rect 151975 51031 152111 51167
rect -3147 50400 -2987 50560
rect -1881 50400 -1721 50560
rect -1497 50331 -1337 50491
rect -2761 49878 -2601 50038
rect -751 49890 -615 50026
rect 151975 49531 152111 49667
rect -3147 48900 -2987 49060
rect -1881 48900 -1721 49060
rect -1497 48831 -1337 48991
rect -2761 48378 -2601 48538
rect -751 48390 -615 48526
rect 151975 48031 152111 48167
rect -3147 47400 -2987 47560
rect -1881 47400 -1721 47560
rect -1497 47331 -1337 47491
rect 151975 46531 152111 46667
rect -3147 45900 -2987 46060
rect -1881 45900 -1721 46060
rect -1497 45831 -1337 45991
rect -2761 45378 -2601 45538
rect -751 45390 -615 45526
rect 151975 45031 152111 45167
rect -3147 44400 -2987 44560
rect -1881 44400 -1721 44560
rect -1497 44331 -1337 44491
rect -2761 43878 -2601 44038
rect -751 43890 -615 44026
rect 151975 43531 152111 43667
rect -3147 42900 -2987 43060
rect -1881 42900 -1721 43060
rect -1497 42831 -1337 42991
rect -2761 42378 -2601 42538
rect -751 42390 -615 42526
rect 151975 42031 152111 42167
rect -3147 41400 -2987 41560
rect -1881 41400 -1721 41560
rect -1497 41331 -1337 41491
rect -2761 40878 -2601 41038
rect -751 40890 -615 41026
rect 151975 40531 152111 40667
rect -3147 39900 -2987 40060
rect -1881 39900 -1721 40060
rect -1497 39831 -1337 39991
rect -2761 39378 -2601 39538
rect -751 39390 -615 39526
rect 151975 39031 152111 39167
rect -3147 38400 -2987 38560
rect -1881 38400 -1721 38560
rect -1497 38331 -1337 38491
rect -2761 37878 -2601 38038
rect -751 37890 -615 38026
rect 151975 37531 152111 37667
rect -3147 36900 -2987 37060
rect -1881 36900 -1721 37060
rect -1497 36831 -1337 36991
rect -2761 36378 -2601 36538
rect -751 36390 -615 36526
rect 151975 36031 152111 36167
rect -3147 35400 -2987 35560
rect -1881 35400 -1721 35560
rect -1497 35331 -1337 35491
rect -2761 34878 -2601 35038
rect -751 34890 -615 35026
rect 151975 34531 152111 34667
rect -3147 33900 -2987 34060
rect -1881 33900 -1721 34060
rect -1497 33831 -1337 33991
rect -2761 33378 -2601 33538
rect -751 33390 -615 33526
rect 151975 33031 152111 33167
rect -3147 32400 -2987 32560
rect -1881 32400 -1721 32560
rect -1497 32331 -1337 32491
rect -2761 31878 -2601 32038
rect -751 31890 -615 32026
rect 151975 31531 152111 31667
rect -3147 30900 -2987 31060
rect -1881 30900 -1721 31060
rect -1497 30831 -1337 30991
rect -2761 30378 -2601 30538
rect -751 30390 -615 30526
rect 151975 30031 152111 30167
rect -3147 29400 -2987 29560
rect -1881 29400 -1721 29560
rect -1497 29331 -1337 29491
rect -2761 28878 -2601 29038
rect -751 28890 -615 29026
rect 151975 28531 152111 28667
rect -1497 27831 -1337 27991
rect -2761 27378 -2601 27538
rect -751 27390 -615 27526
rect 151975 27031 152111 27167
rect -3147 26400 -2987 26560
rect -1881 26400 -1721 26560
rect -1497 26331 -1337 26491
rect -2761 25878 -2601 26038
rect -751 25890 -615 26026
rect 151975 25531 152111 25667
rect -3147 24900 -2987 25060
rect -1881 24900 -1721 25060
rect -1497 24831 -1337 24991
rect -2761 24378 -2601 24538
rect -751 24390 -615 24526
rect 151975 24031 152111 24167
rect -3147 23400 -2987 23560
rect -1881 23400 -1721 23560
rect -1497 23331 -1337 23491
rect -2761 22878 -2601 23038
rect -751 22890 -615 23026
rect 151975 22531 152111 22667
rect -3147 21900 -2987 22060
rect -1881 21900 -1721 22060
rect -1497 21831 -1337 21991
rect -2761 21378 -2601 21538
rect -751 21390 -615 21526
rect 151975 21031 152111 21167
rect -3147 20400 -2987 20560
rect -1881 20400 -1721 20560
rect -1497 20331 -1337 20491
rect -2761 19878 -2601 20038
rect -751 19890 -615 20026
rect 151975 19531 152111 19667
rect -3147 18900 -2987 19060
rect -1881 18900 -1721 19060
rect -1497 18831 -1337 18991
rect -2761 18378 -2601 18538
rect -751 18390 -615 18526
rect 151975 18031 152111 18167
rect -3147 17400 -2987 17560
rect -1881 17400 -1721 17560
rect -1497 17331 -1337 17491
rect -2761 16878 -2601 17038
rect -751 16890 -615 17026
rect 151975 16531 152111 16667
rect -3147 15900 -2987 16060
rect -1881 15900 -1721 16060
rect -1497 15831 -1337 15991
rect -2761 15378 -2601 15538
rect -751 15390 -615 15526
rect 151975 15031 152111 15167
rect -3147 14400 -2987 14560
rect -1881 14400 -1721 14560
rect -1497 14331 -1337 14491
rect -2761 13878 -2601 14038
rect -751 13890 -615 14026
rect 151975 13531 152111 13667
rect -3147 12900 -2987 13060
rect -1881 12900 -1721 13060
rect -1497 12831 -1337 12991
rect -2761 12378 -2601 12538
rect -751 12390 -615 12526
rect 151975 12031 152111 12167
rect -3147 11400 -2987 11560
rect -1881 11400 -1721 11560
rect -1497 11331 -1337 11491
rect -2761 10878 -2601 11038
rect -751 10890 -615 11026
rect 151975 10531 152111 10667
rect -3147 9900 -2987 10060
rect -1881 9900 -1721 10060
rect -2761 9378 -2601 9538
rect -751 9390 -615 9526
rect -3207 8971 -3047 9001
rect -3207 8871 -3102 8971
rect -3102 8871 -3047 8971
rect -3207 8841 -3047 8871
rect 1844 9232 1980 9368
rect 9056 9232 9192 9368
rect 16469 9232 16605 9368
rect 32140 9232 32276 9368
rect 60851 9232 60987 9368
rect 83786 9232 83922 9368
rect 90286 9232 90422 9368
rect 94786 9232 94922 9368
rect 99286 9232 99422 9368
rect 102286 9232 102422 9368
rect 105786 9232 105922 9368
rect 111786 9232 111922 9368
rect 116286 9232 116422 9368
rect 119286 9232 119422 9368
rect 125286 9232 125422 9368
rect 131986 9232 132122 9368
rect 134986 9232 135122 9368
rect 136486 9232 136622 9368
rect 137986 9232 138122 9368
rect 140986 9232 141122 9368
rect 142986 9232 143122 9368
rect 146986 9232 147122 9368
rect 148486 9232 148622 9368
rect 149986 9232 150122 9368
rect 151486 9232 151622 9368
rect 151945 8496 152081 8632
rect 151470 8044 151471 8205
rect 151471 8044 151637 8205
rect 151637 8044 151637 8205
rect 151470 8044 151637 8044
rect 24 7791 184 7821
rect 24 7691 51 7791
rect 51 7691 156 7791
rect 156 7691 184 7791
rect 24 7661 184 7691
rect 1829 7684 1829 7844
rect 1829 7684 1994 7844
rect 1994 7684 1995 7844
rect 9041 7693 9041 7853
rect 9041 7693 9206 7853
rect 9206 7693 9207 7853
rect 9041 7693 9207 7693
rect 1829 7684 1995 7684
rect 16454 7681 16454 7841
rect 16454 7681 16619 7841
rect 16619 7681 16620 7841
rect 32125 7685 32125 7845
rect 32125 7685 32290 7845
rect 32290 7685 32291 7845
rect 60836 7692 60836 7852
rect 60836 7692 61001 7852
rect 61001 7692 61002 7852
rect 83771 7693 83771 7853
rect 83771 7693 83936 7853
rect 83936 7693 83937 7853
rect 83771 7693 83937 7693
rect 90271 7693 90271 7853
rect 90271 7693 90436 7853
rect 90436 7693 90437 7853
rect 90271 7693 90437 7693
rect 94771 7693 94771 7853
rect 94771 7693 94936 7853
rect 94936 7693 94937 7853
rect 94771 7693 94937 7693
rect 99271 7693 99271 7853
rect 99271 7693 99436 7853
rect 99436 7693 99437 7853
rect 99271 7693 99437 7693
rect 102271 7693 102271 7853
rect 102271 7693 102436 7853
rect 102436 7693 102437 7853
rect 102271 7693 102437 7693
rect 105771 7693 105771 7853
rect 105771 7693 105936 7853
rect 105936 7693 105937 7853
rect 105771 7693 105937 7693
rect 111771 7693 111771 7853
rect 111771 7693 111936 7853
rect 111936 7693 111937 7853
rect 111771 7693 111937 7693
rect 116271 7693 116271 7853
rect 116271 7693 116436 7853
rect 116436 7693 116437 7853
rect 116271 7693 116437 7693
rect 119271 7693 119271 7853
rect 119271 7693 119436 7853
rect 119436 7693 119437 7853
rect 119271 7693 119437 7693
rect 125271 7693 125271 7853
rect 125271 7693 125436 7853
rect 125436 7693 125437 7853
rect 125271 7693 125437 7693
rect 131971 7693 131971 7853
rect 131971 7693 132136 7853
rect 132136 7693 132137 7853
rect 131971 7693 132137 7693
rect 134971 7693 134971 7853
rect 134971 7693 135136 7853
rect 135136 7693 135137 7853
rect 134971 7693 135137 7693
rect 136471 7693 136471 7853
rect 136471 7693 136636 7853
rect 136636 7693 136637 7853
rect 136471 7693 136637 7693
rect 137971 7693 137971 7853
rect 137971 7693 138136 7853
rect 138136 7693 138137 7853
rect 137971 7693 138137 7693
rect 140971 7693 140971 7853
rect 140971 7693 141136 7853
rect 141136 7693 141137 7853
rect 140971 7693 141137 7693
rect 142971 7693 142971 7853
rect 142971 7693 143136 7853
rect 143136 7693 143137 7853
rect 142971 7693 143137 7693
rect 146971 7693 146971 7853
rect 146971 7693 147136 7853
rect 147136 7693 147137 7853
rect 146971 7693 147137 7693
rect 148471 7693 148471 7853
rect 148471 7693 148636 7853
rect 148636 7693 148637 7853
rect 148471 7693 148637 7693
rect 149971 7693 149971 7853
rect 149971 7693 150136 7853
rect 150136 7693 150137 7853
rect 149971 7693 150137 7693
rect 151471 7693 151471 7853
rect 151471 7693 151636 7853
rect 151636 7693 151637 7853
rect 151471 7693 151637 7693
rect 60836 7692 61002 7692
rect 151933 7686 152093 7846
rect 32125 7685 32291 7685
rect 16454 7681 16620 7681
<< metal5 >>
rect -1473 163271 -1313 163282
rect -763 163271 -603 163282
rect -1473 163111 152927 163271
rect -2773 161038 -2589 161050
rect -2773 160878 -2761 161038
rect -2601 160878 -2589 161038
rect -2773 160866 -2589 160878
rect -3159 160060 -2975 160072
rect -3159 159900 -3147 160060
rect -2987 159900 -2975 160060
rect -3159 159888 -2975 159900
rect -1893 160060 -1709 160072
rect -1473 160060 -1313 163111
rect -763 163034 -603 163111
rect -763 162318 -603 162342
rect 151224 162318 151384 162497
rect -964 162299 152217 162318
rect -964 162158 151224 162299
rect -1893 159900 -1881 160060
rect -1721 159991 -1313 160060
rect -1721 159900 -1497 159991
rect -1893 159888 -1709 159900
rect -1509 159831 -1497 159900
rect -1337 159831 -1313 159991
rect -1509 159819 -1313 159831
rect -2773 159538 -2589 159550
rect -2773 159378 -2761 159538
rect -2601 159378 -2589 159538
rect -2773 159366 -2589 159378
rect -3159 158560 -2975 158572
rect -3159 158400 -3147 158560
rect -2987 158400 -2975 158560
rect -3159 158388 -2975 158400
rect -1893 158560 -1709 158572
rect -1473 158560 -1313 159819
rect -1893 158400 -1881 158560
rect -1721 158491 -1313 158560
rect -1721 158400 -1497 158491
rect -1893 158388 -1709 158400
rect -1509 158331 -1497 158400
rect -1337 158331 -1313 158491
rect -763 161026 -603 162158
rect 151212 162139 151224 162158
rect 151384 162158 152217 162299
rect 151384 162139 151396 162158
rect 151212 162127 151396 162139
rect -763 160890 -751 161026
rect -615 160890 -603 161026
rect -763 159526 -603 160890
rect -763 159390 -751 159526
rect -615 159390 -603 159526
rect -763 158480 -603 159390
rect -1509 158319 -1313 158331
rect -764 158320 -603 158480
rect -2773 158038 -2589 158050
rect -2773 157878 -2761 158038
rect -2601 157878 -2589 158038
rect -2773 157866 -2589 157878
rect -3159 157060 -2975 157072
rect -3159 156900 -3147 157060
rect -2987 156900 -2975 157060
rect -3159 156888 -2975 156900
rect -1893 157060 -1709 157072
rect -1473 157060 -1313 158319
rect -1893 156900 -1881 157060
rect -1721 156991 -1313 157060
rect -1721 156900 -1497 156991
rect -1893 156888 -1709 156900
rect -1509 156831 -1497 156900
rect -1337 156831 -1313 156991
rect -763 158026 -603 158320
rect -763 157890 -751 158026
rect -615 157890 -603 158026
rect -763 156980 -603 157890
rect -1509 156819 -1313 156831
rect -764 156820 -603 156980
rect -2773 156538 -2589 156550
rect -2773 156378 -2761 156538
rect -2601 156378 -2589 156538
rect -2773 156366 -2589 156378
rect -3159 155560 -2975 155572
rect -3159 155400 -3147 155560
rect -2987 155400 -2975 155560
rect -3159 155388 -2975 155400
rect -1893 155560 -1709 155572
rect -1473 155560 -1313 156819
rect -1893 155400 -1881 155560
rect -1721 155491 -1313 155560
rect -1721 155400 -1497 155491
rect -1893 155388 -1709 155400
rect -1509 155331 -1497 155400
rect -1337 155331 -1313 155491
rect -763 156526 -603 156820
rect -763 156390 -751 156526
rect -615 156390 -603 156526
rect -763 155480 -603 156390
rect -1509 155319 -1313 155331
rect -764 155320 -603 155480
rect -2773 155038 -2589 155050
rect -2773 154878 -2761 155038
rect -2601 154878 -2589 155038
rect -2773 154866 -2589 154878
rect -3159 154060 -2975 154072
rect -3159 153900 -3147 154060
rect -2987 153900 -2975 154060
rect -3159 153888 -2975 153900
rect -1893 154060 -1709 154072
rect -1473 154060 -1313 155319
rect -1893 153900 -1881 154060
rect -1721 153991 -1313 154060
rect -1721 153900 -1497 153991
rect -1893 153888 -1709 153900
rect -1509 153831 -1497 153900
rect -1337 153831 -1313 153991
rect -763 155026 -603 155320
rect -763 154890 -751 155026
rect -615 154890 -603 155026
rect -763 153980 -603 154890
rect -1509 153819 -1313 153831
rect -764 153820 -603 153980
rect -2773 153538 -2589 153550
rect -2773 153378 -2761 153538
rect -2601 153378 -2589 153538
rect -2773 153366 -2589 153378
rect -3159 152560 -2975 152572
rect -3159 152400 -3147 152560
rect -2987 152400 -2975 152560
rect -3159 152388 -2975 152400
rect -1893 152560 -1709 152572
rect -1473 152560 -1313 153819
rect -1893 152400 -1881 152560
rect -1721 152491 -1313 152560
rect -1721 152400 -1497 152491
rect -1893 152388 -1709 152400
rect -1509 152331 -1497 152400
rect -1337 152331 -1313 152491
rect -763 153526 -603 153820
rect -763 153390 -751 153526
rect -615 153390 -603 153526
rect -763 152480 -603 153390
rect -1509 152319 -1313 152331
rect -764 152320 -603 152480
rect -2773 152038 -2589 152050
rect -2773 151878 -2761 152038
rect -2601 151878 -2589 152038
rect -2773 151866 -2589 151878
rect -3159 151060 -2975 151072
rect -3159 150900 -3147 151060
rect -2987 150900 -2975 151060
rect -3159 150888 -2975 150900
rect -1893 151060 -1709 151072
rect -1473 151060 -1313 152319
rect -1893 150900 -1881 151060
rect -1721 150991 -1313 151060
rect -1721 150900 -1497 150991
rect -1893 150888 -1709 150900
rect -1509 150831 -1497 150900
rect -1337 150831 -1313 150991
rect -763 152026 -603 152320
rect -763 151890 -751 152026
rect -615 151890 -603 152026
rect -763 150980 -603 151890
rect -1509 150819 -1313 150831
rect -764 150820 -603 150980
rect -2773 150538 -2589 150550
rect -2773 150378 -2761 150538
rect -2601 150378 -2589 150538
rect -2773 150366 -2589 150378
rect -3159 149560 -2975 149572
rect -3159 149400 -3147 149560
rect -2987 149400 -2975 149560
rect -3159 149388 -2975 149400
rect -1893 149560 -1709 149572
rect -1473 149560 -1313 150819
rect -1893 149400 -1881 149560
rect -1721 149491 -1313 149560
rect -1721 149400 -1497 149491
rect -1893 149388 -1709 149400
rect -1509 149331 -1497 149400
rect -1337 149331 -1313 149491
rect -763 150526 -603 150820
rect -763 150390 -751 150526
rect -615 150390 -603 150526
rect -763 149480 -603 150390
rect -1509 149319 -1313 149331
rect -764 149320 -603 149480
rect -2773 149038 -2589 149050
rect -2773 148878 -2761 149038
rect -2601 148878 -2589 149038
rect -2773 148866 -2589 148878
rect -3159 148060 -2975 148072
rect -3159 147900 -3147 148060
rect -2987 147900 -2975 148060
rect -3159 147888 -2975 147900
rect -1893 148060 -1709 148072
rect -1473 148060 -1313 149319
rect -1893 147900 -1881 148060
rect -1721 147991 -1313 148060
rect -1721 147900 -1497 147991
rect -1893 147888 -1709 147900
rect -1509 147831 -1497 147900
rect -1337 147831 -1313 147991
rect -763 149026 -603 149320
rect -763 148890 -751 149026
rect -615 148890 -603 149026
rect -763 147980 -603 148890
rect -1509 147819 -1313 147831
rect -764 147820 -603 147980
rect -2773 147538 -2589 147550
rect -2773 147378 -2761 147538
rect -2601 147378 -2589 147538
rect -2773 147366 -2589 147378
rect -3159 146560 -2975 146572
rect -3159 146400 -3147 146560
rect -2987 146400 -2975 146560
rect -3159 146388 -2975 146400
rect -1893 146560 -1709 146572
rect -1473 146560 -1313 147819
rect -1893 146400 -1881 146560
rect -1721 146491 -1313 146560
rect -1721 146400 -1497 146491
rect -1893 146388 -1709 146400
rect -1509 146331 -1497 146400
rect -1337 146331 -1313 146491
rect -763 147526 -603 147820
rect -763 147390 -751 147526
rect -615 147390 -603 147526
rect -763 146480 -603 147390
rect -1509 146319 -1313 146331
rect -764 146320 -603 146480
rect -2773 146038 -2589 146050
rect -2773 145878 -2761 146038
rect -2601 145878 -2589 146038
rect -2773 145866 -2589 145878
rect -3159 145060 -2975 145072
rect -3159 144900 -3147 145060
rect -2987 144900 -2975 145060
rect -3159 144888 -2975 144900
rect -1893 145060 -1709 145072
rect -1473 145060 -1313 146319
rect -1893 144900 -1881 145060
rect -1721 144991 -1313 145060
rect -1721 144900 -1497 144991
rect -1893 144888 -1709 144900
rect -1509 144831 -1497 144900
rect -1337 144831 -1313 144991
rect -763 146026 -603 146320
rect -763 145890 -751 146026
rect -615 145890 -603 146026
rect -763 144980 -603 145890
rect -1509 144819 -1313 144831
rect -764 144820 -603 144980
rect -2773 144538 -2589 144550
rect -2773 144378 -2761 144538
rect -2601 144378 -2589 144538
rect -2773 144366 -2589 144378
rect -3159 143560 -2975 143572
rect -3159 143400 -3147 143560
rect -2987 143400 -2975 143560
rect -3159 143388 -2975 143400
rect -1893 143560 -1709 143572
rect -1473 143560 -1313 144819
rect -1893 143400 -1881 143560
rect -1721 143491 -1313 143560
rect -1721 143400 -1497 143491
rect -1893 143388 -1709 143400
rect -1509 143331 -1497 143400
rect -1337 143331 -1313 143491
rect -763 144526 -603 144820
rect -763 144390 -751 144526
rect -615 144390 -603 144526
rect -763 143480 -603 144390
rect -1509 143319 -1313 143331
rect -764 143320 -603 143480
rect -2773 143038 -2589 143050
rect -2773 142878 -2761 143038
rect -2601 142878 -2589 143038
rect -2773 142866 -2589 142878
rect -3159 142060 -2975 142072
rect -3159 141900 -3147 142060
rect -2987 141900 -2975 142060
rect -3159 141888 -2975 141900
rect -1893 142060 -1709 142072
rect -1473 142060 -1313 143319
rect -1893 141900 -1881 142060
rect -1721 141991 -1313 142060
rect -1721 141900 -1497 141991
rect -1893 141888 -1709 141900
rect -1509 141831 -1497 141900
rect -1337 141831 -1313 141991
rect -763 143026 -603 143320
rect -763 142890 -751 143026
rect -615 142890 -603 143026
rect -763 141980 -603 142890
rect -1509 141819 -1313 141831
rect -764 141820 -603 141980
rect -2773 141538 -2589 141550
rect -2773 141378 -2761 141538
rect -2601 141378 -2589 141538
rect -2773 141366 -2589 141378
rect -3159 140560 -2975 140572
rect -3159 140400 -3147 140560
rect -2987 140400 -2975 140560
rect -3159 140388 -2975 140400
rect -1893 140560 -1709 140572
rect -1473 140560 -1313 141819
rect -1893 140400 -1881 140560
rect -1721 140491 -1313 140560
rect -1721 140400 -1497 140491
rect -1893 140388 -1709 140400
rect -1509 140331 -1497 140400
rect -1337 140331 -1313 140491
rect -763 141526 -603 141820
rect -763 141390 -751 141526
rect -615 141390 -603 141526
rect -763 140480 -603 141390
rect -1509 140319 -1313 140331
rect -764 140320 -603 140480
rect -2773 140038 -2589 140050
rect -2773 139878 -2761 140038
rect -2601 139878 -2589 140038
rect -2773 139866 -2589 139878
rect -3159 139060 -2975 139072
rect -3159 138900 -3147 139060
rect -2987 138900 -2975 139060
rect -3159 138888 -2975 138900
rect -1893 139060 -1709 139072
rect -1473 139060 -1313 140319
rect -1893 138900 -1881 139060
rect -1721 138991 -1313 139060
rect -1721 138900 -1497 138991
rect -1893 138888 -1709 138900
rect -1509 138831 -1497 138900
rect -1337 138831 -1313 138991
rect -763 140026 -603 140320
rect -763 139890 -751 140026
rect -615 139890 -603 140026
rect -763 138980 -603 139890
rect -1509 138819 -1313 138831
rect -764 138820 -603 138980
rect -2773 138538 -2589 138550
rect -2773 138378 -2761 138538
rect -2601 138378 -2589 138538
rect -2773 138366 -2589 138378
rect -3159 137560 -2975 137572
rect -3159 137400 -3147 137560
rect -2987 137400 -2975 137560
rect -3159 137388 -2975 137400
rect -1893 137560 -1709 137572
rect -1473 137560 -1313 138819
rect -1893 137400 -1881 137560
rect -1721 137491 -1313 137560
rect -1721 137400 -1497 137491
rect -1893 137388 -1709 137400
rect -1509 137331 -1497 137400
rect -1337 137331 -1313 137491
rect -763 138526 -603 138820
rect -763 138390 -751 138526
rect -615 138390 -603 138526
rect -763 137480 -603 138390
rect -1509 137319 -1313 137331
rect -764 137320 -603 137480
rect -2773 137038 -2589 137050
rect -2773 136878 -2761 137038
rect -2601 136878 -2589 137038
rect -2773 136866 -2589 136878
rect -3159 136060 -2975 136072
rect -3159 135900 -3147 136060
rect -2987 135900 -2975 136060
rect -3159 135888 -2975 135900
rect -1893 136060 -1709 136072
rect -1473 136060 -1313 137319
rect -1893 135900 -1881 136060
rect -1721 135991 -1313 136060
rect -1721 135900 -1497 135991
rect -1893 135888 -1709 135900
rect -1509 135831 -1497 135900
rect -1337 135831 -1313 135991
rect -763 137026 -603 137320
rect -763 136890 -751 137026
rect -615 136890 -603 137026
rect -763 135980 -603 136890
rect -1509 135819 -1313 135831
rect -764 135820 -603 135980
rect -2773 135538 -2589 135550
rect -2773 135378 -2761 135538
rect -2601 135378 -2589 135538
rect -2773 135366 -2589 135378
rect -3159 134560 -2975 134572
rect -3159 134400 -3147 134560
rect -2987 134400 -2975 134560
rect -3159 134388 -2975 134400
rect -1893 134560 -1709 134572
rect -1473 134560 -1313 135819
rect -1893 134400 -1881 134560
rect -1721 134491 -1313 134560
rect -1721 134400 -1497 134491
rect -1893 134388 -1709 134400
rect -1509 134331 -1497 134400
rect -1337 134331 -1313 134491
rect -763 135526 -603 135820
rect -763 135390 -751 135526
rect -615 135390 -603 135526
rect -763 134480 -603 135390
rect -1509 134319 -1313 134331
rect -764 134320 -603 134480
rect -2773 134038 -2589 134050
rect -2773 133878 -2761 134038
rect -2601 133878 -2589 134038
rect -2773 133866 -2589 133878
rect -3159 133060 -2975 133072
rect -3159 132900 -3147 133060
rect -2987 132900 -2975 133060
rect -3159 132888 -2975 132900
rect -1893 133060 -1709 133072
rect -1473 133060 -1313 134319
rect -1893 132900 -1881 133060
rect -1721 132991 -1313 133060
rect -1721 132900 -1497 132991
rect -1893 132888 -1709 132900
rect -1509 132831 -1497 132900
rect -1337 132831 -1313 132991
rect -763 134026 -603 134320
rect -763 133890 -751 134026
rect -615 133890 -603 134026
rect -763 132980 -603 133890
rect -1509 132819 -1313 132831
rect -764 132820 -603 132980
rect -2773 132538 -2589 132550
rect -2773 132378 -2761 132538
rect -2601 132378 -2589 132538
rect -2773 132366 -2589 132378
rect -3159 131560 -2975 131572
rect -3159 131400 -3147 131560
rect -2987 131400 -2975 131560
rect -3159 131388 -2975 131400
rect -1893 131560 -1709 131572
rect -1473 131560 -1313 132819
rect -1893 131400 -1881 131560
rect -1721 131491 -1313 131560
rect -1721 131400 -1497 131491
rect -1893 131388 -1709 131400
rect -1509 131331 -1497 131400
rect -1337 131331 -1313 131491
rect -763 132526 -603 132820
rect -763 132390 -751 132526
rect -615 132390 -603 132526
rect -763 131480 -603 132390
rect -1509 131319 -1313 131331
rect -764 131320 -603 131480
rect -2773 131038 -2589 131050
rect -2773 130878 -2761 131038
rect -2601 130878 -2589 131038
rect -2773 130866 -2589 130878
rect -3159 130060 -2975 130072
rect -3159 129900 -3147 130060
rect -2987 129900 -2975 130060
rect -3159 129888 -2975 129900
rect -1893 130060 -1709 130072
rect -1473 130060 -1313 131319
rect -1893 129900 -1881 130060
rect -1721 129991 -1313 130060
rect -1721 129900 -1497 129991
rect -1893 129888 -1709 129900
rect -1509 129831 -1497 129900
rect -1337 129831 -1313 129991
rect -763 131026 -603 131320
rect -763 130890 -751 131026
rect -615 130890 -603 131026
rect -763 129980 -603 130890
rect -1509 129819 -1313 129831
rect -764 129820 -603 129980
rect -2773 129538 -2589 129550
rect -2773 129378 -2761 129538
rect -2601 129378 -2589 129538
rect -2773 129366 -2589 129378
rect -3159 128560 -2975 128572
rect -3159 128400 -3147 128560
rect -2987 128400 -2975 128560
rect -3159 128388 -2975 128400
rect -1893 128560 -1709 128572
rect -1473 128560 -1313 129819
rect -1893 128400 -1881 128560
rect -1721 128491 -1313 128560
rect -1721 128400 -1497 128491
rect -1893 128388 -1709 128400
rect -1509 128331 -1497 128400
rect -1337 128331 -1313 128491
rect -763 129526 -603 129820
rect -763 129390 -751 129526
rect -615 129390 -603 129526
rect -763 128480 -603 129390
rect -1509 128319 -1313 128331
rect -764 128320 -603 128480
rect -2773 128038 -2589 128050
rect -2773 127878 -2761 128038
rect -2601 127878 -2589 128038
rect -2773 127866 -2589 127878
rect -3159 127060 -2975 127072
rect -3159 126900 -3147 127060
rect -2987 126900 -2975 127060
rect -3159 126888 -2975 126900
rect -1893 127060 -1709 127072
rect -1473 127060 -1313 128319
rect -1893 126900 -1881 127060
rect -1721 126991 -1313 127060
rect -1721 126900 -1497 126991
rect -1893 126888 -1709 126900
rect -1509 126831 -1497 126900
rect -1337 126831 -1313 126991
rect -763 128026 -603 128320
rect -763 127890 -751 128026
rect -615 127890 -603 128026
rect -763 126980 -603 127890
rect -1509 126819 -1313 126831
rect -764 126820 -603 126980
rect -2773 126538 -2589 126550
rect -2773 126378 -2761 126538
rect -2601 126378 -2589 126538
rect -2773 126366 -2589 126378
rect -3159 125560 -2975 125572
rect -3159 125400 -3147 125560
rect -2987 125400 -2975 125560
rect -3159 125388 -2975 125400
rect -1893 125560 -1709 125572
rect -1473 125560 -1313 126819
rect -1893 125400 -1881 125560
rect -1721 125491 -1313 125560
rect -1721 125400 -1497 125491
rect -1893 125388 -1709 125400
rect -1509 125331 -1497 125400
rect -1337 125331 -1313 125491
rect -763 126526 -603 126820
rect -763 126390 -751 126526
rect -615 126390 -603 126526
rect -763 125480 -603 126390
rect -1509 125319 -1313 125331
rect -764 125320 -603 125480
rect -2773 125038 -2589 125050
rect -2773 124878 -2761 125038
rect -2601 124878 -2589 125038
rect -2773 124866 -2589 124878
rect -3159 124060 -2975 124072
rect -3159 123900 -3147 124060
rect -2987 123900 -2975 124060
rect -3159 123888 -2975 123900
rect -1893 124060 -1709 124072
rect -1473 124060 -1313 125319
rect -1893 123900 -1881 124060
rect -1721 123991 -1313 124060
rect -1721 123900 -1497 123991
rect -1893 123888 -1709 123900
rect -1509 123831 -1497 123900
rect -1337 123831 -1313 123991
rect -763 125026 -603 125320
rect -763 124890 -751 125026
rect -615 124890 -603 125026
rect -763 123980 -603 124890
rect -1509 123819 -1313 123831
rect -764 123820 -603 123980
rect -3159 122560 -2975 122572
rect -3159 122400 -3147 122560
rect -2987 122400 -2975 122560
rect -3159 122388 -2975 122400
rect -1893 122560 -1709 122572
rect -1473 122560 -1313 123819
rect -1893 122400 -1881 122560
rect -1721 122491 -1313 122560
rect -1721 122400 -1497 122491
rect -1893 122388 -1709 122400
rect -1509 122331 -1497 122400
rect -1337 122331 -1313 122491
rect -763 122480 -603 123820
rect -1509 122319 -1313 122331
rect -764 122320 -603 122480
rect -2773 122038 -2589 122050
rect -2773 121878 -2761 122038
rect -2601 121878 -2589 122038
rect -2773 121866 -2589 121878
rect -3159 121060 -2975 121072
rect -3159 120900 -3147 121060
rect -2987 120900 -2975 121060
rect -3159 120888 -2975 120900
rect -1893 121060 -1709 121072
rect -1473 121060 -1313 122319
rect -1893 120900 -1881 121060
rect -1721 120991 -1313 121060
rect -1721 120900 -1497 120991
rect -1893 120888 -1709 120900
rect -1509 120831 -1497 120900
rect -1337 120831 -1313 120991
rect -763 122026 -603 122320
rect -763 121890 -751 122026
rect -615 121890 -603 122026
rect -763 120980 -603 121890
rect -1509 120819 -1313 120831
rect -764 120820 -603 120980
rect -2773 120538 -2589 120550
rect -2773 120378 -2761 120538
rect -2601 120378 -2589 120538
rect -2773 120366 -2589 120378
rect -3159 119560 -2975 119572
rect -3159 119400 -3147 119560
rect -2987 119400 -2975 119560
rect -3159 119388 -2975 119400
rect -1893 119560 -1709 119572
rect -1473 119560 -1313 120819
rect -1893 119400 -1881 119560
rect -1721 119491 -1313 119560
rect -1721 119400 -1497 119491
rect -1893 119388 -1709 119400
rect -1509 119331 -1497 119400
rect -1337 119331 -1313 119491
rect -763 120526 -603 120820
rect -763 120390 -751 120526
rect -615 120390 -603 120526
rect -763 119480 -603 120390
rect -1509 119319 -1313 119331
rect -764 119320 -603 119480
rect -2773 119038 -2589 119050
rect -2773 118878 -2761 119038
rect -2601 118878 -2589 119038
rect -2773 118866 -2589 118878
rect -3159 118060 -2975 118072
rect -3159 117900 -3147 118060
rect -2987 117900 -2975 118060
rect -3159 117888 -2975 117900
rect -1893 118060 -1709 118072
rect -1473 118060 -1313 119319
rect -1893 117900 -1881 118060
rect -1721 117991 -1313 118060
rect -1721 117900 -1497 117991
rect -1893 117888 -1709 117900
rect -1509 117831 -1497 117900
rect -1337 117831 -1313 117991
rect -763 119026 -603 119320
rect -763 118890 -751 119026
rect -615 118890 -603 119026
rect -763 117980 -603 118890
rect -1509 117819 -1313 117831
rect -764 117820 -603 117980
rect -2773 117538 -2589 117550
rect -2773 117378 -2761 117538
rect -2601 117378 -2589 117538
rect -2773 117366 -2589 117378
rect -3159 116560 -2975 116572
rect -3159 116400 -3147 116560
rect -2987 116400 -2975 116560
rect -3159 116388 -2975 116400
rect -1893 116560 -1709 116572
rect -1473 116560 -1313 117819
rect -1893 116400 -1881 116560
rect -1721 116491 -1313 116560
rect -1721 116400 -1497 116491
rect -1893 116388 -1709 116400
rect -1509 116331 -1497 116400
rect -1337 116331 -1313 116491
rect -763 117526 -603 117820
rect -763 117390 -751 117526
rect -615 117390 -603 117526
rect -763 116480 -603 117390
rect -1509 116319 -1313 116331
rect -764 116320 -603 116480
rect -2773 116038 -2589 116050
rect -2773 115878 -2761 116038
rect -2601 115878 -2589 116038
rect -2773 115866 -2589 115878
rect -3159 115060 -2975 115072
rect -3159 114900 -3147 115060
rect -2987 114900 -2975 115060
rect -3159 114888 -2975 114900
rect -1893 115060 -1709 115072
rect -1473 115060 -1313 116319
rect -1893 114900 -1881 115060
rect -1721 114991 -1313 115060
rect -1721 114900 -1497 114991
rect -1893 114888 -1709 114900
rect -1509 114831 -1497 114900
rect -1337 114831 -1313 114991
rect -763 116026 -603 116320
rect -763 115890 -751 116026
rect -615 115890 -603 116026
rect -763 114980 -603 115890
rect -1509 114819 -1313 114831
rect -764 114820 -603 114980
rect -2773 114538 -2589 114550
rect -2773 114378 -2761 114538
rect -2601 114378 -2589 114538
rect -2773 114366 -2589 114378
rect -3159 113560 -2975 113572
rect -3159 113400 -3147 113560
rect -2987 113400 -2975 113560
rect -3159 113388 -2975 113400
rect -1893 113560 -1709 113572
rect -1473 113560 -1313 114819
rect -1893 113400 -1881 113560
rect -1721 113491 -1313 113560
rect -1721 113400 -1497 113491
rect -1893 113388 -1709 113400
rect -1509 113331 -1497 113400
rect -1337 113331 -1313 113491
rect -763 114526 -603 114820
rect -763 114390 -751 114526
rect -615 114390 -603 114526
rect -763 113480 -603 114390
rect -1509 113319 -1313 113331
rect -764 113320 -603 113480
rect -2773 113038 -2589 113050
rect -2773 112878 -2761 113038
rect -2601 112878 -2589 113038
rect -2773 112866 -2589 112878
rect -3159 112060 -2975 112072
rect -3159 111900 -3147 112060
rect -2987 111900 -2975 112060
rect -3159 111888 -2975 111900
rect -1893 112060 -1709 112072
rect -1473 112060 -1313 113319
rect -1893 111900 -1881 112060
rect -1721 111991 -1313 112060
rect -1721 111900 -1497 111991
rect -1893 111888 -1709 111900
rect -1509 111831 -1497 111900
rect -1337 111831 -1313 111991
rect -763 113026 -603 113320
rect -763 112890 -751 113026
rect -615 112890 -603 113026
rect -763 111980 -603 112890
rect -1509 111819 -1313 111831
rect -764 111820 -603 111980
rect -2773 111538 -2589 111550
rect -2773 111378 -2761 111538
rect -2601 111378 -2589 111538
rect -2773 111366 -2589 111378
rect -3159 110560 -2975 110572
rect -3159 110400 -3147 110560
rect -2987 110400 -2975 110560
rect -3159 110388 -2975 110400
rect -1893 110560 -1709 110572
rect -1473 110560 -1313 111819
rect -1893 110400 -1881 110560
rect -1721 110491 -1313 110560
rect -1721 110400 -1497 110491
rect -1893 110388 -1709 110400
rect -1509 110331 -1497 110400
rect -1337 110331 -1313 110491
rect -763 111526 -603 111820
rect -763 111390 -751 111526
rect -615 111390 -603 111526
rect -763 110480 -603 111390
rect -1509 110319 -1313 110331
rect -764 110320 -603 110480
rect -2773 110038 -2589 110050
rect -2773 109878 -2761 110038
rect -2601 109878 -2589 110038
rect -2773 109866 -2589 109878
rect -3159 109060 -2975 109072
rect -3159 108900 -3147 109060
rect -2987 108900 -2975 109060
rect -3159 108888 -2975 108900
rect -1893 109060 -1709 109072
rect -1473 109060 -1313 110319
rect -1893 108900 -1881 109060
rect -1721 108991 -1313 109060
rect -1721 108900 -1497 108991
rect -1893 108888 -1709 108900
rect -1509 108831 -1497 108900
rect -1337 108831 -1313 108991
rect -763 110026 -603 110320
rect -763 109890 -751 110026
rect -615 109890 -603 110026
rect -763 108980 -603 109890
rect -1509 108819 -1313 108831
rect -764 108820 -603 108980
rect -2773 108538 -2589 108550
rect -2773 108378 -2761 108538
rect -2601 108378 -2589 108538
rect -2773 108366 -2589 108378
rect -3159 107560 -2975 107572
rect -3159 107400 -3147 107560
rect -2987 107400 -2975 107560
rect -3159 107388 -2975 107400
rect -1893 107560 -1709 107572
rect -1473 107560 -1313 108819
rect -1893 107400 -1881 107560
rect -1721 107491 -1313 107560
rect -1721 107400 -1497 107491
rect -1893 107388 -1709 107400
rect -1509 107331 -1497 107400
rect -1337 107331 -1313 107491
rect -763 108526 -603 108820
rect -763 108390 -751 108526
rect -615 108390 -603 108526
rect -763 107480 -603 108390
rect -1509 107319 -1313 107331
rect -764 107320 -603 107480
rect -2773 107038 -2589 107050
rect -2773 106878 -2761 107038
rect -2601 106878 -2589 107038
rect -2773 106866 -2589 106878
rect -3159 106060 -2975 106072
rect -3159 105900 -3147 106060
rect -2987 105900 -2975 106060
rect -3159 105888 -2975 105900
rect -1893 106060 -1709 106072
rect -1473 106060 -1313 107319
rect -1893 105900 -1881 106060
rect -1721 105991 -1313 106060
rect -1721 105900 -1497 105991
rect -1893 105888 -1709 105900
rect -1509 105831 -1497 105900
rect -1337 105831 -1313 105991
rect -763 107026 -603 107320
rect -763 106890 -751 107026
rect -615 106890 -603 107026
rect -763 105980 -603 106890
rect -1509 105819 -1313 105831
rect -764 105820 -603 105980
rect -2773 105538 -2589 105550
rect -2773 105378 -2761 105538
rect -2601 105378 -2589 105538
rect -2773 105366 -2589 105378
rect -1473 104560 -1313 105819
rect -1560 104491 -1313 104560
rect -1560 104400 -1497 104491
rect -1509 104331 -1497 104400
rect -1337 104331 -1313 104491
rect -763 105526 -603 105820
rect -763 105390 -751 105526
rect -615 105390 -603 105526
rect -763 104480 -603 105390
rect -1509 104319 -1313 104331
rect -764 104320 -603 104480
rect -2773 104038 -2589 104050
rect -2773 103878 -2761 104038
rect -2601 103878 -2589 104038
rect -2773 103866 -2589 103878
rect -3159 103060 -2975 103072
rect -3159 102900 -3147 103060
rect -2987 102900 -2975 103060
rect -3159 102888 -2975 102900
rect -1893 103060 -1709 103072
rect -1473 103060 -1313 104319
rect -1893 102900 -1881 103060
rect -1721 102991 -1313 103060
rect -1721 102900 -1497 102991
rect -1893 102888 -1709 102900
rect -1509 102831 -1497 102900
rect -1337 102831 -1313 102991
rect -763 104026 -603 104320
rect -763 103890 -751 104026
rect -615 103890 -603 104026
rect -763 102980 -603 103890
rect -1509 102819 -1313 102831
rect -764 102820 -603 102980
rect -2773 102538 -2589 102550
rect -2773 102378 -2761 102538
rect -2601 102378 -2589 102538
rect -2773 102366 -2589 102378
rect -3159 101560 -2975 101572
rect -3159 101400 -3147 101560
rect -2987 101400 -2975 101560
rect -3159 101388 -2975 101400
rect -1893 101560 -1709 101572
rect -1473 101560 -1313 102819
rect -1893 101400 -1881 101560
rect -1721 101491 -1313 101560
rect -1721 101400 -1497 101491
rect -1893 101388 -1709 101400
rect -1509 101331 -1497 101400
rect -1337 101331 -1313 101491
rect -763 102526 -603 102820
rect -763 102390 -751 102526
rect -615 102390 -603 102526
rect -763 101480 -603 102390
rect -1509 101319 -1313 101331
rect -764 101320 -603 101480
rect -2773 101038 -2589 101050
rect -2773 100878 -2761 101038
rect -2601 100878 -2589 101038
rect -2773 100866 -2589 100878
rect -3159 100060 -2975 100072
rect -3159 99900 -3147 100060
rect -2987 99900 -2975 100060
rect -3159 99888 -2975 99900
rect -1893 100060 -1709 100072
rect -1473 100060 -1313 101319
rect -1893 99900 -1881 100060
rect -1721 99991 -1313 100060
rect -1721 99900 -1497 99991
rect -1893 99888 -1709 99900
rect -1509 99831 -1497 99900
rect -1337 99831 -1313 99991
rect -763 101026 -603 101320
rect -763 100890 -751 101026
rect -615 100890 -603 101026
rect -763 99980 -603 100890
rect -1509 99819 -1313 99831
rect -764 99820 -603 99980
rect -2773 99538 -2589 99550
rect -2773 99378 -2761 99538
rect -2601 99378 -2589 99538
rect -2773 99366 -2589 99378
rect -3159 98560 -2975 98572
rect -3159 98400 -3147 98560
rect -2987 98400 -2975 98560
rect -3159 98388 -2975 98400
rect -1893 98560 -1709 98572
rect -1473 98560 -1313 99819
rect -1893 98400 -1881 98560
rect -1721 98491 -1313 98560
rect -1721 98400 -1497 98491
rect -1893 98388 -1709 98400
rect -1509 98331 -1497 98400
rect -1337 98331 -1313 98491
rect -763 99526 -603 99820
rect -763 99390 -751 99526
rect -615 99390 -603 99526
rect -763 98480 -603 99390
rect -1509 98319 -1313 98331
rect -764 98320 -603 98480
rect -2773 98038 -2589 98050
rect -2773 97878 -2761 98038
rect -2601 97878 -2589 98038
rect -2773 97866 -2589 97878
rect -3159 97060 -2975 97072
rect -3159 96900 -3147 97060
rect -2987 96900 -2975 97060
rect -3159 96888 -2975 96900
rect -1893 97060 -1709 97072
rect -1473 97060 -1313 98319
rect -1893 96900 -1881 97060
rect -1721 96991 -1313 97060
rect -1721 96900 -1497 96991
rect -1893 96888 -1709 96900
rect -1509 96831 -1497 96900
rect -1337 96831 -1313 96991
rect -763 98026 -603 98320
rect -763 97890 -751 98026
rect -615 97890 -603 98026
rect -763 96980 -603 97890
rect -1509 96819 -1313 96831
rect -764 96820 -603 96980
rect -2773 96538 -2589 96550
rect -2773 96378 -2761 96538
rect -2601 96378 -2589 96538
rect -2773 96366 -2589 96378
rect -3159 95560 -2975 95572
rect -3159 95400 -3147 95560
rect -2987 95400 -2975 95560
rect -3159 95388 -2975 95400
rect -1893 95560 -1709 95572
rect -1473 95560 -1313 96819
rect -1893 95400 -1881 95560
rect -1721 95491 -1313 95560
rect -1721 95400 -1497 95491
rect -1893 95388 -1709 95400
rect -1509 95331 -1497 95400
rect -1337 95331 -1313 95491
rect -763 96526 -603 96820
rect -763 96390 -751 96526
rect -615 96390 -603 96526
rect -763 95480 -603 96390
rect -1509 95319 -1313 95331
rect -764 95320 -603 95480
rect -2773 95038 -2589 95050
rect -2773 94878 -2761 95038
rect -2601 94878 -2589 95038
rect -2773 94866 -2589 94878
rect -3159 94060 -2975 94072
rect -3159 93900 -3147 94060
rect -2987 93900 -2975 94060
rect -3159 93888 -2975 93900
rect -1893 94060 -1709 94072
rect -1473 94060 -1313 95319
rect -1893 93900 -1881 94060
rect -1721 93991 -1313 94060
rect -1721 93900 -1497 93991
rect -1893 93888 -1709 93900
rect -1509 93831 -1497 93900
rect -1337 93831 -1313 93991
rect -763 95026 -603 95320
rect -763 94890 -751 95026
rect -615 94890 -603 95026
rect -763 93980 -603 94890
rect -1509 93819 -1313 93831
rect -764 93820 -603 93980
rect -2773 93538 -2589 93550
rect -2773 93378 -2761 93538
rect -2601 93378 -2589 93538
rect -2773 93366 -2589 93378
rect -3159 92560 -2975 92572
rect -3159 92400 -3147 92560
rect -2987 92400 -2975 92560
rect -3159 92388 -2975 92400
rect -1893 92560 -1709 92572
rect -1473 92560 -1313 93819
rect -1893 92400 -1881 92560
rect -1721 92491 -1313 92560
rect -1721 92400 -1497 92491
rect -1893 92388 -1709 92400
rect -1509 92331 -1497 92400
rect -1337 92331 -1313 92491
rect -763 93526 -603 93820
rect -763 93390 -751 93526
rect -615 93390 -603 93526
rect -763 92480 -603 93390
rect -1509 92319 -1313 92331
rect -764 92320 -603 92480
rect -2773 92038 -2589 92050
rect -2773 91878 -2761 92038
rect -2601 91878 -2589 92038
rect -2773 91866 -2589 91878
rect -3159 91060 -2975 91072
rect -3159 90900 -3147 91060
rect -2987 90900 -2975 91060
rect -3159 90888 -2975 90900
rect -1893 91060 -1709 91072
rect -1473 91060 -1313 92319
rect -1893 90900 -1881 91060
rect -1721 90991 -1313 91060
rect -1721 90900 -1497 90991
rect -1893 90888 -1709 90900
rect -1509 90831 -1497 90900
rect -1337 90831 -1313 90991
rect -763 92026 -603 92320
rect -763 91890 -751 92026
rect -615 91890 -603 92026
rect -763 90980 -603 91890
rect -1509 90819 -1313 90831
rect -764 90820 -603 90980
rect -2773 90538 -2589 90550
rect -2773 90378 -2761 90538
rect -2601 90378 -2589 90538
rect -2773 90366 -2589 90378
rect -3159 89560 -2975 89572
rect -3159 89400 -3147 89560
rect -2987 89400 -2975 89560
rect -3159 89388 -2975 89400
rect -1893 89560 -1709 89572
rect -1473 89560 -1313 90819
rect -1893 89400 -1881 89560
rect -1721 89491 -1313 89560
rect -1721 89400 -1497 89491
rect -1893 89388 -1709 89400
rect -1509 89331 -1497 89400
rect -1337 89331 -1313 89491
rect -763 90526 -603 90820
rect -763 90390 -751 90526
rect -615 90390 -603 90526
rect -763 89480 -603 90390
rect -1509 89319 -1313 89331
rect -764 89320 -603 89480
rect -2773 89038 -2589 89050
rect -2773 88878 -2761 89038
rect -2601 88878 -2589 89038
rect -2773 88866 -2589 88878
rect -3159 88060 -2975 88072
rect -3159 87900 -3147 88060
rect -2987 87900 -2975 88060
rect -3159 87888 -2975 87900
rect -1893 88060 -1709 88072
rect -1473 88060 -1313 89319
rect -1893 87900 -1881 88060
rect -1721 87991 -1313 88060
rect -1721 87900 -1497 87991
rect -1893 87888 -1709 87900
rect -1509 87831 -1497 87900
rect -1337 87831 -1313 87991
rect -763 89026 -603 89320
rect -763 88890 -751 89026
rect -615 88890 -603 89026
rect -763 87980 -603 88890
rect -1509 87819 -1313 87831
rect -764 87820 -603 87980
rect -2773 87538 -2589 87550
rect -2773 87378 -2761 87538
rect -2601 87378 -2589 87538
rect -2773 87366 -2589 87378
rect -3159 86560 -2975 86572
rect -3159 86400 -3147 86560
rect -2987 86400 -2975 86560
rect -3159 86388 -2975 86400
rect -1893 86560 -1709 86572
rect -1473 86560 -1313 87819
rect -1893 86400 -1881 86560
rect -1721 86491 -1313 86560
rect -1721 86400 -1497 86491
rect -1893 86388 -1709 86400
rect -1509 86331 -1497 86400
rect -1337 86331 -1313 86491
rect -763 87526 -603 87820
rect -763 87390 -751 87526
rect -615 87390 -603 87526
rect -763 86480 -603 87390
rect -1509 86319 -1313 86331
rect -764 86320 -603 86480
rect -2773 86038 -2589 86050
rect -2773 85878 -2761 86038
rect -2601 85878 -2589 86038
rect -2773 85866 -2589 85878
rect -3159 85060 -2975 85072
rect -3159 84900 -3147 85060
rect -2987 84900 -2975 85060
rect -3159 84888 -2975 84900
rect -1893 85060 -1709 85072
rect -1473 85060 -1313 86319
rect -1893 84900 -1881 85060
rect -1721 84991 -1313 85060
rect -1721 84900 -1497 84991
rect -1893 84888 -1709 84900
rect -1509 84831 -1497 84900
rect -1337 84831 -1313 84991
rect -763 86026 -603 86320
rect -763 85890 -751 86026
rect -615 85890 -603 86026
rect -763 84980 -603 85890
rect -1509 84819 -1313 84831
rect -764 84820 -603 84980
rect -2773 84538 -2589 84550
rect -2773 84378 -2761 84538
rect -2601 84378 -2589 84538
rect -2773 84366 -2589 84378
rect -3159 83560 -2975 83572
rect -3159 83400 -3147 83560
rect -2987 83400 -2975 83560
rect -3159 83388 -2975 83400
rect -1893 83560 -1709 83572
rect -1473 83560 -1313 84819
rect -1893 83400 -1881 83560
rect -1721 83491 -1313 83560
rect -1721 83400 -1497 83491
rect -1893 83388 -1709 83400
rect -1509 83331 -1497 83400
rect -1337 83331 -1313 83491
rect -763 84526 -603 84820
rect -763 84390 -751 84526
rect -615 84390 -603 84526
rect -763 83480 -603 84390
rect -1509 83319 -1313 83331
rect -764 83320 -603 83480
rect -2773 83038 -2589 83050
rect -2773 82878 -2761 83038
rect -2601 82878 -2589 83038
rect -2773 82866 -2589 82878
rect -3159 82060 -2975 82072
rect -3159 81900 -3147 82060
rect -2987 81900 -2975 82060
rect -3159 81888 -2975 81900
rect -1893 82060 -1709 82072
rect -1473 82060 -1313 83319
rect -1893 81900 -1881 82060
rect -1721 81991 -1313 82060
rect -1721 81900 -1497 81991
rect -1893 81888 -1709 81900
rect -1509 81831 -1497 81900
rect -1337 81831 -1313 81991
rect -763 83026 -603 83320
rect -763 82890 -751 83026
rect -615 82890 -603 83026
rect -763 81980 -603 82890
rect -1509 81819 -1313 81831
rect -764 81820 -603 81980
rect -2773 81538 -2589 81550
rect -2773 81378 -2761 81538
rect -2601 81378 -2589 81538
rect -2773 81366 -2589 81378
rect -3159 80560 -2975 80572
rect -3159 80400 -3147 80560
rect -2987 80400 -2975 80560
rect -3159 80388 -2975 80400
rect -1893 80560 -1709 80572
rect -1473 80560 -1313 81819
rect -1893 80400 -1881 80560
rect -1721 80491 -1313 80560
rect -1721 80400 -1497 80491
rect -1893 80388 -1709 80400
rect -1509 80331 -1497 80400
rect -1337 80331 -1313 80491
rect -763 81526 -603 81820
rect -763 81390 -751 81526
rect -615 81390 -603 81526
rect -763 80480 -603 81390
rect -1509 80319 -1313 80331
rect -764 80320 -603 80480
rect -2773 80038 -2589 80050
rect -2773 79878 -2761 80038
rect -2601 79878 -2589 80038
rect -2773 79866 -2589 79878
rect -3159 79060 -2975 79072
rect -3159 78900 -3147 79060
rect -2987 78900 -2975 79060
rect -3159 78888 -2975 78900
rect -1893 79060 -1709 79072
rect -1473 79060 -1313 80319
rect -1893 78900 -1881 79060
rect -1721 78991 -1313 79060
rect -1721 78900 -1497 78991
rect -1893 78888 -1709 78900
rect -1509 78831 -1497 78900
rect -1337 78831 -1313 78991
rect -763 80026 -603 80320
rect -763 79890 -751 80026
rect -615 79890 -603 80026
rect -763 78980 -603 79890
rect -1509 78819 -1313 78831
rect -764 78820 -603 78980
rect -2773 78538 -2589 78550
rect -2773 78378 -2761 78538
rect -2601 78378 -2589 78538
rect -2773 78366 -2589 78378
rect -3159 77560 -2975 77572
rect -3159 77400 -3147 77560
rect -2987 77400 -2975 77560
rect -3159 77388 -2975 77400
rect -1893 77560 -1709 77572
rect -1473 77560 -1313 78819
rect -1893 77400 -1881 77560
rect -1721 77491 -1313 77560
rect -1721 77400 -1497 77491
rect -1893 77388 -1709 77400
rect -1509 77331 -1497 77400
rect -1337 77331 -1313 77491
rect -763 78526 -603 78820
rect -763 78390 -751 78526
rect -615 78390 -603 78526
rect -763 77480 -603 78390
rect -1509 77319 -1313 77331
rect -764 77320 -603 77480
rect -2773 77038 -2589 77050
rect -2773 76878 -2761 77038
rect -2601 76878 -2589 77038
rect -2773 76866 -2589 76878
rect -3159 76060 -2975 76072
rect -3159 75900 -3147 76060
rect -2987 75900 -2975 76060
rect -3159 75888 -2975 75900
rect -1893 76060 -1709 76072
rect -1473 76060 -1313 77319
rect -1893 75900 -1881 76060
rect -1721 75991 -1313 76060
rect -1721 75900 -1497 75991
rect -1893 75888 -1709 75900
rect -1509 75831 -1497 75900
rect -1337 75831 -1313 75991
rect -763 77026 -603 77320
rect -763 76890 -751 77026
rect -615 76890 -603 77026
rect -763 75980 -603 76890
rect -1509 75819 -1313 75831
rect -764 75820 -603 75980
rect -2773 75538 -2589 75550
rect -2773 75378 -2761 75538
rect -2601 75378 -2589 75538
rect -2773 75366 -2589 75378
rect -3159 74560 -2975 74572
rect -3159 74400 -3147 74560
rect -2987 74400 -2975 74560
rect -3159 74388 -2975 74400
rect -1893 74560 -1709 74572
rect -1473 74560 -1313 75819
rect -1893 74400 -1881 74560
rect -1721 74491 -1313 74560
rect -1721 74400 -1497 74491
rect -1893 74388 -1709 74400
rect -1509 74331 -1497 74400
rect -1337 74331 -1313 74491
rect -763 75526 -603 75820
rect -763 75390 -751 75526
rect -615 75390 -603 75526
rect -763 74480 -603 75390
rect -1509 74319 -1313 74331
rect -764 74320 -603 74480
rect -2773 74038 -2589 74050
rect -2773 73878 -2761 74038
rect -2601 73878 -2589 74038
rect -2773 73866 -2589 73878
rect -3159 73060 -2975 73072
rect -3159 72900 -3147 73060
rect -2987 72900 -2975 73060
rect -3159 72888 -2975 72900
rect -1893 73060 -1709 73072
rect -1473 73060 -1313 74319
rect -1893 72900 -1881 73060
rect -1721 72991 -1313 73060
rect -1721 72900 -1497 72991
rect -1893 72888 -1709 72900
rect -1509 72831 -1497 72900
rect -1337 72831 -1313 72991
rect -763 74026 -603 74320
rect -763 73890 -751 74026
rect -615 73890 -603 74026
rect -763 72980 -603 73890
rect -1509 72819 -1313 72831
rect -764 72820 -603 72980
rect -2773 72538 -2589 72550
rect -2773 72378 -2761 72538
rect -2601 72378 -2589 72538
rect -2773 72366 -2589 72378
rect -3159 71560 -2975 71572
rect -3159 71400 -3147 71560
rect -2987 71400 -2975 71560
rect -3159 71388 -2975 71400
rect -1893 71560 -1709 71572
rect -1473 71560 -1313 72819
rect -1893 71400 -1881 71560
rect -1721 71491 -1313 71560
rect -1721 71400 -1497 71491
rect -1893 71388 -1709 71400
rect -1509 71331 -1497 71400
rect -1337 71331 -1313 71491
rect -763 72526 -603 72820
rect -763 72390 -751 72526
rect -615 72390 -603 72526
rect -763 71480 -603 72390
rect -1509 71319 -1313 71331
rect -764 71320 -603 71480
rect -2773 71038 -2589 71050
rect -2773 70878 -2761 71038
rect -2601 70878 -2589 71038
rect -2773 70866 -2589 70878
rect -3159 70060 -2975 70072
rect -3159 69900 -3147 70060
rect -2987 69900 -2975 70060
rect -3159 69888 -2975 69900
rect -1893 70060 -1709 70072
rect -1473 70060 -1313 71319
rect -1893 69900 -1881 70060
rect -1721 69991 -1313 70060
rect -1721 69900 -1497 69991
rect -1893 69888 -1709 69900
rect -1509 69831 -1497 69900
rect -1337 69831 -1313 69991
rect -763 71026 -603 71320
rect -763 70890 -751 71026
rect -615 70890 -603 71026
rect -763 69980 -603 70890
rect -1509 69819 -1313 69831
rect -764 69820 -603 69980
rect -2773 69538 -2589 69550
rect -2773 69378 -2761 69538
rect -2601 69378 -2589 69538
rect -2773 69366 -2589 69378
rect -3159 68560 -2975 68572
rect -3159 68400 -3147 68560
rect -2987 68400 -2975 68560
rect -3159 68388 -2975 68400
rect -1893 68560 -1709 68572
rect -1473 68560 -1313 69819
rect -1893 68400 -1881 68560
rect -1721 68491 -1313 68560
rect -1721 68400 -1497 68491
rect -1893 68388 -1709 68400
rect -1509 68331 -1497 68400
rect -1337 68331 -1313 68491
rect -763 69526 -603 69820
rect -763 69390 -751 69526
rect -615 69390 -603 69526
rect -763 68480 -603 69390
rect -1509 68319 -1313 68331
rect -764 68320 -603 68480
rect -2773 68038 -2589 68050
rect -2773 67878 -2761 68038
rect -2601 67878 -2589 68038
rect -2773 67866 -2589 67878
rect -3159 67060 -2975 67072
rect -3159 66900 -3147 67060
rect -2987 66900 -2975 67060
rect -3159 66888 -2975 66900
rect -1893 67060 -1709 67072
rect -1473 67060 -1313 68319
rect -1893 66900 -1881 67060
rect -1721 66991 -1313 67060
rect -1721 66900 -1497 66991
rect -1893 66888 -1709 66900
rect -1509 66831 -1497 66900
rect -1337 66831 -1313 66991
rect -763 68026 -603 68320
rect -763 67890 -751 68026
rect -615 67890 -603 68026
rect -763 66980 -603 67890
rect -1509 66819 -1313 66831
rect -764 66820 -603 66980
rect -2773 66538 -2589 66550
rect -2773 66378 -2761 66538
rect -2601 66378 -2589 66538
rect -2773 66366 -2589 66378
rect -3159 65560 -2975 65572
rect -3159 65400 -3147 65560
rect -2987 65400 -2975 65560
rect -3159 65388 -2975 65400
rect -1893 65560 -1709 65572
rect -1473 65560 -1313 66819
rect -1893 65400 -1881 65560
rect -1721 65491 -1313 65560
rect -1721 65400 -1497 65491
rect -1893 65388 -1709 65400
rect -1509 65331 -1497 65400
rect -1337 65331 -1313 65491
rect -763 66526 -603 66820
rect -763 66390 -751 66526
rect -615 66390 -603 66526
rect -763 65480 -603 66390
rect -1509 65319 -1313 65331
rect -764 65320 -603 65480
rect -2773 65038 -2589 65050
rect -2773 64878 -2761 65038
rect -2601 64878 -2589 65038
rect -2773 64866 -2589 64878
rect -3159 64060 -2975 64072
rect -3159 63900 -3147 64060
rect -2987 63900 -2975 64060
rect -3159 63888 -2975 63900
rect -1893 64060 -1709 64072
rect -1473 64060 -1313 65319
rect -1893 63900 -1881 64060
rect -1721 63991 -1313 64060
rect -1721 63900 -1497 63991
rect -1893 63888 -1709 63900
rect -1509 63831 -1497 63900
rect -1337 63831 -1313 63991
rect -763 65026 -603 65320
rect -763 64890 -751 65026
rect -615 64890 -603 65026
rect -763 63980 -603 64890
rect -1509 63819 -1313 63831
rect -764 63820 -603 63980
rect -2773 63538 -2589 63550
rect -2773 63378 -2761 63538
rect -2601 63378 -2589 63538
rect -2773 63366 -2589 63378
rect -3159 62560 -2975 62572
rect -3159 62400 -3147 62560
rect -2987 62400 -2975 62560
rect -3159 62388 -2975 62400
rect -1893 62560 -1709 62572
rect -1473 62560 -1313 63819
rect -1893 62400 -1881 62560
rect -1721 62491 -1313 62560
rect -1721 62400 -1497 62491
rect -1893 62388 -1709 62400
rect -1509 62331 -1497 62400
rect -1337 62331 -1313 62491
rect -763 63526 -603 63820
rect -763 63390 -751 63526
rect -615 63390 -603 63526
rect -763 62480 -603 63390
rect -1509 62319 -1313 62331
rect -764 62320 -603 62480
rect -2773 62038 -2589 62050
rect -2773 61878 -2761 62038
rect -2601 61878 -2589 62038
rect -2773 61866 -2589 61878
rect -3159 61060 -2975 61072
rect -3159 60900 -3147 61060
rect -2987 60900 -2975 61060
rect -3159 60888 -2975 60900
rect -1893 61060 -1709 61072
rect -1473 61060 -1313 62319
rect -1893 60900 -1881 61060
rect -1721 60991 -1313 61060
rect -1721 60900 -1497 60991
rect -1893 60888 -1709 60900
rect -1509 60831 -1497 60900
rect -1337 60831 -1313 60991
rect -763 62026 -603 62320
rect -763 61890 -751 62026
rect -615 61890 -603 62026
rect -763 60980 -603 61890
rect -1509 60819 -1313 60831
rect -764 60820 -603 60980
rect -2773 60538 -2589 60550
rect -2773 60378 -2761 60538
rect -2601 60378 -2589 60538
rect -2773 60366 -2589 60378
rect -3159 59560 -2975 59572
rect -3159 59400 -3147 59560
rect -2987 59400 -2975 59560
rect -3159 59388 -2975 59400
rect -1893 59560 -1709 59572
rect -1473 59560 -1313 60819
rect -1893 59400 -1881 59560
rect -1721 59491 -1313 59560
rect -1721 59400 -1497 59491
rect -1893 59388 -1709 59400
rect -1509 59331 -1497 59400
rect -1337 59331 -1313 59491
rect -763 60526 -603 60820
rect -763 60390 -751 60526
rect -615 60390 -603 60526
rect -763 59480 -603 60390
rect -1509 59319 -1313 59331
rect -764 59320 -603 59480
rect -2773 59038 -2589 59050
rect -2773 58878 -2761 59038
rect -2601 58878 -2589 59038
rect -2773 58866 -2589 58878
rect -3159 58060 -2975 58072
rect -3159 57900 -3147 58060
rect -2987 57900 -2975 58060
rect -3159 57888 -2975 57900
rect -1893 58060 -1709 58072
rect -1473 58060 -1313 59319
rect -1893 57900 -1881 58060
rect -1721 57991 -1313 58060
rect -1721 57900 -1497 57991
rect -1893 57888 -1709 57900
rect -1509 57831 -1497 57900
rect -1337 57831 -1313 57991
rect -763 59026 -603 59320
rect -763 58890 -751 59026
rect -615 58890 -603 59026
rect -763 57980 -603 58890
rect -1509 57819 -1313 57831
rect -764 57820 -603 57980
rect -2773 57538 -2589 57550
rect -2773 57378 -2761 57538
rect -2601 57378 -2589 57538
rect -2773 57366 -2589 57378
rect -3159 56560 -2975 56572
rect -3159 56400 -3147 56560
rect -2987 56400 -2975 56560
rect -3159 56388 -2975 56400
rect -1893 56560 -1709 56572
rect -1473 56560 -1313 57819
rect -1893 56400 -1881 56560
rect -1721 56491 -1313 56560
rect -1721 56400 -1497 56491
rect -1893 56388 -1709 56400
rect -1509 56331 -1497 56400
rect -1337 56331 -1313 56491
rect -763 57526 -603 57820
rect -763 57390 -751 57526
rect -615 57390 -603 57526
rect -763 56480 -603 57390
rect -1509 56319 -1313 56331
rect -764 56320 -603 56480
rect -2773 56038 -2589 56050
rect -2773 55878 -2761 56038
rect -2601 55878 -2589 56038
rect -2773 55866 -2589 55878
rect -3159 55060 -2975 55072
rect -3159 54900 -3147 55060
rect -2987 54900 -2975 55060
rect -3159 54888 -2975 54900
rect -1893 55060 -1709 55072
rect -1473 55060 -1313 56319
rect -1893 54900 -1881 55060
rect -1721 54991 -1313 55060
rect -1721 54900 -1497 54991
rect -1893 54888 -1709 54900
rect -1509 54831 -1497 54900
rect -1337 54831 -1313 54991
rect -763 56026 -603 56320
rect -763 55890 -751 56026
rect -615 55890 -603 56026
rect -763 54980 -603 55890
rect -1509 54819 -1313 54831
rect -764 54820 -603 54980
rect -2773 54538 -2589 54550
rect -2773 54378 -2761 54538
rect -2601 54378 -2589 54538
rect -2773 54366 -2589 54378
rect -3159 53560 -2975 53572
rect -3159 53400 -3147 53560
rect -2987 53400 -2975 53560
rect -3159 53388 -2975 53400
rect -1893 53560 -1709 53572
rect -1473 53560 -1313 54819
rect -1893 53400 -1881 53560
rect -1721 53491 -1313 53560
rect -1721 53400 -1497 53491
rect -1893 53388 -1709 53400
rect -1509 53331 -1497 53400
rect -1337 53331 -1313 53491
rect -763 54526 -603 54820
rect -763 54390 -751 54526
rect -615 54390 -603 54526
rect -763 53480 -603 54390
rect -1509 53319 -1313 53331
rect -764 53320 -603 53480
rect -2773 53038 -2589 53050
rect -2773 52878 -2761 53038
rect -2601 52878 -2589 53038
rect -2773 52866 -2589 52878
rect -3159 52060 -2975 52072
rect -3159 51900 -3147 52060
rect -2987 51900 -2975 52060
rect -3159 51888 -2975 51900
rect -1893 52060 -1709 52072
rect -1473 52060 -1313 53319
rect -1893 51900 -1881 52060
rect -1721 51991 -1313 52060
rect -1721 51900 -1497 51991
rect -1893 51888 -1709 51900
rect -1509 51831 -1497 51900
rect -1337 51831 -1313 51991
rect -763 53026 -603 53320
rect -763 52890 -751 53026
rect -615 52890 -603 53026
rect -763 51980 -603 52890
rect -1509 51819 -1313 51831
rect -764 51820 -603 51980
rect -2773 51538 -2589 51550
rect -2773 51378 -2761 51538
rect -2601 51378 -2589 51538
rect -2773 51366 -2589 51378
rect -3159 50560 -2975 50572
rect -3159 50400 -3147 50560
rect -2987 50400 -2975 50560
rect -3159 50388 -2975 50400
rect -1893 50560 -1709 50572
rect -1473 50560 -1313 51819
rect -1893 50400 -1881 50560
rect -1721 50491 -1313 50560
rect -1721 50400 -1497 50491
rect -1893 50388 -1709 50400
rect -1509 50331 -1497 50400
rect -1337 50331 -1313 50491
rect -763 51526 -603 51820
rect -763 51390 -751 51526
rect -615 51390 -603 51526
rect -763 50480 -603 51390
rect -1509 50319 -1313 50331
rect -764 50320 -603 50480
rect -2773 50038 -2589 50050
rect -2773 49878 -2761 50038
rect -2601 49878 -2589 50038
rect -2773 49866 -2589 49878
rect -3159 49060 -2975 49072
rect -3159 48900 -3147 49060
rect -2987 48900 -2975 49060
rect -3159 48888 -2975 48900
rect -1893 49060 -1709 49072
rect -1473 49060 -1313 50319
rect -1893 48900 -1881 49060
rect -1721 48991 -1313 49060
rect -1721 48900 -1497 48991
rect -1893 48888 -1709 48900
rect -1509 48831 -1497 48900
rect -1337 48831 -1313 48991
rect -763 50026 -603 50320
rect -763 49890 -751 50026
rect -615 49890 -603 50026
rect -763 48980 -603 49890
rect -1509 48819 -1313 48831
rect -764 48820 -603 48980
rect -2773 48538 -2589 48550
rect -2773 48378 -2761 48538
rect -2601 48378 -2589 48538
rect -2773 48366 -2589 48378
rect -3159 47560 -2975 47572
rect -3159 47400 -3147 47560
rect -2987 47400 -2975 47560
rect -3159 47388 -2975 47400
rect -1893 47560 -1709 47572
rect -1473 47560 -1313 48819
rect -1893 47400 -1881 47560
rect -1721 47491 -1313 47560
rect -1721 47400 -1497 47491
rect -1893 47388 -1709 47400
rect -1509 47331 -1497 47400
rect -1337 47331 -1313 47491
rect -763 48526 -603 48820
rect -763 48390 -751 48526
rect -615 48390 -603 48526
rect -763 47480 -603 48390
rect -1509 47319 -1313 47331
rect -764 47320 -603 47480
rect -3159 46060 -2975 46072
rect -3159 45900 -3147 46060
rect -2987 45900 -2975 46060
rect -3159 45888 -2975 45900
rect -1893 46060 -1709 46072
rect -1473 46060 -1313 47319
rect -1893 45900 -1881 46060
rect -1721 45991 -1313 46060
rect -1721 45900 -1497 45991
rect -1893 45888 -1709 45900
rect -1509 45831 -1497 45900
rect -1337 45831 -1313 45991
rect -763 45980 -603 47320
rect -1509 45819 -1313 45831
rect -764 45820 -603 45980
rect -2773 45538 -2589 45550
rect -2773 45378 -2761 45538
rect -2601 45378 -2589 45538
rect -2773 45366 -2589 45378
rect -3159 44560 -2975 44572
rect -3159 44400 -3147 44560
rect -2987 44400 -2975 44560
rect -3159 44388 -2975 44400
rect -1893 44560 -1709 44572
rect -1473 44560 -1313 45819
rect -1893 44400 -1881 44560
rect -1721 44491 -1313 44560
rect -1721 44400 -1497 44491
rect -1893 44388 -1709 44400
rect -1509 44331 -1497 44400
rect -1337 44331 -1313 44491
rect -763 45526 -603 45820
rect -763 45390 -751 45526
rect -615 45390 -603 45526
rect -763 44480 -603 45390
rect -1509 44319 -1313 44331
rect -764 44320 -603 44480
rect -2773 44038 -2589 44050
rect -2773 43878 -2761 44038
rect -2601 43878 -2589 44038
rect -2773 43866 -2589 43878
rect -3159 43060 -2975 43072
rect -3159 42900 -3147 43060
rect -2987 42900 -2975 43060
rect -3159 42888 -2975 42900
rect -1893 43060 -1709 43072
rect -1473 43060 -1313 44319
rect -1893 42900 -1881 43060
rect -1721 42991 -1313 43060
rect -1721 42900 -1497 42991
rect -1893 42888 -1709 42900
rect -1509 42831 -1497 42900
rect -1337 42831 -1313 42991
rect -763 44026 -603 44320
rect -763 43890 -751 44026
rect -615 43890 -603 44026
rect -763 42980 -603 43890
rect -1509 42819 -1313 42831
rect -764 42820 -603 42980
rect -2773 42538 -2589 42550
rect -2773 42378 -2761 42538
rect -2601 42378 -2589 42538
rect -2773 42366 -2589 42378
rect -3159 41560 -2975 41572
rect -3159 41400 -3147 41560
rect -2987 41400 -2975 41560
rect -3159 41388 -2975 41400
rect -1893 41560 -1709 41572
rect -1473 41560 -1313 42819
rect -1893 41400 -1881 41560
rect -1721 41491 -1313 41560
rect -1721 41400 -1497 41491
rect -1893 41388 -1709 41400
rect -1509 41331 -1497 41400
rect -1337 41331 -1313 41491
rect -763 42526 -603 42820
rect -763 42390 -751 42526
rect -615 42390 -603 42526
rect -763 41480 -603 42390
rect -1509 41319 -1313 41331
rect -764 41320 -603 41480
rect -2773 41038 -2589 41050
rect -2773 40878 -2761 41038
rect -2601 40878 -2589 41038
rect -2773 40866 -2589 40878
rect -3159 40060 -2975 40072
rect -3159 39900 -3147 40060
rect -2987 39900 -2975 40060
rect -3159 39888 -2975 39900
rect -1893 40060 -1709 40072
rect -1473 40060 -1313 41319
rect -1893 39900 -1881 40060
rect -1721 39991 -1313 40060
rect -1721 39900 -1497 39991
rect -1893 39888 -1709 39900
rect -1509 39831 -1497 39900
rect -1337 39831 -1313 39991
rect -763 41026 -603 41320
rect -763 40890 -751 41026
rect -615 40890 -603 41026
rect -763 39980 -603 40890
rect -1509 39819 -1313 39831
rect -764 39820 -603 39980
rect -2773 39538 -2589 39550
rect -2773 39378 -2761 39538
rect -2601 39378 -2589 39538
rect -2773 39366 -2589 39378
rect -3159 38560 -2975 38572
rect -3159 38400 -3147 38560
rect -2987 38400 -2975 38560
rect -3159 38388 -2975 38400
rect -1893 38560 -1709 38572
rect -1473 38560 -1313 39819
rect -1893 38400 -1881 38560
rect -1721 38491 -1313 38560
rect -1721 38400 -1497 38491
rect -1893 38388 -1709 38400
rect -1509 38331 -1497 38400
rect -1337 38331 -1313 38491
rect -763 39526 -603 39820
rect -763 39390 -751 39526
rect -615 39390 -603 39526
rect -763 38480 -603 39390
rect -1509 38319 -1313 38331
rect -764 38320 -603 38480
rect -2773 38038 -2589 38050
rect -2773 37878 -2761 38038
rect -2601 37878 -2589 38038
rect -2773 37866 -2589 37878
rect -3159 37060 -2975 37072
rect -3159 36900 -3147 37060
rect -2987 36900 -2975 37060
rect -3159 36888 -2975 36900
rect -1893 37060 -1709 37072
rect -1473 37060 -1313 38319
rect -1893 36900 -1881 37060
rect -1721 36991 -1313 37060
rect -1721 36900 -1497 36991
rect -1893 36888 -1709 36900
rect -1509 36831 -1497 36900
rect -1337 36831 -1313 36991
rect -763 38026 -603 38320
rect -763 37890 -751 38026
rect -615 37890 -603 38026
rect -763 36980 -603 37890
rect -1509 36819 -1313 36831
rect -764 36820 -603 36980
rect -2773 36538 -2589 36550
rect -2773 36378 -2761 36538
rect -2601 36378 -2589 36538
rect -2773 36366 -2589 36378
rect -3159 35560 -2975 35572
rect -3159 35400 -3147 35560
rect -2987 35400 -2975 35560
rect -3159 35388 -2975 35400
rect -1893 35560 -1709 35572
rect -1473 35560 -1313 36819
rect -1893 35400 -1881 35560
rect -1721 35491 -1313 35560
rect -1721 35400 -1497 35491
rect -1893 35388 -1709 35400
rect -1509 35331 -1497 35400
rect -1337 35331 -1313 35491
rect -763 36526 -603 36820
rect -763 36390 -751 36526
rect -615 36390 -603 36526
rect -763 35480 -603 36390
rect -1509 35319 -1313 35331
rect -764 35320 -603 35480
rect -2773 35038 -2589 35050
rect -2773 34878 -2761 35038
rect -2601 34878 -2589 35038
rect -2773 34866 -2589 34878
rect -3159 34060 -2975 34072
rect -3159 33900 -3147 34060
rect -2987 33900 -2975 34060
rect -3159 33888 -2975 33900
rect -1893 34060 -1709 34072
rect -1473 34060 -1313 35319
rect -1893 33900 -1881 34060
rect -1721 33991 -1313 34060
rect -1721 33900 -1497 33991
rect -1893 33888 -1709 33900
rect -1509 33831 -1497 33900
rect -1337 33831 -1313 33991
rect -763 35026 -603 35320
rect -763 34890 -751 35026
rect -615 34890 -603 35026
rect -763 33980 -603 34890
rect -1509 33819 -1313 33831
rect -764 33820 -603 33980
rect -2773 33538 -2589 33550
rect -2773 33378 -2761 33538
rect -2601 33378 -2589 33538
rect -2773 33366 -2589 33378
rect -3159 32560 -2975 32572
rect -3159 32400 -3147 32560
rect -2987 32400 -2975 32560
rect -3159 32388 -2975 32400
rect -1893 32560 -1709 32572
rect -1473 32560 -1313 33819
rect -1893 32400 -1881 32560
rect -1721 32491 -1313 32560
rect -1721 32400 -1497 32491
rect -1893 32388 -1709 32400
rect -1509 32331 -1497 32400
rect -1337 32331 -1313 32491
rect -763 33526 -603 33820
rect -763 33390 -751 33526
rect -615 33390 -603 33526
rect -763 32480 -603 33390
rect -1509 32319 -1313 32331
rect -764 32320 -603 32480
rect -2773 32038 -2589 32050
rect -2773 31878 -2761 32038
rect -2601 31878 -2589 32038
rect -2773 31866 -2589 31878
rect -3159 31060 -2975 31072
rect -3159 30900 -3147 31060
rect -2987 30900 -2975 31060
rect -3159 30888 -2975 30900
rect -1893 31060 -1709 31072
rect -1473 31060 -1313 32319
rect -1893 30900 -1881 31060
rect -1721 30991 -1313 31060
rect -1721 30900 -1497 30991
rect -1893 30888 -1709 30900
rect -1509 30831 -1497 30900
rect -1337 30831 -1313 30991
rect -763 32026 -603 32320
rect -763 31890 -751 32026
rect -615 31890 -603 32026
rect -763 30980 -603 31890
rect -1509 30819 -1313 30831
rect -764 30820 -603 30980
rect -2773 30538 -2589 30550
rect -2773 30378 -2761 30538
rect -2601 30378 -2589 30538
rect -2773 30366 -2589 30378
rect -3159 29560 -2975 29572
rect -3159 29400 -3147 29560
rect -2987 29400 -2975 29560
rect -3159 29388 -2975 29400
rect -1893 29560 -1709 29572
rect -1473 29560 -1313 30819
rect -1893 29400 -1881 29560
rect -1721 29491 -1313 29560
rect -1721 29400 -1497 29491
rect -1893 29388 -1709 29400
rect -1509 29331 -1497 29400
rect -1337 29331 -1313 29491
rect -763 30526 -603 30820
rect -763 30390 -751 30526
rect -615 30390 -603 30526
rect -763 29480 -603 30390
rect -1509 29319 -1313 29331
rect -764 29320 -603 29480
rect -2773 29038 -2589 29050
rect -2773 28878 -2761 29038
rect -2601 28878 -2589 29038
rect -2773 28866 -2589 28878
rect -1473 28060 -1313 29319
rect -1560 27991 -1313 28060
rect -1560 27900 -1497 27991
rect -1509 27831 -1497 27900
rect -1337 27831 -1313 27991
rect -763 29026 -603 29320
rect -763 28890 -751 29026
rect -615 28890 -603 29026
rect -763 27980 -603 28890
rect -1509 27819 -1313 27831
rect -764 27820 -603 27980
rect -2773 27538 -2589 27550
rect -2773 27378 -2761 27538
rect -2601 27378 -2589 27538
rect -2773 27366 -2589 27378
rect -3159 26560 -2975 26572
rect -3159 26400 -3147 26560
rect -2987 26400 -2975 26560
rect -3159 26388 -2975 26400
rect -1893 26560 -1709 26572
rect -1473 26560 -1313 27819
rect -1893 26400 -1881 26560
rect -1721 26491 -1313 26560
rect -1721 26400 -1497 26491
rect -1893 26388 -1709 26400
rect -1509 26331 -1497 26400
rect -1337 26331 -1313 26491
rect -763 27526 -603 27820
rect -763 27390 -751 27526
rect -615 27390 -603 27526
rect -763 26480 -603 27390
rect -1509 26319 -1313 26331
rect -764 26320 -603 26480
rect -2773 26038 -2589 26050
rect -2773 25878 -2761 26038
rect -2601 25878 -2589 26038
rect -2773 25866 -2589 25878
rect -3159 25060 -2975 25072
rect -3159 24900 -3147 25060
rect -2987 24900 -2975 25060
rect -3159 24888 -2975 24900
rect -1893 25060 -1709 25072
rect -1473 25060 -1313 26319
rect -1893 24900 -1881 25060
rect -1721 24991 -1313 25060
rect -1721 24900 -1497 24991
rect -1893 24888 -1709 24900
rect -1509 24831 -1497 24900
rect -1337 24831 -1313 24991
rect -763 26026 -603 26320
rect -763 25890 -751 26026
rect -615 25890 -603 26026
rect -763 24980 -603 25890
rect -1509 24819 -1313 24831
rect -764 24820 -603 24980
rect -2773 24538 -2589 24550
rect -2773 24378 -2761 24538
rect -2601 24378 -2589 24538
rect -2773 24366 -2589 24378
rect -3159 23560 -2975 23572
rect -3159 23400 -3147 23560
rect -2987 23400 -2975 23560
rect -3159 23388 -2975 23400
rect -1893 23560 -1709 23572
rect -1473 23560 -1313 24819
rect -1893 23400 -1881 23560
rect -1721 23491 -1313 23560
rect -1721 23400 -1497 23491
rect -1893 23388 -1709 23400
rect -1509 23331 -1497 23400
rect -1337 23331 -1313 23491
rect -763 24526 -603 24820
rect -763 24390 -751 24526
rect -615 24390 -603 24526
rect -763 23480 -603 24390
rect -1509 23319 -1313 23331
rect -764 23320 -603 23480
rect -2773 23038 -2589 23050
rect -2773 22878 -2761 23038
rect -2601 22878 -2589 23038
rect -2773 22866 -2589 22878
rect -3159 22060 -2975 22072
rect -3159 21900 -3147 22060
rect -2987 21900 -2975 22060
rect -3159 21888 -2975 21900
rect -1893 22060 -1709 22072
rect -1473 22060 -1313 23319
rect -1893 21900 -1881 22060
rect -1721 21991 -1313 22060
rect -1721 21900 -1497 21991
rect -1893 21888 -1709 21900
rect -1509 21831 -1497 21900
rect -1337 21831 -1313 21991
rect -763 23026 -603 23320
rect -763 22890 -751 23026
rect -615 22890 -603 23026
rect -763 21980 -603 22890
rect -1509 21819 -1313 21831
rect -764 21820 -603 21980
rect -2773 21538 -2589 21550
rect -2773 21378 -2761 21538
rect -2601 21378 -2589 21538
rect -2773 21366 -2589 21378
rect -3159 20560 -2975 20572
rect -3159 20400 -3147 20560
rect -2987 20400 -2975 20560
rect -3159 20388 -2975 20400
rect -1893 20560 -1709 20572
rect -1473 20560 -1313 21819
rect -1893 20400 -1881 20560
rect -1721 20491 -1313 20560
rect -1721 20400 -1497 20491
rect -1893 20388 -1709 20400
rect -1509 20331 -1497 20400
rect -1337 20331 -1313 20491
rect -763 21526 -603 21820
rect -763 21390 -751 21526
rect -615 21390 -603 21526
rect -763 20480 -603 21390
rect -1509 20319 -1313 20331
rect -764 20320 -603 20480
rect -2773 20038 -2589 20050
rect -2773 19878 -2761 20038
rect -2601 19878 -2589 20038
rect -2773 19866 -2589 19878
rect -3159 19060 -2975 19072
rect -3159 18900 -3147 19060
rect -2987 18900 -2975 19060
rect -3159 18888 -2975 18900
rect -1893 19060 -1709 19072
rect -1473 19060 -1313 20319
rect -1893 18900 -1881 19060
rect -1721 18991 -1313 19060
rect -1721 18900 -1497 18991
rect -1893 18888 -1709 18900
rect -1509 18831 -1497 18900
rect -1337 18831 -1313 18991
rect -763 20026 -603 20320
rect -763 19890 -751 20026
rect -615 19890 -603 20026
rect -763 18980 -603 19890
rect -1509 18819 -1313 18831
rect -764 18820 -603 18980
rect -2773 18538 -2589 18550
rect -2773 18378 -2761 18538
rect -2601 18378 -2589 18538
rect -2773 18366 -2589 18378
rect -3159 17560 -2975 17572
rect -3159 17400 -3147 17560
rect -2987 17400 -2975 17560
rect -3159 17388 -2975 17400
rect -1893 17560 -1709 17572
rect -1473 17560 -1313 18819
rect -1893 17400 -1881 17560
rect -1721 17491 -1313 17560
rect -1721 17400 -1497 17491
rect -1893 17388 -1709 17400
rect -1509 17331 -1497 17400
rect -1337 17331 -1313 17491
rect -763 18526 -603 18820
rect -763 18390 -751 18526
rect -615 18390 -603 18526
rect -763 17480 -603 18390
rect -1509 17319 -1313 17331
rect -764 17320 -603 17480
rect -2773 17038 -2589 17050
rect -2773 16878 -2761 17038
rect -2601 16878 -2589 17038
rect -2773 16866 -2589 16878
rect -3159 16060 -2975 16072
rect -3159 15900 -3147 16060
rect -2987 15900 -2975 16060
rect -3159 15888 -2975 15900
rect -1893 16060 -1709 16072
rect -1473 16060 -1313 17319
rect -1893 15900 -1881 16060
rect -1721 15991 -1313 16060
rect -1721 15900 -1497 15991
rect -1893 15888 -1709 15900
rect -1509 15831 -1497 15900
rect -1337 15831 -1313 15991
rect -763 17026 -603 17320
rect -763 16890 -751 17026
rect -615 16890 -603 17026
rect -763 15980 -603 16890
rect -1509 15819 -1313 15831
rect -764 15820 -603 15980
rect -2773 15538 -2589 15550
rect -2773 15378 -2761 15538
rect -2601 15378 -2589 15538
rect -2773 15366 -2589 15378
rect -3159 14560 -2975 14572
rect -3159 14400 -3147 14560
rect -2987 14400 -2975 14560
rect -3159 14388 -2975 14400
rect -1893 14560 -1709 14572
rect -1473 14560 -1313 15819
rect -1893 14400 -1881 14560
rect -1721 14491 -1313 14560
rect -1721 14400 -1497 14491
rect -1893 14388 -1709 14400
rect -1509 14331 -1497 14400
rect -1337 14331 -1313 14491
rect -763 15526 -603 15820
rect -763 15390 -751 15526
rect -615 15390 -603 15526
rect -763 14480 -603 15390
rect -1509 14319 -1313 14331
rect -764 14320 -603 14480
rect -2773 14038 -2589 14050
rect -2773 13878 -2761 14038
rect -2601 13878 -2589 14038
rect -2773 13866 -2589 13878
rect -3159 13060 -2975 13072
rect -3159 12900 -3147 13060
rect -2987 12900 -2975 13060
rect -3159 12888 -2975 12900
rect -1893 13060 -1709 13072
rect -1473 13060 -1313 14319
rect -1893 12900 -1881 13060
rect -1721 12991 -1313 13060
rect -1721 12900 -1497 12991
rect -1893 12888 -1709 12900
rect -1509 12831 -1497 12900
rect -1337 12831 -1313 12991
rect -763 14026 -603 14320
rect -763 13890 -751 14026
rect -615 13890 -603 14026
rect -763 12980 -603 13890
rect -1509 12819 -1313 12831
rect -764 12820 -603 12980
rect -2773 12538 -2589 12550
rect -2773 12378 -2761 12538
rect -2601 12378 -2589 12538
rect -2773 12366 -2589 12378
rect -3159 11560 -2975 11572
rect -3159 11400 -3147 11560
rect -2987 11400 -2975 11560
rect -3159 11388 -2975 11400
rect -1893 11560 -1709 11572
rect -1473 11560 -1313 12819
rect -1893 11400 -1881 11560
rect -1721 11491 -1313 11560
rect -1721 11400 -1497 11491
rect -1893 11388 -1709 11400
rect -1509 11331 -1497 11400
rect -1337 11331 -1313 11491
rect -763 12526 -603 12820
rect -763 12390 -751 12526
rect -615 12390 -603 12526
rect -763 11480 -603 12390
rect -1509 11319 -1313 11331
rect -764 11320 -603 11480
rect -2773 11038 -2589 11050
rect -2773 10878 -2761 11038
rect -2601 10878 -2589 11038
rect -2773 10866 -2589 10878
rect -3159 10060 -2975 10072
rect -3159 9900 -3147 10060
rect -2987 9900 -2975 10060
rect -3159 9888 -2975 9900
rect -1893 10060 -1709 10072
rect -1473 10060 -1313 11319
rect -1893 9900 -1881 10060
rect -1721 9900 -1313 10060
rect -763 11026 -603 11320
rect -763 10890 -751 11026
rect -615 10890 -603 11026
rect -763 9980 -603 10890
rect -1893 9888 -1709 9900
rect -2773 9538 -2589 9550
rect -2773 9378 -2761 9538
rect -2601 9378 -2589 9538
rect -2773 9366 -2589 9378
rect -3207 9013 -3047 9093
rect -3219 9001 -3035 9013
rect -3219 8841 -3207 9001
rect -3047 8841 -3035 9001
rect -3219 8829 -3035 8841
rect -3207 8687 -3047 8829
rect -1473 8644 -1313 9900
rect -764 9820 -603 9980
rect -763 9526 -603 9820
rect -763 9390 -751 9526
rect -615 9390 -603 9526
rect 151963 160667 152123 162158
rect 151963 160531 151975 160667
rect 152111 160531 152123 160667
rect 151963 159167 152123 160531
rect 151963 159031 151975 159167
rect 152111 159031 152123 159167
rect 151963 157667 152123 159031
rect 151963 157531 151975 157667
rect 152111 157531 152123 157667
rect 151963 156167 152123 157531
rect 151963 156031 151975 156167
rect 152111 156031 152123 156167
rect 151963 154667 152123 156031
rect 151963 154531 151975 154667
rect 152111 154531 152123 154667
rect 151963 153167 152123 154531
rect 151963 153031 151975 153167
rect 152111 153031 152123 153167
rect 151963 151667 152123 153031
rect 151963 151531 151975 151667
rect 152111 151531 152123 151667
rect 151963 150167 152123 151531
rect 151963 150031 151975 150167
rect 152111 150031 152123 150167
rect 151963 148667 152123 150031
rect 151963 148531 151975 148667
rect 152111 148531 152123 148667
rect 151963 147167 152123 148531
rect 151963 147031 151975 147167
rect 152111 147031 152123 147167
rect 151963 145667 152123 147031
rect 151963 145531 151975 145667
rect 152111 145531 152123 145667
rect 151963 144167 152123 145531
rect 151963 144031 151975 144167
rect 152111 144031 152123 144167
rect 151963 142667 152123 144031
rect 151963 142531 151975 142667
rect 152111 142531 152123 142667
rect 151963 141167 152123 142531
rect 151963 141031 151975 141167
rect 152111 141031 152123 141167
rect 151963 139667 152123 141031
rect 151963 139531 151975 139667
rect 152111 139531 152123 139667
rect 151963 138167 152123 139531
rect 151963 138031 151975 138167
rect 152111 138031 152123 138167
rect 151963 136667 152123 138031
rect 151963 136531 151975 136667
rect 152111 136531 152123 136667
rect 151963 135167 152123 136531
rect 151963 135031 151975 135167
rect 152111 135031 152123 135167
rect 151963 133667 152123 135031
rect 151963 133531 151975 133667
rect 152111 133531 152123 133667
rect 151963 132167 152123 133531
rect 151963 132031 151975 132167
rect 152111 132031 152123 132167
rect 151963 130667 152123 132031
rect 151963 130531 151975 130667
rect 152111 130531 152123 130667
rect 151963 129167 152123 130531
rect 151963 129031 151975 129167
rect 152111 129031 152123 129167
rect 151963 127667 152123 129031
rect 151963 127531 151975 127667
rect 152111 127531 152123 127667
rect 151963 126167 152123 127531
rect 151963 126031 151975 126167
rect 152111 126031 152123 126167
rect 151963 124667 152123 126031
rect 151963 124531 151975 124667
rect 152111 124531 152123 124667
rect 151963 123167 152123 124531
rect 151963 123031 151975 123167
rect 152111 123031 152123 123167
rect 151963 121667 152123 123031
rect 151963 121531 151975 121667
rect 152111 121531 152123 121667
rect 151963 120167 152123 121531
rect 151963 120031 151975 120167
rect 152111 120031 152123 120167
rect 151963 118667 152123 120031
rect 151963 118531 151975 118667
rect 152111 118531 152123 118667
rect 151963 117167 152123 118531
rect 151963 117031 151975 117167
rect 152111 117031 152123 117167
rect 151963 115667 152123 117031
rect 151963 115531 151975 115667
rect 152111 115531 152123 115667
rect 151963 114167 152123 115531
rect 151963 114031 151975 114167
rect 152111 114031 152123 114167
rect 151963 112667 152123 114031
rect 151963 112531 151975 112667
rect 152111 112531 152123 112667
rect 151963 111167 152123 112531
rect 151963 111031 151975 111167
rect 152111 111031 152123 111167
rect 151963 109667 152123 111031
rect 151963 109531 151975 109667
rect 152111 109531 152123 109667
rect 151963 108167 152123 109531
rect 151963 108031 151975 108167
rect 152111 108031 152123 108167
rect 151963 106667 152123 108031
rect 151963 106531 151975 106667
rect 152111 106531 152123 106667
rect 151963 105167 152123 106531
rect 151963 105031 151975 105167
rect 152111 105031 152123 105167
rect 151963 103667 152123 105031
rect 151963 103531 151975 103667
rect 152111 103531 152123 103667
rect 151963 102167 152123 103531
rect 151963 102031 151975 102167
rect 152111 102031 152123 102167
rect 151963 100667 152123 102031
rect 151963 100531 151975 100667
rect 152111 100531 152123 100667
rect 151963 99167 152123 100531
rect 151963 99031 151975 99167
rect 152111 99031 152123 99167
rect 151963 97667 152123 99031
rect 151963 97531 151975 97667
rect 152111 97531 152123 97667
rect 151963 96167 152123 97531
rect 151963 96031 151975 96167
rect 152111 96031 152123 96167
rect 151963 94667 152123 96031
rect 151963 94531 151975 94667
rect 152111 94531 152123 94667
rect 151963 93167 152123 94531
rect 151963 93031 151975 93167
rect 152111 93031 152123 93167
rect 151963 91667 152123 93031
rect 151963 91531 151975 91667
rect 152111 91531 152123 91667
rect 151963 90167 152123 91531
rect 151963 90031 151975 90167
rect 152111 90031 152123 90167
rect 151963 88667 152123 90031
rect 151963 88531 151975 88667
rect 152111 88531 152123 88667
rect 151963 87167 152123 88531
rect 151963 87031 151975 87167
rect 152111 87031 152123 87167
rect 151963 85667 152123 87031
rect 151963 85531 151975 85667
rect 152111 85531 152123 85667
rect 151963 84167 152123 85531
rect 151963 84031 151975 84167
rect 152111 84031 152123 84167
rect 151963 82667 152123 84031
rect 151963 82531 151975 82667
rect 152111 82531 152123 82667
rect 151963 81167 152123 82531
rect 151963 81031 151975 81167
rect 152111 81031 152123 81167
rect 151963 79667 152123 81031
rect 151963 79531 151975 79667
rect 152111 79531 152123 79667
rect 151963 78167 152123 79531
rect 151963 78031 151975 78167
rect 152111 78031 152123 78167
rect 151963 76667 152123 78031
rect 151963 76531 151975 76667
rect 152111 76531 152123 76667
rect 151963 75167 152123 76531
rect 151963 75031 151975 75167
rect 152111 75031 152123 75167
rect 151963 73667 152123 75031
rect 151963 73531 151975 73667
rect 152111 73531 152123 73667
rect 151963 72167 152123 73531
rect 151963 72031 151975 72167
rect 152111 72031 152123 72167
rect 151963 70667 152123 72031
rect 151963 70531 151975 70667
rect 152111 70531 152123 70667
rect 151963 69167 152123 70531
rect 151963 69031 151975 69167
rect 152111 69031 152123 69167
rect 151963 67667 152123 69031
rect 151963 67531 151975 67667
rect 152111 67531 152123 67667
rect 151963 66167 152123 67531
rect 151963 66031 151975 66167
rect 152111 66031 152123 66167
rect 151963 64667 152123 66031
rect 151963 64531 151975 64667
rect 152111 64531 152123 64667
rect 151963 63167 152123 64531
rect 151963 63031 151975 63167
rect 152111 63031 152123 63167
rect 151963 61667 152123 63031
rect 151963 61531 151975 61667
rect 152111 61531 152123 61667
rect 151963 60167 152123 61531
rect 151963 60031 151975 60167
rect 152111 60031 152123 60167
rect 151963 58667 152123 60031
rect 151963 58531 151975 58667
rect 152111 58531 152123 58667
rect 151963 57167 152123 58531
rect 151963 57031 151975 57167
rect 152111 57031 152123 57167
rect 151963 55667 152123 57031
rect 151963 55531 151975 55667
rect 152111 55531 152123 55667
rect 151963 54167 152123 55531
rect 151963 54031 151975 54167
rect 152111 54031 152123 54167
rect 151963 52667 152123 54031
rect 151963 52531 151975 52667
rect 152111 52531 152123 52667
rect 151963 51167 152123 52531
rect 151963 51031 151975 51167
rect 152111 51031 152123 51167
rect 151963 49667 152123 51031
rect 151963 49531 151975 49667
rect 152111 49531 152123 49667
rect 151963 48167 152123 49531
rect 151963 48031 151975 48167
rect 152111 48031 152123 48167
rect 151963 46667 152123 48031
rect 151963 46531 151975 46667
rect 152111 46531 152123 46667
rect 151963 45167 152123 46531
rect 151963 45031 151975 45167
rect 152111 45031 152123 45167
rect 151963 43667 152123 45031
rect 151963 43531 151975 43667
rect 152111 43531 152123 43667
rect 151963 42167 152123 43531
rect 151963 42031 151975 42167
rect 152111 42031 152123 42167
rect 151963 40667 152123 42031
rect 151963 40531 151975 40667
rect 152111 40531 152123 40667
rect 151963 39167 152123 40531
rect 151963 39031 151975 39167
rect 152111 39031 152123 39167
rect 151963 37667 152123 39031
rect 151963 37531 151975 37667
rect 152111 37531 152123 37667
rect 151963 36167 152123 37531
rect 151963 36031 151975 36167
rect 152111 36031 152123 36167
rect 151963 34667 152123 36031
rect 151963 34531 151975 34667
rect 152111 34531 152123 34667
rect 151963 33167 152123 34531
rect 151963 33031 151975 33167
rect 152111 33031 152123 33167
rect 151963 31667 152123 33031
rect 151963 31531 151975 31667
rect 152111 31531 152123 31667
rect 151963 30167 152123 31531
rect 151963 30031 151975 30167
rect 152111 30031 152123 30167
rect 151963 28667 152123 30031
rect 151963 28531 151975 28667
rect 152111 28531 152123 28667
rect 151963 27167 152123 28531
rect 151963 27031 151975 27167
rect 152111 27031 152123 27167
rect 151963 25667 152123 27031
rect 151963 25531 151975 25667
rect 152111 25531 152123 25667
rect 151963 24167 152123 25531
rect 151963 24031 151975 24167
rect 152111 24031 152123 24167
rect 151963 22667 152123 24031
rect 151963 22531 151975 22667
rect 152111 22531 152123 22667
rect 151963 21167 152123 22531
rect 151963 21031 151975 21167
rect 152111 21031 152123 21167
rect 151963 19667 152123 21031
rect 151963 19531 151975 19667
rect 152111 19531 152123 19667
rect 151963 18167 152123 19531
rect 151963 18031 151975 18167
rect 152111 18031 152123 18167
rect 151963 16667 152123 18031
rect 151963 16531 151975 16667
rect 152111 16531 152123 16667
rect 151963 15167 152123 16531
rect 151963 15031 151975 15167
rect 152111 15031 152123 15167
rect 151963 13667 152123 15031
rect 151963 13531 151975 13667
rect 152111 13531 152123 13667
rect 151963 12167 152123 13531
rect 151963 12031 151975 12167
rect 152111 12031 152123 12167
rect 151963 10667 152123 12031
rect 151963 10531 151975 10667
rect 152111 10531 152123 10667
rect -763 9380 -603 9390
rect 144786 9380 144976 9395
rect 151963 9380 152123 10531
rect -789 9368 152131 9380
rect -789 9232 1844 9368
rect 1980 9232 9056 9368
rect 9192 9232 16469 9368
rect 16605 9232 32140 9368
rect 32276 9232 60851 9368
rect 60987 9232 83786 9368
rect 83922 9232 90286 9368
rect 90422 9232 94786 9368
rect 94922 9232 99286 9368
rect 99422 9232 102286 9368
rect 102422 9232 105786 9368
rect 105922 9232 111786 9368
rect 111922 9232 116286 9368
rect 116422 9232 119286 9368
rect 119422 9232 125286 9368
rect 125422 9232 131986 9368
rect 132122 9232 134986 9368
rect 135122 9232 136486 9368
rect 136622 9232 137986 9368
rect 138122 9232 140986 9368
rect 141122 9232 142986 9368
rect 143122 9232 146986 9368
rect 147122 9232 148486 9368
rect 148622 9232 149986 9368
rect 150122 9232 151486 9368
rect 151622 9232 152131 9368
rect -789 9220 152131 9232
rect 144786 9211 144976 9220
rect 151963 9052 152123 9220
rect 152718 8644 152878 163111
rect -1491 8632 152878 8644
rect -1491 8496 151945 8632
rect 152081 8496 152878 8632
rect -1491 8484 152878 8496
rect -1473 8452 -1313 8484
rect 322 8437 482 8484
rect 1822 8437 1982 8484
rect 3322 8437 3482 8484
rect 4822 8437 4982 8484
rect 6322 8437 6482 8484
rect 7822 8437 7982 8484
rect 9322 8437 9482 8484
rect 10822 8437 10982 8484
rect 12322 8437 12482 8484
rect 13822 8437 13982 8484
rect 15322 8437 15482 8484
rect 16822 8437 16982 8484
rect 18322 8437 18482 8484
rect 19822 8437 19982 8484
rect 21322 8437 21482 8484
rect 22822 8437 22982 8484
rect 24322 8437 24482 8484
rect 25822 8437 25982 8484
rect 27322 8437 27482 8484
rect 28822 8437 28982 8484
rect 30322 8437 30482 8484
rect 31822 8437 31982 8484
rect 33322 8437 33482 8484
rect 34822 8437 34982 8484
rect 36322 8437 36482 8484
rect 37822 8437 37982 8484
rect 39322 8437 39482 8484
rect 40822 8437 40982 8484
rect 42322 8437 42482 8484
rect 43822 8437 43982 8484
rect 45322 8437 45482 8484
rect 46822 8437 46982 8484
rect 48322 8437 48482 8484
rect 49822 8437 49982 8484
rect 51322 8437 51482 8484
rect 52822 8437 52982 8484
rect 54322 8437 54482 8484
rect 55822 8437 55982 8484
rect 57322 8437 57482 8484
rect 58822 8437 58982 8484
rect 60322 8437 60482 8484
rect 61822 8437 61982 8484
rect 63322 8437 63482 8484
rect 64822 8437 64982 8484
rect 66322 8437 66482 8484
rect 67822 8437 67982 8484
rect 69322 8437 69482 8484
rect 70822 8437 70982 8484
rect 72322 8437 72482 8484
rect 73822 8437 73982 8484
rect 75322 8437 75482 8484
rect 76822 8437 76982 8484
rect 78322 8437 78482 8484
rect 79822 8437 79982 8484
rect 81322 8437 81482 8484
rect 82822 8437 82982 8484
rect 84322 8437 84482 8484
rect 85822 8437 85982 8484
rect 87322 8437 87482 8484
rect 88822 8437 88982 8484
rect 90322 8437 90482 8484
rect 91822 8437 91982 8484
rect 93322 8437 93482 8484
rect 94822 8437 94982 8484
rect 96322 8437 96482 8484
rect 97822 8437 97982 8484
rect 99322 8437 99482 8484
rect 100822 8437 100982 8484
rect 102322 8437 102482 8484
rect 103822 8437 103982 8484
rect 105322 8437 105482 8484
rect 106822 8437 106982 8484
rect 108322 8437 108482 8484
rect 109822 8437 109982 8484
rect 111322 8437 111482 8484
rect 112822 8437 112982 8484
rect 114322 8437 114482 8484
rect 115822 8437 115982 8484
rect 117322 8437 117482 8484
rect 118822 8437 118982 8484
rect 120322 8437 120482 8484
rect 121822 8437 121982 8484
rect 123322 8437 123482 8484
rect 124822 8437 124982 8484
rect 126322 8437 126482 8484
rect 127822 8437 127982 8484
rect 129322 8437 129482 8484
rect 130822 8437 130982 8484
rect 132322 8437 132482 8484
rect 135322 8437 135482 8484
rect 136822 8437 136982 8484
rect 138322 8437 138482 8484
rect 139822 8437 139982 8484
rect 141322 8437 141482 8484
rect 142822 8437 142982 8484
rect 144322 8437 144482 8484
rect 145822 8437 145982 8484
rect 147322 8437 147482 8484
rect 148822 8437 148982 8484
rect 150322 8437 150482 8484
rect 151458 8205 151649 8217
rect 151458 8044 151470 8205
rect 151637 8044 151649 8205
rect 151458 8032 151649 8044
rect 153437 8024 153597 8421
rect 1817 7844 2007 7856
rect 12 7821 196 7833
rect 12 7661 24 7821
rect 184 7661 418 7821
rect 1817 7684 1829 7844
rect 1995 7684 2007 7844
rect 1817 7672 2007 7684
rect 9029 7853 9219 7865
rect 9029 7693 9041 7853
rect 9207 7693 9219 7853
rect 9029 7681 9219 7693
rect 16442 7841 16632 7853
rect 16442 7681 16454 7841
rect 16620 7681 16632 7841
rect 16442 7669 16632 7681
rect 32113 7845 32303 7857
rect 32113 7685 32125 7845
rect 32291 7685 32303 7845
rect 32113 7673 32303 7685
rect 60824 7852 61014 7864
rect 60824 7692 60836 7852
rect 61002 7692 61014 7852
rect 60824 7680 61014 7692
rect 83759 7853 83949 7865
rect 83759 7693 83771 7853
rect 83937 7693 83949 7853
rect 83759 7681 83949 7693
rect 90259 7853 90449 7865
rect 90259 7693 90271 7853
rect 90437 7693 90449 7853
rect 90259 7681 90449 7693
rect 94759 7853 94949 7865
rect 94759 7693 94771 7853
rect 94937 7693 94949 7853
rect 94759 7681 94949 7693
rect 99259 7853 99449 7865
rect 99259 7693 99271 7853
rect 99437 7693 99449 7853
rect 99259 7681 99449 7693
rect 102259 7853 102449 7865
rect 102259 7693 102271 7853
rect 102437 7693 102449 7853
rect 102259 7681 102449 7693
rect 105759 7853 105949 7865
rect 105759 7693 105771 7853
rect 105937 7693 105949 7853
rect 105759 7681 105949 7693
rect 111759 7853 111949 7865
rect 111759 7693 111771 7853
rect 111937 7693 111949 7853
rect 111759 7681 111949 7693
rect 116259 7853 116449 7865
rect 116259 7693 116271 7853
rect 116437 7693 116449 7853
rect 116259 7681 116449 7693
rect 119259 7853 119449 7865
rect 119259 7693 119271 7853
rect 119437 7693 119449 7853
rect 119259 7681 119449 7693
rect 125259 7853 125449 7865
rect 125259 7693 125271 7853
rect 125437 7693 125449 7853
rect 125259 7681 125449 7693
rect 131959 7853 132149 7865
rect 131959 7693 131971 7853
rect 132137 7693 132149 7853
rect 131959 7681 132149 7693
rect 134959 7853 135149 7865
rect 134959 7693 134971 7853
rect 135137 7693 135149 7853
rect 134959 7681 135149 7693
rect 136459 7853 136649 7865
rect 136459 7693 136471 7853
rect 136637 7693 136649 7853
rect 136459 7681 136649 7693
rect 137959 7853 138149 7865
rect 137959 7693 137971 7853
rect 138137 7693 138149 7853
rect 137959 7681 138149 7693
rect 140959 7853 141149 7865
rect 140959 7693 140971 7853
rect 141137 7693 141149 7853
rect 140959 7681 141149 7693
rect 142959 7853 143149 7865
rect 142959 7693 142971 7853
rect 143137 7693 143149 7853
rect 142959 7681 143149 7693
rect 146959 7853 147149 7865
rect 146959 7693 146971 7853
rect 147137 7693 147149 7853
rect 146959 7681 147149 7693
rect 148459 7853 148649 7865
rect 148459 7693 148471 7853
rect 148637 7693 148649 7853
rect 148459 7681 148649 7693
rect 149959 7853 150149 7865
rect 149959 7693 149971 7853
rect 150137 7693 150149 7853
rect 149959 7681 150149 7693
rect 151459 7853 151649 7865
rect 151459 7693 151471 7853
rect 151637 7693 151649 7853
rect 151459 7681 151649 7693
rect 151921 7846 152105 7858
rect 151921 7686 151933 7846
rect 152093 7686 152105 7846
rect 151921 7674 152105 7686
rect 12 7649 196 7661
use pixel_array100x100  pixel_array100x100_0
timestamp 1655251759
transform 1 0 1054 0 1 158689
box -1500 -149300 150370 2875
use shift_register  shift_register_0
timestamp 1757709129
transform 0 1 -10536 -1 0 161992
box -538 -2 153994 8000
use shift_registerC  shift_registerC_0
timestamp 1757709129
transform 1 0 29 0 1 295
box -538 -2 153994 8000
<< labels >>
rlabel metal5 -1421 9375 -1417 9380 1 VDD
<< end >>
