magic
tech sky130A
magscale 1 2
timestamp 1758069660
<< error_p >>
rect -855 71 -797 77
rect -737 71 -679 77
rect -619 71 -561 77
rect -501 71 -443 77
rect -383 71 -325 77
rect -265 71 -207 77
rect -147 71 -89 77
rect -29 71 29 77
rect 89 71 147 77
rect 207 71 265 77
rect 325 71 383 77
rect 443 71 501 77
rect 561 71 619 77
rect 679 71 737 77
rect 797 71 855 77
rect -855 37 -843 71
rect -737 37 -725 71
rect -619 37 -607 71
rect -501 37 -489 71
rect -383 37 -371 71
rect -265 37 -253 71
rect -147 37 -135 71
rect -29 37 -17 71
rect 89 37 101 71
rect 207 37 219 71
rect 325 37 337 71
rect 443 37 455 71
rect 561 37 573 71
rect 679 37 691 71
rect 797 37 809 71
rect -855 31 -797 37
rect -737 31 -679 37
rect -619 31 -561 37
rect -501 31 -443 37
rect -383 31 -325 37
rect -265 31 -207 37
rect -147 31 -89 37
rect -29 31 29 37
rect 89 31 147 37
rect 207 31 265 37
rect 325 31 383 37
rect 443 31 501 37
rect 561 31 619 37
rect 679 31 737 37
rect 797 31 855 37
rect -855 -37 -797 -31
rect -737 -37 -679 -31
rect -619 -37 -561 -31
rect -501 -37 -443 -31
rect -383 -37 -325 -31
rect -265 -37 -207 -31
rect -147 -37 -89 -31
rect -29 -37 29 -31
rect 89 -37 147 -31
rect 207 -37 265 -31
rect 325 -37 383 -31
rect 443 -37 501 -31
rect 561 -37 619 -31
rect 679 -37 737 -31
rect 797 -37 855 -31
rect -855 -71 -843 -37
rect -737 -71 -725 -37
rect -619 -71 -607 -37
rect -501 -71 -489 -37
rect -383 -71 -371 -37
rect -265 -71 -253 -37
rect -147 -71 -135 -37
rect -29 -71 -17 -37
rect 89 -71 101 -37
rect 207 -71 219 -37
rect 325 -71 337 -37
rect 443 -71 455 -37
rect 561 -71 573 -37
rect 679 -71 691 -37
rect 797 -71 809 -37
rect -855 -77 -797 -71
rect -737 -77 -679 -71
rect -619 -77 -561 -71
rect -501 -77 -443 -71
rect -383 -77 -325 -71
rect -265 -77 -207 -71
rect -147 -77 -89 -71
rect -29 -77 29 -71
rect 89 -77 147 -71
rect 207 -77 265 -71
rect 325 -77 383 -71
rect 443 -77 501 -71
rect 561 -77 619 -71
rect 679 -77 737 -71
rect 797 -77 855 -71
<< pwell >>
rect -1052 -919 1052 919
<< nmos >>
rect -856 109 -796 709
rect -738 109 -678 709
rect -620 109 -560 709
rect -502 109 -442 709
rect -384 109 -324 709
rect -266 109 -206 709
rect -148 109 -88 709
rect -30 109 30 709
rect 88 109 148 709
rect 206 109 266 709
rect 324 109 384 709
rect 442 109 502 709
rect 560 109 620 709
rect 678 109 738 709
rect 796 109 856 709
rect -856 -709 -796 -109
rect -738 -709 -678 -109
rect -620 -709 -560 -109
rect -502 -709 -442 -109
rect -384 -709 -324 -109
rect -266 -709 -206 -109
rect -148 -709 -88 -109
rect -30 -709 30 -109
rect 88 -709 148 -109
rect 206 -709 266 -109
rect 324 -709 384 -109
rect 442 -709 502 -109
rect 560 -709 620 -109
rect 678 -709 738 -109
rect 796 -709 856 -109
<< ndiff >>
rect -914 697 -856 709
rect -914 121 -902 697
rect -868 121 -856 697
rect -914 109 -856 121
rect -796 697 -738 709
rect -796 121 -784 697
rect -750 121 -738 697
rect -796 109 -738 121
rect -678 697 -620 709
rect -678 121 -666 697
rect -632 121 -620 697
rect -678 109 -620 121
rect -560 697 -502 709
rect -560 121 -548 697
rect -514 121 -502 697
rect -560 109 -502 121
rect -442 697 -384 709
rect -442 121 -430 697
rect -396 121 -384 697
rect -442 109 -384 121
rect -324 697 -266 709
rect -324 121 -312 697
rect -278 121 -266 697
rect -324 109 -266 121
rect -206 697 -148 709
rect -206 121 -194 697
rect -160 121 -148 697
rect -206 109 -148 121
rect -88 697 -30 709
rect -88 121 -76 697
rect -42 121 -30 697
rect -88 109 -30 121
rect 30 697 88 709
rect 30 121 42 697
rect 76 121 88 697
rect 30 109 88 121
rect 148 697 206 709
rect 148 121 160 697
rect 194 121 206 697
rect 148 109 206 121
rect 266 697 324 709
rect 266 121 278 697
rect 312 121 324 697
rect 266 109 324 121
rect 384 697 442 709
rect 384 121 396 697
rect 430 121 442 697
rect 384 109 442 121
rect 502 697 560 709
rect 502 121 514 697
rect 548 121 560 697
rect 502 109 560 121
rect 620 697 678 709
rect 620 121 632 697
rect 666 121 678 697
rect 620 109 678 121
rect 738 697 796 709
rect 738 121 750 697
rect 784 121 796 697
rect 738 109 796 121
rect 856 697 914 709
rect 856 121 868 697
rect 902 121 914 697
rect 856 109 914 121
rect -914 -121 -856 -109
rect -914 -697 -902 -121
rect -868 -697 -856 -121
rect -914 -709 -856 -697
rect -796 -121 -738 -109
rect -796 -697 -784 -121
rect -750 -697 -738 -121
rect -796 -709 -738 -697
rect -678 -121 -620 -109
rect -678 -697 -666 -121
rect -632 -697 -620 -121
rect -678 -709 -620 -697
rect -560 -121 -502 -109
rect -560 -697 -548 -121
rect -514 -697 -502 -121
rect -560 -709 -502 -697
rect -442 -121 -384 -109
rect -442 -697 -430 -121
rect -396 -697 -384 -121
rect -442 -709 -384 -697
rect -324 -121 -266 -109
rect -324 -697 -312 -121
rect -278 -697 -266 -121
rect -324 -709 -266 -697
rect -206 -121 -148 -109
rect -206 -697 -194 -121
rect -160 -697 -148 -121
rect -206 -709 -148 -697
rect -88 -121 -30 -109
rect -88 -697 -76 -121
rect -42 -697 -30 -121
rect -88 -709 -30 -697
rect 30 -121 88 -109
rect 30 -697 42 -121
rect 76 -697 88 -121
rect 30 -709 88 -697
rect 148 -121 206 -109
rect 148 -697 160 -121
rect 194 -697 206 -121
rect 148 -709 206 -697
rect 266 -121 324 -109
rect 266 -697 278 -121
rect 312 -697 324 -121
rect 266 -709 324 -697
rect 384 -121 442 -109
rect 384 -697 396 -121
rect 430 -697 442 -121
rect 384 -709 442 -697
rect 502 -121 560 -109
rect 502 -697 514 -121
rect 548 -697 560 -121
rect 502 -709 560 -697
rect 620 -121 678 -109
rect 620 -697 632 -121
rect 666 -697 678 -121
rect 620 -709 678 -697
rect 738 -121 796 -109
rect 738 -697 750 -121
rect 784 -697 796 -121
rect 738 -709 796 -697
rect 856 -121 914 -109
rect 856 -697 868 -121
rect 902 -697 914 -121
rect 856 -709 914 -697
<< ndiffc >>
rect -902 121 -868 697
rect -784 121 -750 697
rect -666 121 -632 697
rect -548 121 -514 697
rect -430 121 -396 697
rect -312 121 -278 697
rect -194 121 -160 697
rect -76 121 -42 697
rect 42 121 76 697
rect 160 121 194 697
rect 278 121 312 697
rect 396 121 430 697
rect 514 121 548 697
rect 632 121 666 697
rect 750 121 784 697
rect 868 121 902 697
rect -902 -697 -868 -121
rect -784 -697 -750 -121
rect -666 -697 -632 -121
rect -548 -697 -514 -121
rect -430 -697 -396 -121
rect -312 -697 -278 -121
rect -194 -697 -160 -121
rect -76 -697 -42 -121
rect 42 -697 76 -121
rect 160 -697 194 -121
rect 278 -697 312 -121
rect 396 -697 430 -121
rect 514 -697 548 -121
rect 632 -697 666 -121
rect 750 -697 784 -121
rect 868 -697 902 -121
<< psubdiff >>
rect -1016 849 -920 883
rect 920 849 1016 883
rect -1016 787 -982 849
rect 982 787 1016 849
rect -1016 -849 -982 -787
rect 982 -849 1016 -787
rect -1016 -883 -920 -849
rect 920 -883 1016 -849
<< psubdiffcont >>
rect -920 849 920 883
rect -1016 -787 -982 787
rect 982 -787 1016 787
rect -920 -883 920 -849
<< poly >>
rect -859 731 -793 797
rect -741 731 -675 797
rect -623 731 -557 797
rect -505 731 -439 797
rect -387 731 -321 797
rect -269 731 -203 797
rect -151 731 -85 797
rect -33 731 33 797
rect 85 731 151 797
rect 203 731 269 797
rect 321 731 387 797
rect 439 731 505 797
rect 557 731 623 797
rect 675 731 741 797
rect 793 731 859 797
rect -856 709 -796 731
rect -738 709 -678 731
rect -620 709 -560 731
rect -502 709 -442 731
rect -384 709 -324 731
rect -266 709 -206 731
rect -148 709 -88 731
rect -30 709 30 731
rect 88 709 148 731
rect 206 709 266 731
rect 324 709 384 731
rect 442 709 502 731
rect 560 709 620 731
rect 678 709 738 731
rect 796 709 856 731
rect -856 87 -796 109
rect -738 87 -678 109
rect -620 87 -560 109
rect -502 87 -442 109
rect -384 87 -324 109
rect -266 87 -206 109
rect -148 87 -88 109
rect -30 87 30 109
rect 88 87 148 109
rect 206 87 266 109
rect 324 87 384 109
rect 442 87 502 109
rect 560 87 620 109
rect 678 87 738 109
rect 796 87 856 109
rect -859 71 -793 87
rect -859 37 -843 71
rect -809 37 -793 71
rect -859 21 -793 37
rect -741 71 -675 87
rect -741 37 -725 71
rect -691 37 -675 71
rect -741 21 -675 37
rect -623 71 -557 87
rect -623 37 -607 71
rect -573 37 -557 71
rect -623 21 -557 37
rect -505 71 -439 87
rect -505 37 -489 71
rect -455 37 -439 71
rect -505 21 -439 37
rect -387 71 -321 87
rect -387 37 -371 71
rect -337 37 -321 71
rect -387 21 -321 37
rect -269 71 -203 87
rect -269 37 -253 71
rect -219 37 -203 71
rect -269 21 -203 37
rect -151 71 -85 87
rect -151 37 -135 71
rect -101 37 -85 71
rect -151 21 -85 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 85 71 151 87
rect 85 37 101 71
rect 135 37 151 71
rect 85 21 151 37
rect 203 71 269 87
rect 203 37 219 71
rect 253 37 269 71
rect 203 21 269 37
rect 321 71 387 87
rect 321 37 337 71
rect 371 37 387 71
rect 321 21 387 37
rect 439 71 505 87
rect 439 37 455 71
rect 489 37 505 71
rect 439 21 505 37
rect 557 71 623 87
rect 557 37 573 71
rect 607 37 623 71
rect 557 21 623 37
rect 675 71 741 87
rect 675 37 691 71
rect 725 37 741 71
rect 675 21 741 37
rect 793 71 859 87
rect 793 37 809 71
rect 843 37 859 71
rect 793 21 859 37
rect -859 -37 -793 -21
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -859 -87 -793 -71
rect -741 -37 -675 -21
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -741 -87 -675 -71
rect -623 -37 -557 -21
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -623 -87 -557 -71
rect -505 -37 -439 -21
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -505 -87 -439 -71
rect -387 -37 -321 -21
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -387 -87 -321 -71
rect -269 -37 -203 -21
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -269 -87 -203 -71
rect -151 -37 -85 -21
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -151 -87 -85 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 85 -37 151 -21
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 85 -87 151 -71
rect 203 -37 269 -21
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 203 -87 269 -71
rect 321 -37 387 -21
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 321 -87 387 -71
rect 439 -37 505 -21
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 439 -87 505 -71
rect 557 -37 623 -21
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 557 -87 623 -71
rect 675 -37 741 -21
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 675 -87 741 -71
rect 793 -37 859 -21
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 793 -87 859 -71
rect -856 -109 -796 -87
rect -738 -109 -678 -87
rect -620 -109 -560 -87
rect -502 -109 -442 -87
rect -384 -109 -324 -87
rect -266 -109 -206 -87
rect -148 -109 -88 -87
rect -30 -109 30 -87
rect 88 -109 148 -87
rect 206 -109 266 -87
rect 324 -109 384 -87
rect 442 -109 502 -87
rect 560 -109 620 -87
rect 678 -109 738 -87
rect 796 -109 856 -87
rect -856 -731 -796 -709
rect -738 -731 -678 -709
rect -620 -731 -560 -709
rect -502 -731 -442 -709
rect -384 -731 -324 -709
rect -266 -731 -206 -709
rect -148 -731 -88 -709
rect -30 -731 30 -709
rect 88 -731 148 -709
rect 206 -731 266 -709
rect 324 -731 384 -709
rect 442 -731 502 -709
rect 560 -731 620 -709
rect 678 -731 738 -709
rect 796 -731 856 -709
rect -859 -797 -793 -731
rect -741 -797 -675 -731
rect -623 -797 -557 -731
rect -505 -797 -439 -731
rect -387 -797 -321 -731
rect -269 -797 -203 -731
rect -151 -797 -85 -731
rect -33 -797 33 -731
rect 85 -797 151 -731
rect 203 -797 269 -731
rect 321 -797 387 -731
rect 439 -797 505 -731
rect 557 -797 623 -731
rect 675 -797 741 -731
rect 793 -797 859 -731
<< polycont >>
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
<< locali >>
rect -1016 849 -920 883
rect 920 849 1016 883
rect -1016 787 -982 849
rect 982 787 1016 849
rect -902 697 -868 713
rect -902 105 -868 121
rect -784 697 -750 713
rect -784 105 -750 121
rect -666 697 -632 713
rect -666 105 -632 121
rect -548 697 -514 713
rect -548 105 -514 121
rect -430 697 -396 713
rect -430 105 -396 121
rect -312 697 -278 713
rect -312 105 -278 121
rect -194 697 -160 713
rect -194 105 -160 121
rect -76 697 -42 713
rect -76 105 -42 121
rect 42 697 76 713
rect 42 105 76 121
rect 160 697 194 713
rect 160 105 194 121
rect 278 697 312 713
rect 278 105 312 121
rect 396 697 430 713
rect 396 105 430 121
rect 514 697 548 713
rect 514 105 548 121
rect 632 697 666 713
rect 632 105 666 121
rect 750 697 784 713
rect 750 105 784 121
rect 868 697 902 713
rect 868 105 902 121
rect -859 37 -843 71
rect -809 37 -793 71
rect -741 37 -725 71
rect -691 37 -675 71
rect -623 37 -607 71
rect -573 37 -557 71
rect -505 37 -489 71
rect -455 37 -439 71
rect -387 37 -371 71
rect -337 37 -321 71
rect -269 37 -253 71
rect -219 37 -203 71
rect -151 37 -135 71
rect -101 37 -85 71
rect -33 37 -17 71
rect 17 37 33 71
rect 85 37 101 71
rect 135 37 151 71
rect 203 37 219 71
rect 253 37 269 71
rect 321 37 337 71
rect 371 37 387 71
rect 439 37 455 71
rect 489 37 505 71
rect 557 37 573 71
rect 607 37 623 71
rect 675 37 691 71
rect 725 37 741 71
rect 793 37 809 71
rect 843 37 859 71
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 793 -71 809 -37
rect 843 -71 859 -37
rect -902 -121 -868 -105
rect -902 -713 -868 -697
rect -784 -121 -750 -105
rect -784 -713 -750 -697
rect -666 -121 -632 -105
rect -666 -713 -632 -697
rect -548 -121 -514 -105
rect -548 -713 -514 -697
rect -430 -121 -396 -105
rect -430 -713 -396 -697
rect -312 -121 -278 -105
rect -312 -713 -278 -697
rect -194 -121 -160 -105
rect -194 -713 -160 -697
rect -76 -121 -42 -105
rect -76 -713 -42 -697
rect 42 -121 76 -105
rect 42 -713 76 -697
rect 160 -121 194 -105
rect 160 -713 194 -697
rect 278 -121 312 -105
rect 278 -713 312 -697
rect 396 -121 430 -105
rect 396 -713 430 -697
rect 514 -121 548 -105
rect 514 -713 548 -697
rect 632 -121 666 -105
rect 632 -713 666 -697
rect 750 -121 784 -105
rect 750 -713 784 -697
rect 868 -121 902 -105
rect 868 -713 902 -697
rect -1016 -849 -982 -787
rect 982 -849 1016 -787
rect -1016 -883 -920 -849
rect 920 -883 1016 -849
<< viali >>
rect -902 121 -868 697
rect -784 121 -750 697
rect -666 121 -632 697
rect -548 121 -514 697
rect -430 121 -396 697
rect -312 121 -278 697
rect -194 121 -160 697
rect -76 121 -42 697
rect 42 121 76 697
rect 160 121 194 697
rect 278 121 312 697
rect 396 121 430 697
rect 514 121 548 697
rect 632 121 666 697
rect 750 121 784 697
rect 868 121 902 697
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect -902 -697 -868 -121
rect -784 -697 -750 -121
rect -666 -697 -632 -121
rect -548 -697 -514 -121
rect -430 -697 -396 -121
rect -312 -697 -278 -121
rect -194 -697 -160 -121
rect -76 -697 -42 -121
rect 42 -697 76 -121
rect 160 -697 194 -121
rect 278 -697 312 -121
rect 396 -697 430 -121
rect 514 -697 548 -121
rect 632 -697 666 -121
rect 750 -697 784 -121
rect 868 -697 902 -121
<< metal1 >>
rect -908 697 -862 709
rect -908 121 -902 697
rect -868 121 -862 697
rect -908 109 -862 121
rect -790 697 -744 709
rect -790 121 -784 697
rect -750 121 -744 697
rect -790 109 -744 121
rect -672 697 -626 709
rect -672 121 -666 697
rect -632 121 -626 697
rect -672 109 -626 121
rect -554 697 -508 709
rect -554 121 -548 697
rect -514 121 -508 697
rect -554 109 -508 121
rect -436 697 -390 709
rect -436 121 -430 697
rect -396 121 -390 697
rect -436 109 -390 121
rect -318 697 -272 709
rect -318 121 -312 697
rect -278 121 -272 697
rect -318 109 -272 121
rect -200 697 -154 709
rect -200 121 -194 697
rect -160 121 -154 697
rect -200 109 -154 121
rect -82 697 -36 709
rect -82 121 -76 697
rect -42 121 -36 697
rect -82 109 -36 121
rect 36 697 82 709
rect 36 121 42 697
rect 76 121 82 697
rect 36 109 82 121
rect 154 697 200 709
rect 154 121 160 697
rect 194 121 200 697
rect 154 109 200 121
rect 272 697 318 709
rect 272 121 278 697
rect 312 121 318 697
rect 272 109 318 121
rect 390 697 436 709
rect 390 121 396 697
rect 430 121 436 697
rect 390 109 436 121
rect 508 697 554 709
rect 508 121 514 697
rect 548 121 554 697
rect 508 109 554 121
rect 626 697 672 709
rect 626 121 632 697
rect 666 121 672 697
rect 626 109 672 121
rect 744 697 790 709
rect 744 121 750 697
rect 784 121 790 697
rect 744 109 790 121
rect 862 697 908 709
rect 862 121 868 697
rect 902 121 908 697
rect 862 109 908 121
rect -855 71 -797 77
rect -855 37 -843 71
rect -809 37 -797 71
rect -855 31 -797 37
rect -737 71 -679 77
rect -737 37 -725 71
rect -691 37 -679 71
rect -737 31 -679 37
rect -619 71 -561 77
rect -619 37 -607 71
rect -573 37 -561 71
rect -619 31 -561 37
rect -501 71 -443 77
rect -501 37 -489 71
rect -455 37 -443 71
rect -501 31 -443 37
rect -383 71 -325 77
rect -383 37 -371 71
rect -337 37 -325 71
rect -383 31 -325 37
rect -265 71 -207 77
rect -265 37 -253 71
rect -219 37 -207 71
rect -265 31 -207 37
rect -147 71 -89 77
rect -147 37 -135 71
rect -101 37 -89 71
rect -147 31 -89 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 89 71 147 77
rect 89 37 101 71
rect 135 37 147 71
rect 89 31 147 37
rect 207 71 265 77
rect 207 37 219 71
rect 253 37 265 71
rect 207 31 265 37
rect 325 71 383 77
rect 325 37 337 71
rect 371 37 383 71
rect 325 31 383 37
rect 443 71 501 77
rect 443 37 455 71
rect 489 37 501 71
rect 443 31 501 37
rect 561 71 619 77
rect 561 37 573 71
rect 607 37 619 71
rect 561 31 619 37
rect 679 71 737 77
rect 679 37 691 71
rect 725 37 737 71
rect 679 31 737 37
rect 797 71 855 77
rect 797 37 809 71
rect 843 37 855 71
rect 797 31 855 37
rect -855 -37 -797 -31
rect -855 -71 -843 -37
rect -809 -71 -797 -37
rect -855 -77 -797 -71
rect -737 -37 -679 -31
rect -737 -71 -725 -37
rect -691 -71 -679 -37
rect -737 -77 -679 -71
rect -619 -37 -561 -31
rect -619 -71 -607 -37
rect -573 -71 -561 -37
rect -619 -77 -561 -71
rect -501 -37 -443 -31
rect -501 -71 -489 -37
rect -455 -71 -443 -37
rect -501 -77 -443 -71
rect -383 -37 -325 -31
rect -383 -71 -371 -37
rect -337 -71 -325 -37
rect -383 -77 -325 -71
rect -265 -37 -207 -31
rect -265 -71 -253 -37
rect -219 -71 -207 -37
rect -265 -77 -207 -71
rect -147 -37 -89 -31
rect -147 -71 -135 -37
rect -101 -71 -89 -37
rect -147 -77 -89 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 89 -37 147 -31
rect 89 -71 101 -37
rect 135 -71 147 -37
rect 89 -77 147 -71
rect 207 -37 265 -31
rect 207 -71 219 -37
rect 253 -71 265 -37
rect 207 -77 265 -71
rect 325 -37 383 -31
rect 325 -71 337 -37
rect 371 -71 383 -37
rect 325 -77 383 -71
rect 443 -37 501 -31
rect 443 -71 455 -37
rect 489 -71 501 -37
rect 443 -77 501 -71
rect 561 -37 619 -31
rect 561 -71 573 -37
rect 607 -71 619 -37
rect 561 -77 619 -71
rect 679 -37 737 -31
rect 679 -71 691 -37
rect 725 -71 737 -37
rect 679 -77 737 -71
rect 797 -37 855 -31
rect 797 -71 809 -37
rect 843 -71 855 -37
rect 797 -77 855 -71
rect -908 -121 -862 -109
rect -908 -697 -902 -121
rect -868 -697 -862 -121
rect -908 -709 -862 -697
rect -790 -121 -744 -109
rect -790 -697 -784 -121
rect -750 -697 -744 -121
rect -790 -709 -744 -697
rect -672 -121 -626 -109
rect -672 -697 -666 -121
rect -632 -697 -626 -121
rect -672 -709 -626 -697
rect -554 -121 -508 -109
rect -554 -697 -548 -121
rect -514 -697 -508 -121
rect -554 -709 -508 -697
rect -436 -121 -390 -109
rect -436 -697 -430 -121
rect -396 -697 -390 -121
rect -436 -709 -390 -697
rect -318 -121 -272 -109
rect -318 -697 -312 -121
rect -278 -697 -272 -121
rect -318 -709 -272 -697
rect -200 -121 -154 -109
rect -200 -697 -194 -121
rect -160 -697 -154 -121
rect -200 -709 -154 -697
rect -82 -121 -36 -109
rect -82 -697 -76 -121
rect -42 -697 -36 -121
rect -82 -709 -36 -697
rect 36 -121 82 -109
rect 36 -697 42 -121
rect 76 -697 82 -121
rect 36 -709 82 -697
rect 154 -121 200 -109
rect 154 -697 160 -121
rect 194 -697 200 -121
rect 154 -709 200 -697
rect 272 -121 318 -109
rect 272 -697 278 -121
rect 312 -697 318 -121
rect 272 -709 318 -697
rect 390 -121 436 -109
rect 390 -697 396 -121
rect 430 -697 436 -121
rect 390 -709 436 -697
rect 508 -121 554 -109
rect 508 -697 514 -121
rect 548 -697 554 -121
rect 508 -709 554 -697
rect 626 -121 672 -109
rect 626 -697 632 -121
rect 666 -697 672 -121
rect 626 -709 672 -697
rect 744 -121 790 -109
rect 744 -697 750 -121
rect 784 -697 790 -121
rect 744 -709 790 -697
rect 862 -121 908 -109
rect 862 -697 868 -121
rect 902 -697 908 -121
rect 862 -709 908 -697
<< properties >>
string FIXED_BBOX -999 -866 999 866
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 0.3 m 2 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
