magic
tech sky130A
timestamp 1758143371
<< metal5 >>
rect 59500 56600 60000 56800
rect 58800 56400 60000 56600
rect 58300 56300 60000 56400
rect 57800 56100 60000 56300
rect 57300 55900 60000 56100
rect 56700 55800 59800 55900
rect 56200 55600 59300 55800
rect 55500 55400 58800 55600
rect 54800 55300 58300 55400
rect 54300 55100 57800 55300
rect 53700 54900 57200 55100
rect 53000 54800 56700 54900
rect 52300 54600 56000 54800
rect 51700 54400 55500 54600
rect 0 54300 500 54400
rect 51000 54300 54800 54400
rect 0 54100 1200 54300
rect 50300 54100 54300 54300
rect 0 53900 1800 54100
rect 49500 53900 53700 54100
rect 0 53800 2500 53900
rect 48800 53800 53000 53900
rect 500 53600 3200 53800
rect 48000 53600 52300 53800
rect 1000 53400 3800 53600
rect 47200 53400 51700 53600
rect 1700 53300 4700 53400
rect 46500 53300 51000 53400
rect 2200 53100 5500 53300
rect 45700 53100 50200 53300
rect 2800 52900 6300 53100
rect 36700 52900 37000 53100
rect 44700 52900 49500 53100
rect 3500 52800 7300 52900
rect 36000 52800 37700 52900
rect 43800 52800 48700 52900
rect 4200 52600 8300 52800
rect 35700 52600 38000 52800
rect 42800 52600 48000 52800
rect 5000 52400 9500 52600
rect 35500 52400 38200 52600
rect 41800 52400 47200 52600
rect 5700 52300 10700 52400
rect 35200 52300 38300 52400
rect 40800 52300 46300 52400
rect 6700 52100 12000 52300
rect 34800 52100 38500 52300
rect 39500 52100 45500 52300
rect 7500 51900 13500 52100
rect 26700 51900 28300 52100
rect 34700 51900 44500 52100
rect 8500 51800 15200 51900
rect 26300 51800 28700 51900
rect 34500 51800 43700 51900
rect 9700 51600 17200 51800
rect 26000 51600 29200 51800
rect 34500 51600 42700 51800
rect 10700 51400 19700 51600
rect 25800 51400 29500 51600
rect 32700 51400 41500 51600
rect 12000 51300 23500 51400
rect 25700 51300 40500 51400
rect 13300 51100 39200 51300
rect 15000 50900 38300 51100
rect 16700 50800 38200 50900
rect 19000 50600 37700 50800
rect 22000 50400 31300 50600
rect 33800 50400 36800 50600
rect 25300 50300 30300 50400
rect 25500 50100 30300 50300
rect 25700 49900 30300 50100
rect 33800 50300 36500 50400
rect 33800 49900 36300 50300
rect 26000 49800 30500 49900
rect 27500 49600 30500 49800
rect 27700 49400 30500 49600
rect 27800 48800 30500 49400
rect 33700 49800 36300 49900
rect 33700 48900 36200 49800
rect 27800 47600 30700 48800
rect 27700 47100 30700 47600
rect 27500 46400 30700 47100
rect 27300 45800 30700 46400
rect 27200 45300 30700 45800
rect 27000 44800 30700 45300
rect 26800 44100 30700 44800
rect 26700 43800 30700 44100
rect 33700 48100 36300 48900
rect 33700 47600 36500 48100
rect 33700 46900 36700 47600
rect 33700 46300 36800 46900
rect 33700 45800 37000 46300
rect 33700 45300 37200 45800
rect 33700 44600 37300 45300
rect 33700 43900 37500 44600
rect 26700 43400 30500 43800
rect 26500 42400 30500 43400
rect 33700 42900 37700 43900
rect 33700 42600 37800 42900
rect 26300 40800 30500 42400
rect 33800 41400 37800 42600
rect 26300 38100 30300 40800
rect 33800 40300 38000 41400
rect 34000 38800 38000 40300
rect 33800 38600 38000 38800
rect 26300 37100 30500 38100
rect 33800 37800 37800 38600
rect 33700 37600 37800 37800
rect 33200 37400 37800 37600
rect 32700 37300 37800 37400
rect 32500 37100 37800 37300
rect 17800 36900 19200 37100
rect 16700 36800 19800 36900
rect 16200 36600 20300 36800
rect 15500 36400 20700 36600
rect 26300 36400 30700 37100
rect 32200 36900 37800 37100
rect 32000 36800 37800 36900
rect 31800 36600 37800 36800
rect 31700 36400 37800 36600
rect 15200 36300 21000 36400
rect 26500 36300 30700 36400
rect 14800 36100 21200 36300
rect 14500 35900 21300 36100
rect 14200 35800 21700 35900
rect 26500 35800 30800 36300
rect 31500 36100 37800 36400
rect 31300 35900 37800 36100
rect 13800 35600 21800 35800
rect 13700 35400 22000 35600
rect 26500 35400 31000 35800
rect 31300 35600 37700 35900
rect 31200 35400 37700 35600
rect 13500 35300 22200 35400
rect 26500 35300 37700 35400
rect 13300 35100 17200 35300
rect 19300 35100 22300 35300
rect 13200 34900 16300 35100
rect 19800 34900 22500 35100
rect 26700 34900 37700 35300
rect 13000 34800 15800 34900
rect 20200 34800 22700 34900
rect 12800 34600 15500 34800
rect 20500 34600 22800 34800
rect 12800 34400 15200 34600
rect 20700 34400 23000 34600
rect 26700 34400 37500 34900
rect 12700 34300 15000 34400
rect 20800 34300 23200 34400
rect 12500 34100 14800 34300
rect 21000 34100 23300 34300
rect 12500 33900 14500 34100
rect 21200 33900 23300 34100
rect 26800 33900 37700 34400
rect 12300 33800 14300 33900
rect 21300 33800 23500 33900
rect 12300 33600 14200 33800
rect 21500 33600 23700 33800
rect 27000 33600 37800 33900
rect 12200 33400 14000 33600
rect 21700 33400 23800 33600
rect 27000 33400 38000 33600
rect 12200 33300 13800 33400
rect 21800 33300 23800 33400
rect 27200 33300 38200 33400
rect 12200 33100 13700 33300
rect 21800 33100 24000 33300
rect 12000 32900 13700 33100
rect 22000 32900 24000 33100
rect 27300 33100 38300 33300
rect 27300 32900 38500 33100
rect 12000 32800 13500 32900
rect 22000 32800 24200 32900
rect 27500 32800 38500 32900
rect 12000 32600 13300 32800
rect 11800 32400 13300 32600
rect 22200 32600 24200 32800
rect 27700 32600 38700 32800
rect 11800 32300 13200 32400
rect 22200 32300 24300 32600
rect 27800 32400 38700 32600
rect 28000 32300 38700 32400
rect 11800 31800 13000 32300
rect 22300 31800 24500 32300
rect 28000 31900 38500 32300
rect 28000 31800 38300 31900
rect 11800 31300 12800 31800
rect 11800 30900 12700 31300
rect 22500 30900 24700 31800
rect 27800 31600 38300 31800
rect 27800 31400 38200 31600
rect 27800 31300 38000 31400
rect 27800 31100 35800 31300
rect 36200 31100 37700 31300
rect 12000 30600 12500 30900
rect 22700 28900 24700 30900
rect 27700 30900 35800 31100
rect 27700 30600 36000 30900
rect 27700 30100 36200 30600
rect 27500 29400 36300 30100
rect 27300 29100 36300 29400
rect 22500 28300 24500 28900
rect 27300 28600 36500 29100
rect 27200 28400 36500 28600
rect 22500 28100 24300 28300
rect 22300 27600 24300 28100
rect 27200 27900 36700 28400
rect 22200 27100 24200 27600
rect 27000 27100 36700 27900
rect 22200 26900 24000 27100
rect 22000 26600 24000 26900
rect 26800 26800 36700 27100
rect 22000 26100 23800 26600
rect 26800 26300 36500 26800
rect 22000 25800 23700 26100
rect 21800 25300 23700 25800
rect 26800 25900 36300 26300
rect 26800 25600 36200 25900
rect 21800 24300 23500 25300
rect 26700 25100 36000 25600
rect 26700 24800 35800 25100
rect 26700 24600 35700 24800
rect 26800 24400 35700 24600
rect 22000 23800 23500 24300
rect 26700 24300 35500 24400
rect 26700 24100 35300 24300
rect 26700 23900 35200 24100
rect 22000 23300 23700 23800
rect 22200 23100 23700 23300
rect 26700 23600 35000 23900
rect 26700 23400 34800 23600
rect 26700 23100 34700 23400
rect 22200 22800 23800 23100
rect 26500 22800 34500 23100
rect 22300 22600 24000 22800
rect 22300 22300 24200 22600
rect 26500 22400 34300 22800
rect 22500 22100 24300 22300
rect 22500 21900 24500 22100
rect 22700 21800 24800 21900
rect 26300 21800 34200 22400
rect 22800 21600 25000 21800
rect 26200 21600 34200 21800
rect 22800 21400 25300 21600
rect 26200 21400 34500 21600
rect 23000 21300 25700 21400
rect 26200 21300 34700 21400
rect 23200 21100 35000 21300
rect 23300 20900 35200 21100
rect 23700 20800 35500 20900
rect 23800 20600 35800 20800
rect 24000 20400 36200 20600
rect 24300 20300 36300 20400
rect 24500 20100 36700 20300
rect 24700 19900 37000 20100
rect 25000 19800 37200 19900
rect 25200 19600 37500 19800
rect 25000 19400 37800 19600
rect 25000 19300 38200 19400
rect 24800 19100 38300 19300
rect 24800 18900 38700 19100
rect 24700 18800 39000 18900
rect 24700 18600 39200 18800
rect 24500 18400 39500 18600
rect 24500 18300 39700 18400
rect 24300 18100 40000 18300
rect 24300 17900 40200 18100
rect 24200 17800 40300 17900
rect 24200 17600 40500 17800
rect 24000 17300 29300 17600
rect 29500 17400 40700 17600
rect 30000 17300 40800 17400
rect 23800 17100 29200 17300
rect 30500 17100 41000 17300
rect 23700 16900 29000 17100
rect 31000 16900 41000 17100
rect 23500 16800 29000 16900
rect 31800 16800 41200 16900
rect 23300 16600 28800 16800
rect 32700 16600 41200 16800
rect 23000 16400 28800 16600
rect 33700 16400 41300 16600
rect 19800 16300 28700 16400
rect 34700 16300 41300 16400
rect 18000 16100 28500 16300
rect 35500 16100 41300 16300
rect 17200 15900 28500 16100
rect 36200 15900 41500 16100
rect 16700 15800 28300 15900
rect 36700 15800 41500 15900
rect 16300 15600 28300 15800
rect 37200 15600 41500 15800
rect 16200 15400 28200 15600
rect 37500 15400 41500 15600
rect 16000 15100 28000 15400
rect 37700 15300 41500 15400
rect 37700 15100 41700 15300
rect 16000 14900 27800 15100
rect 15800 14800 27700 14900
rect 15800 14400 27500 14800
rect 15800 14300 27300 14400
rect 37800 14300 41700 15100
rect 15800 14100 27200 14300
rect 15800 13900 27000 14100
rect 38000 13900 41700 14300
rect 15800 13800 26800 13900
rect 15800 13600 26700 13800
rect 15800 13400 26300 13600
rect 15800 13300 26000 13400
rect 38000 13300 41800 13900
rect 15800 13100 25800 13300
rect 16000 12900 25500 13100
rect 16000 12800 24700 12900
rect 16000 12100 19000 12800
rect 20000 12600 23700 12800
rect 20800 12400 21800 12600
rect 38200 12400 41800 13300
rect 16200 11600 19000 12100
rect 16200 11400 19200 11600
rect 38300 11400 41800 12400
rect 16300 11300 19200 11400
rect 16300 10900 19300 11300
rect 16500 10800 19500 10900
rect 16500 10600 19700 10800
rect 38500 10600 41800 11400
rect 44700 11300 46700 11400
rect 43800 11100 46800 11300
rect 43200 10900 47000 11100
rect 42500 10800 47000 10900
rect 42200 10600 46800 10800
rect 16700 10400 19800 10600
rect 38500 10400 46800 10600
rect 16700 10300 20000 10400
rect 38500 10300 46700 10400
rect 16800 10100 20200 10300
rect 38700 10100 46500 10300
rect 16800 9900 20500 10100
rect 38700 9900 46300 10100
rect 17200 9800 20700 9900
rect 38700 9800 46000 9900
rect 17300 9600 20800 9800
rect 38700 9600 45700 9800
rect 17800 9400 21000 9600
rect 38700 9400 45200 9600
rect 18500 9300 21200 9400
rect 38800 9300 44800 9400
rect 19000 9100 21300 9300
rect 38800 9100 44300 9300
rect 19200 8900 21500 9100
rect 38800 8900 43800 9100
rect 19500 8800 21700 8900
rect 38800 8800 43300 8900
rect 19700 8600 21700 8800
rect 39000 8600 42800 8800
rect 20200 8400 21800 8600
rect 39000 8400 42300 8600
rect 20700 8300 21800 8400
rect 39200 8300 41800 8400
rect 21200 8100 21800 8300
rect 39300 8100 41300 8300
rect 39700 7900 40700 8100
<< end >>
