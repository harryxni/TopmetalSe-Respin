magic
tech sky130A
magscale 1 2
timestamp 1758069660
<< pwell >>
rect -211 -285 211 285
<< nmos >>
rect -15 -75 15 75
<< ndiff >>
rect -73 63 -15 75
rect -73 -63 -61 63
rect -27 -63 -15 63
rect -73 -75 -15 -63
rect 15 63 73 75
rect 15 -63 27 63
rect 61 -63 73 63
rect 15 -75 73 -63
<< ndiffc >>
rect -61 -63 -27 63
rect 27 -63 61 63
<< psubdiff >>
rect -175 215 -79 249
rect 79 215 175 249
rect -175 153 -141 215
rect 141 153 175 215
rect -175 -215 -141 -153
rect 141 -215 175 -153
rect -175 -249 -79 -215
rect 79 -249 175 -215
<< psubdiffcont >>
rect -79 215 79 249
rect -175 -153 -141 153
rect 141 -153 175 153
rect -79 -249 79 -215
<< poly >>
rect -69 151 69 167
rect -69 117 -53 151
rect -19 117 19 151
rect 53 117 69 151
rect -69 97 69 117
rect -15 75 15 97
rect -15 -97 15 -75
rect -33 -163 33 -97
<< polycont >>
rect -53 117 -19 151
rect 19 117 53 151
<< locali >>
rect -175 215 -79 249
rect 79 215 175 249
rect -175 153 -141 215
rect 141 153 175 215
rect -69 117 -53 151
rect -19 117 19 151
rect 53 117 69 151
rect -61 63 -27 79
rect -61 -79 -27 -63
rect 27 63 61 79
rect 27 -79 61 -63
rect -175 -215 -141 -153
rect 141 -215 175 -153
rect -175 -249 -79 -215
rect 79 -249 175 -215
<< viali >>
rect -53 117 -19 151
rect 19 117 53 151
rect -61 -63 -27 63
rect 27 -63 61 63
<< metal1 >>
rect -81 117 -71 169
rect -19 117 19 169
rect 71 117 81 169
rect -81 111 81 117
rect -67 63 -21 75
rect -67 -63 -61 63
rect -27 -63 -21 63
rect -67 -75 -21 -63
rect 21 63 67 75
rect 21 -63 27 63
rect 61 -63 67 63
rect 21 -75 67 -63
<< via1 >>
rect -71 151 -19 169
rect -71 117 -53 151
rect -53 117 -19 151
rect 19 151 71 169
rect 19 117 53 151
rect 53 117 71 151
<< metal2 >>
rect -71 169 71 179
rect -19 117 19 169
rect -71 107 71 117
<< properties >>
string FIXED_BBOX -158 -232 158 232
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w .75 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
