magic
tech sky130A
timestamp 1758153220
<< nwell >>
rect 505 -566 965 -255
<< pmoslvt >>
rect 640 -480 740 -380
<< nmoslvt >>
rect 1180 -705 1280 -585
rect 1435 -705 1535 -585
rect 1615 -665 2415 -465
rect 2615 -665 3415 -465
<< ndiff >>
rect 1615 -405 2415 -395
rect 1615 -455 1625 -405
rect 2405 -455 2415 -405
rect 1615 -465 2415 -455
rect 2615 -405 3415 -395
rect 2615 -455 2625 -405
rect 3405 -455 3415 -405
rect 2615 -465 3415 -455
rect 1180 -555 1280 -550
rect 1180 -575 1190 -555
rect 1270 -575 1280 -555
rect 1180 -585 1280 -575
rect 1435 -555 1535 -550
rect 1435 -575 1445 -555
rect 1525 -575 1535 -555
rect 1435 -585 1535 -575
rect 1615 -675 2415 -665
rect 1180 -715 1280 -705
rect 1180 -735 1190 -715
rect 1270 -735 1280 -715
rect 1180 -740 1280 -735
rect 1435 -715 1535 -705
rect 1435 -735 1445 -715
rect 1525 -735 1535 -715
rect 1615 -725 1625 -675
rect 2405 -725 2415 -675
rect 1615 -730 2415 -725
rect 2615 -675 3415 -665
rect 2615 -725 2625 -675
rect 3405 -725 3415 -675
rect 2615 -730 3415 -725
rect 1435 -740 1535 -735
<< pdiff >>
rect 595 -390 640 -380
rect 595 -470 600 -390
rect 630 -470 640 -390
rect 595 -480 640 -470
rect 740 -390 795 -380
rect 740 -470 750 -390
rect 780 -470 795 -390
rect 740 -480 795 -470
<< ndiffc >>
rect 1625 -455 2405 -405
rect 2625 -455 3405 -405
rect 1190 -575 1270 -555
rect 1445 -575 1525 -555
rect 1190 -735 1270 -715
rect 1445 -735 1525 -715
rect 1625 -725 2405 -675
rect 2625 -725 3405 -675
<< pdiffc >>
rect 600 -470 630 -390
rect 750 -470 780 -390
<< psubdiff >>
rect 2615 -745 3415 -730
rect 2615 -790 2630 -745
rect 3400 -790 3415 -745
rect 2615 -800 3415 -790
<< nsubdiff >>
rect 545 -395 595 -380
rect 545 -465 555 -395
rect 580 -465 595 -395
rect 545 -480 595 -465
<< psubdiffcont >>
rect 2630 -790 3400 -745
<< nsubdiffcont >>
rect 555 -465 580 -395
<< poly >>
rect 640 -380 740 -365
rect 640 -495 740 -480
rect 640 -525 680 -495
rect 640 -555 645 -525
rect 675 -555 680 -525
rect 640 -565 680 -555
rect 1165 -665 1180 -585
rect 1115 -670 1180 -665
rect 1115 -700 1125 -670
rect 1155 -700 1180 -670
rect 1115 -705 1180 -700
rect 1280 -705 1295 -585
rect 1420 -665 1435 -585
rect 1370 -670 1435 -665
rect 1370 -700 1380 -670
rect 1410 -700 1435 -670
rect 1370 -705 1435 -700
rect 1535 -705 1550 -585
rect 1600 -665 1615 -465
rect 2415 -590 2430 -465
rect 2415 -600 2510 -590
rect 2415 -655 2445 -600
rect 2500 -655 2510 -600
rect 2415 -665 2510 -655
rect 2600 -665 2615 -465
rect 3415 -590 3430 -465
rect 3415 -600 3510 -590
rect 3415 -655 3445 -600
rect 3500 -655 3510 -600
rect 3415 -665 3510 -655
<< polycont >>
rect 645 -555 675 -525
rect 1125 -700 1155 -670
rect 1380 -700 1410 -670
rect 2445 -655 2500 -600
rect 3445 -655 3500 -600
<< locali >>
rect 545 -305 595 -300
rect 545 -385 595 -370
rect 545 -390 640 -385
rect 545 -395 600 -390
rect 545 -465 555 -395
rect 580 -465 600 -395
rect 545 -470 600 -465
rect 630 -470 640 -390
rect 545 -475 640 -470
rect 740 -390 790 -385
rect 740 -470 750 -390
rect 780 -470 790 -390
rect 1615 -405 2575 -395
rect 1615 -455 1625 -405
rect 2405 -455 2575 -405
rect 2615 -405 3575 -395
rect 2615 -455 2625 -405
rect 3405 -455 3575 -405
rect 740 -475 790 -470
rect 750 -520 790 -475
rect 545 -525 790 -520
rect 545 -560 555 -525
rect 600 -555 645 -525
rect 675 -555 735 -525
rect 600 -560 735 -555
rect 545 -565 790 -560
rect 1125 -575 1190 -545
rect 1270 -575 1280 -545
rect 1380 -575 1445 -545
rect 1525 -575 1535 -545
rect 1125 -665 1155 -575
rect 1380 -665 1410 -575
rect 2520 -600 2575 -455
rect 3520 -600 3575 -455
rect 2430 -655 2445 -600
rect 2500 -605 2575 -600
rect 2560 -650 2575 -605
rect 2500 -655 2575 -650
rect 3430 -655 3445 -600
rect 3500 -605 3575 -600
rect 3560 -650 3575 -605
rect 3500 -655 3575 -650
rect 1090 -670 1155 -665
rect 1110 -700 1125 -670
rect 1090 -705 1155 -700
rect 1300 -670 1410 -665
rect 1300 -700 1310 -670
rect 1365 -700 1380 -670
rect 1300 -705 1410 -700
rect 1615 -675 2410 -665
rect 1125 -710 1155 -705
rect 1180 -715 1280 -705
rect 1380 -710 1410 -705
rect 1180 -735 1190 -715
rect 1270 -735 1280 -715
rect 1180 -775 1280 -735
rect 1180 -840 1185 -775
rect 1275 -840 1280 -775
rect 1180 -845 1280 -840
rect 1435 -715 1535 -705
rect 1435 -735 1445 -715
rect 1525 -735 1535 -715
rect 1435 -775 1535 -735
rect 1435 -840 1440 -775
rect 1530 -840 1535 -775
rect 1435 -845 1535 -840
rect 1615 -725 1625 -675
rect 2405 -725 2410 -675
rect 1615 -730 2410 -725
rect 2615 -675 3410 -665
rect 2615 -725 2625 -675
rect 3405 -725 3410 -675
rect 1615 -775 2415 -730
rect 1615 -960 1625 -775
rect 2405 -960 2415 -775
rect 1615 -970 2415 -960
rect 2615 -738 3410 -725
rect 2615 -745 3415 -738
rect 2615 -770 2630 -745
rect 3400 -770 3415 -745
rect 2615 -965 2625 -770
rect 3405 -965 3415 -770
rect 2615 -975 3415 -965
<< viali >>
rect 545 -370 595 -305
rect 1625 -450 2405 -405
rect 2625 -450 3405 -405
rect 555 -560 600 -525
rect 735 -560 790 -525
rect 1190 -555 1270 -545
rect 1190 -565 1270 -555
rect 1445 -555 1525 -545
rect 1445 -570 1525 -555
rect 2445 -650 2500 -605
rect 2500 -650 2560 -605
rect 3445 -650 3500 -605
rect 3500 -650 3560 -605
rect 1055 -700 1110 -670
rect 1310 -700 1365 -670
rect 1185 -840 1275 -775
rect 1440 -840 1530 -775
rect 1625 -960 2405 -775
rect 2625 -790 2630 -770
rect 2630 -790 3400 -770
rect 3400 -790 3405 -770
rect 2625 -965 3405 -790
<< metal1 >>
rect 430 -305 965 -110
rect 430 -370 545 -305
rect 595 -370 965 -305
rect 430 -375 965 -370
rect 1180 -340 1280 -337
rect 410 -525 610 -520
rect 410 -560 420 -525
rect 600 -560 610 -525
rect 410 -565 610 -560
rect 725 -525 965 -520
rect 725 -560 730 -525
rect 955 -560 965 -525
rect 725 -565 965 -560
rect 1180 -545 1280 -440
rect 1180 -565 1190 -545
rect 1270 -565 1280 -545
rect 1180 -575 1280 -565
rect 1435 -340 1535 -337
rect 1435 -545 1535 -440
rect 1615 -400 2415 -395
rect 1615 -450 1625 -400
rect 2405 -450 2415 -400
rect 1615 -455 2415 -450
rect 2615 -400 3415 -395
rect 2615 -450 2625 -400
rect 3405 -450 3415 -400
rect 2615 -455 3415 -450
rect 1435 -570 1445 -545
rect 1525 -570 1535 -545
rect 1435 -575 1535 -570
rect 2430 -605 2575 -600
rect 2430 -650 2445 -605
rect 2565 -650 2575 -605
rect 2430 -655 2575 -650
rect 3430 -605 3575 -600
rect 3430 -650 3445 -605
rect 3565 -650 3575 -605
rect 3430 -655 3575 -650
rect 1045 -670 1155 -665
rect 1045 -700 1050 -670
rect 1140 -700 1155 -670
rect 1045 -705 1155 -700
rect 1300 -670 1410 -665
rect 1300 -700 1305 -670
rect 1395 -700 1410 -670
rect 1300 -705 1410 -700
rect 765 -770 3590 -765
rect 765 -775 2625 -770
rect 765 -840 1185 -775
rect 1275 -840 1440 -775
rect 1530 -840 1625 -775
rect 765 -960 1625 -840
rect 2405 -960 2625 -775
rect 765 -965 2625 -960
rect 3405 -965 3590 -770
rect 765 -1085 3590 -965
<< via1 >>
rect 1180 -440 1280 -340
rect 420 -560 555 -525
rect 555 -560 600 -525
rect 730 -560 735 -525
rect 735 -560 790 -525
rect 790 -560 955 -525
rect 1435 -440 1535 -340
rect 1625 -405 2405 -400
rect 1625 -450 2405 -405
rect 2625 -405 3405 -400
rect 2625 -450 3405 -405
rect 2445 -650 2560 -605
rect 2560 -650 2565 -605
rect 3445 -650 3560 -605
rect 3560 -650 3565 -605
rect 1050 -700 1055 -670
rect 1055 -700 1110 -670
rect 1110 -700 1140 -670
rect 1305 -700 1310 -670
rect 1310 -700 1365 -670
rect 1365 -700 1395 -670
<< metal2 >>
rect 1175 -340 1285 -335
rect 1175 -440 1180 -340
rect 1280 -440 1285 -340
rect 1175 -445 1285 -440
rect 1430 -340 1540 -335
rect 1430 -440 1435 -340
rect 1535 -440 1540 -340
rect 1430 -445 1540 -440
rect 1615 -400 2415 -395
rect 1615 -450 1625 -400
rect 2405 -450 2415 -400
rect 1615 -455 2415 -450
rect 2615 -400 3415 -395
rect 2615 -450 2625 -400
rect 3405 -450 3415 -400
rect 2615 -455 3415 -450
rect 395 -525 610 -520
rect 395 -560 420 -525
rect 600 -560 610 -525
rect 395 -565 610 -560
rect 725 -525 965 -520
rect 725 -560 730 -525
rect 955 -560 965 -525
rect 725 -565 965 -560
rect 2430 -605 2575 -600
rect 2430 -650 2445 -605
rect 2565 -650 2575 -605
rect 2430 -655 2575 -650
rect 3430 -605 3575 -600
rect 3430 -650 3445 -605
rect 3565 -650 3575 -605
rect 3430 -655 3575 -650
rect 1045 -670 1155 -665
rect 1045 -700 1050 -670
rect 1140 -700 1155 -670
rect 1045 -705 1155 -700
rect 1300 -670 1410 -665
rect 1300 -700 1305 -670
rect 1395 -700 1410 -670
rect 1300 -705 1410 -700
rect 1045 -1117 1090 -705
rect 1300 -1112 1345 -705
rect 2520 -1102 2575 -655
rect 3520 -1102 3575 -655
<< via2 >>
rect 1180 -440 1280 -340
rect 1435 -440 1535 -340
rect 1625 -450 2405 -400
rect 2625 -450 3405 -400
rect 735 -560 955 -525
<< metal3 >>
rect 1180 -335 1280 -185
rect 1435 -335 1535 -185
rect 1175 -340 1285 -335
rect 1175 -440 1180 -340
rect 1280 -440 1285 -340
rect 1175 -445 1285 -440
rect 1430 -340 1540 -335
rect 1430 -440 1435 -340
rect 1535 -440 1540 -340
rect 1430 -445 1540 -440
rect 1615 -400 2415 -340
rect 1615 -450 1625 -400
rect 2405 -450 2415 -400
rect 1615 -455 2415 -450
rect 2615 -400 3415 -340
rect 2615 -450 2625 -400
rect 3405 -450 3415 -400
rect 2615 -455 3415 -450
rect 725 -525 965 -520
rect 725 -560 735 -525
rect 955 -560 965 -525
rect 725 -565 965 -560
rect 920 -1118 965 -565
<< labels >>
rlabel metal1 435 -335 435 -335 1 VDD
port 1 n
rlabel metal2 1065 -815 1065 -815 1 NB1
port 4 n
rlabel metal2 1320 -815 1320 -815 1 NB2
port 5 n
rlabel metal2 2545 -815 2545 -815 1 OUT_IB
port 6 n
rlabel metal2 3550 -815 3550 -815 1 AMP_IB
port 7 n
rlabel metal1 825 -770 825 -770 1 GND
port 12 n
rlabel metal3 920 -1118 965 -1100 1 SF_IB
port 13 n
<< end >>
