magic
tech sky130A
magscale 1 2
timestamp 1718072386
<< nmoslvt >>
rect -1350 9870 650 9900
rect -120 -850 1880 -820
<< ndiff >>
rect -950 10620 650 10670
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10260 650 10290
rect -1350 10230 650 10260
rect -1350 9940 -1300 10230
rect 600 9940 650 10230
rect -1350 9900 650 9940
rect -1350 9830 650 9870
rect -1350 9660 -1270 9830
rect 600 9660 650 9830
rect -1350 9640 650 9660
rect 280 -140 1880 -120
rect 280 -420 300 -140
rect 1860 -420 1880 -140
rect 280 -430 1880 -420
rect -120 -480 1880 -430
rect -120 -770 30 -480
rect 1810 -770 1880 -480
rect -120 -820 1880 -770
rect -120 -870 1880 -850
rect -120 -1050 -100 -870
rect 620 -880 1880 -870
rect 1860 -1050 1880 -880
rect -120 -1080 1880 -1050
<< ndiffc >>
rect -930 10290 630 10620
rect -1300 9940 600 10230
rect -1270 9660 600 9830
rect 300 -420 1860 -140
rect 30 -770 1810 -480
rect -100 -880 620 -870
rect -100 -1050 1860 -880
<< psubdiff >>
rect -1350 9590 650 9640
rect -1350 9480 -1270 9590
rect 600 9480 650 9590
rect -1350 9440 650 9480
rect -120 -1110 1880 -1080
rect -120 -1300 310 -1110
rect 280 -1360 310 -1300
rect 1850 -1360 1880 -1110
rect 280 -1560 1880 -1360
<< psubdiffcont >>
rect -1270 9480 600 9590
rect 310 -1360 1850 -1110
<< poly >>
rect -1610 10040 -1460 10060
rect -1610 9880 -1600 10040
rect -1470 9900 -1460 10040
rect -1470 9880 -1350 9900
rect -1610 9868 -1527 9880
rect -1493 9870 -1350 9880
rect 650 9870 680 9900
rect -1493 9868 -1460 9870
rect -1610 9850 -1460 9868
rect -217 -818 -163 -802
rect -217 -852 -207 -818
rect -173 -820 -163 -818
rect -173 -850 -120 -820
rect 1880 -850 1910 -820
rect -173 -852 -163 -850
rect -217 -868 -163 -852
<< polycont >>
rect -1600 9880 -1470 10040
rect -1527 9868 -1493 9880
rect -207 -852 -173 -818
<< locali >>
rect -950 10620 650 10650
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10270 650 10290
rect -950 10260 620 10270
rect -1320 10230 620 10260
rect -1610 10055 -1460 10060
rect -1610 9985 -1605 10055
rect -1535 10040 -1460 10055
rect -1610 9880 -1600 9985
rect -1470 9880 -1460 10040
rect -1320 9940 -1300 10230
rect 600 9940 620 10230
rect -1320 9930 620 9940
rect -1610 9868 -1527 9880
rect -1493 9868 -1460 9880
rect -1610 9850 -1460 9868
rect -1320 9830 630 9850
rect -1320 9660 -1270 9830
rect 600 9660 630 9830
rect -1320 9590 630 9660
rect -1320 9270 -1270 9590
rect 600 9270 630 9590
rect -1320 9200 630 9270
rect -400 -250 -90 -240
rect -400 -400 -390 -250
rect -110 -400 -90 -250
rect -400 -410 -90 -400
rect -219 -818 -160 -410
rect 280 -420 300 60
rect 1860 -420 1880 60
rect 280 -430 1880 -420
rect -60 -480 1870 -430
rect -60 -770 30 -480
rect 1810 -770 1870 -480
rect -60 -800 1870 -770
rect -223 -852 -207 -818
rect -173 -852 -157 -818
rect -219 -869 -160 -852
rect -120 -1050 -100 -870
rect 620 -880 1880 -870
rect 1860 -1050 1880 -880
rect -120 -1110 1880 -1050
rect -120 -1300 310 -1110
rect 1850 -1300 1880 -1110
rect 280 -1530 300 -1300
rect 1860 -1530 1880 -1300
rect 280 -1550 1880 -1530
<< viali >>
rect -930 10290 630 10620
rect -1605 10040 -1535 10055
rect -1605 9985 -1600 10040
rect -1600 9880 -1470 10040
rect -1270 9480 600 9590
rect -1270 9270 600 9480
rect -390 -400 -110 -250
rect 300 -140 1860 60
rect 300 -420 1860 -140
rect 300 -1360 310 -1300
rect 310 -1360 1850 -1300
rect 1850 -1360 1860 -1300
rect 300 -1530 1860 -1360
<< metal1 >>
rect 23020 11280 27441 11570
rect -950 10620 650 10630
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10270 650 10290
rect -1611 10060 -1529 10067
rect -2280 10055 -1460 10060
rect -2280 9985 -1605 10055
rect -1535 10040 -1460 10055
rect -2280 9890 -1600 9985
rect -1610 9880 -1600 9890
rect -1470 9880 -1460 10040
rect -1610 9850 -1460 9880
rect -1320 9590 630 9630
rect -1320 9270 -1270 9590
rect 600 9270 630 9590
rect -1320 9200 630 9270
rect 280 60 1880 180
rect -500 -250 100 -240
rect -500 -400 -490 -250
rect -500 -410 -390 -400
rect -110 -410 100 -250
rect 280 -420 300 60
rect 1860 -420 1880 60
rect 280 -430 1880 -420
rect -950 -1290 2500 -1280
rect -950 -1550 -920 -1290
rect 2280 -1550 2500 -1290
rect -950 -1560 2500 -1550
rect -237 -1565 -34 -1560
<< via1 >>
rect -930 10290 630 10620
rect -1270 9270 600 9590
rect -490 -400 -390 -250
rect -390 -400 -110 -250
rect -390 -410 -110 -400
rect 300 -420 1860 60
rect -920 -1300 2280 -1290
rect -920 -1530 300 -1300
rect 300 -1530 1860 -1300
rect 1860 -1530 2280 -1300
rect -920 -1550 2280 -1530
<< metal2 >>
rect -950 10620 650 10630
rect -950 10290 -930 10620
rect 630 10290 650 10620
rect -950 10270 650 10290
rect -950 10269 529 10270
rect -1320 9590 630 9630
rect -1320 9270 -1270 9590
rect 600 9270 630 9590
rect -1320 9200 630 9270
rect 1300 8370 2520 8450
rect 1300 7710 1320 8370
rect 2490 7710 2520 8370
rect 1300 7620 2520 7710
rect 280 3859 1890 3870
rect -1688 3611 2174 3859
rect 280 60 1890 3611
rect -1190 -250 -100 -240
rect -1190 -400 -490 -250
rect -1190 -410 -390 -400
rect -110 -410 -100 -250
rect 280 -420 300 60
rect 1860 -420 1890 60
rect 280 -430 1890 -420
rect -920 -1100 -326 -1036
rect -920 -1280 -878 -1100
rect -950 -1290 -878 -1280
rect -356 -1280 -326 -1100
rect -356 -1290 2490 -1280
rect -950 -1550 -920 -1290
rect 2280 -1550 2490 -1290
rect -950 -1560 -878 -1550
rect -920 -1690 -878 -1560
rect -356 -1560 2490 -1550
rect -356 -1690 -326 -1560
rect -237 -1565 -34 -1560
rect -920 -1796 -326 -1690
<< via2 >>
rect -1270 9270 600 9590
rect 1320 7710 2490 8370
rect -878 -1290 -356 -1100
rect -920 -1550 2280 -1290
rect -878 -1690 -356 -1550
<< metal3 >>
rect -1320 9590 630 9630
rect -1320 9270 -1270 9590
rect 600 9270 630 9590
rect -1320 9200 630 9270
rect -950 -1100 -265 9200
rect 1300 8370 2520 8450
rect 1300 7710 1320 8370
rect 2490 7710 2520 8370
rect 1300 7620 2520 7710
rect -950 -1290 -878 -1100
rect -356 -1256 -265 -1100
rect -356 -1280 -156 -1256
rect -356 -1290 2490 -1280
rect -950 -1550 -920 -1290
rect 2280 -1550 2490 -1290
rect -950 -1690 -878 -1550
rect -356 -1560 2490 -1550
rect -356 -1565 -34 -1560
rect -356 -1636 -156 -1565
rect -356 -1690 -265 -1636
rect -950 -2669 -265 -1690
<< via3 >>
rect 1320 7710 2490 8370
<< metal4 >>
rect -2205 12835 26620 13665
rect -2205 9860 -1375 12835
rect -2205 9180 -1400 9860
rect -2205 8455 -1375 9180
rect -2205 8370 2515 8455
rect -2205 7710 1320 8370
rect 2490 7710 2515 8370
rect -2205 7625 2515 7710
rect 25795 7690 26620 12835
rect 24850 6830 26620 7690
use opamp_v1  opamp_v1_0 fulgor_opamp/
timestamp 1718072386
transform 1 0 -1719 0 1 8388
box 2069 -10028 26971 3199
<< labels >>
rlabel metal4 26418 7258 26418 7258 1 AOUT
port 2 n
rlabel metal1 -2240 9968 -2240 9968 1 AMP_IB
port 4 n
rlabel metal2 -1576 3762 -1576 3762 1 ARRAY_OUT
port 5 n
rlabel metal3 -950 -2669 -265 -1984 1 VSS
port 6 n
rlabel metal1 27151 11280 27441 11570 1 VDD
port 7 n
rlabel metal2 -1078 -314 -1078 -314 1 OUT_IB
port 3 n
<< end >>
