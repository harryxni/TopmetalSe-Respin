magic
tech sky130A
timestamp 1758079492
<< end >>
