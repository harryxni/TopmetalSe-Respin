module shift_register (GND,
    VDD,
    clk,
    data_in,
    data_out,
    ena,
    rst,
    ROW_SEL);
 input GND;
 input VDD;
 input clk;
 input data_in;
 output data_out;
 input ena;
 input rst;
 output [99:0] ROW_SEL;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_0 (.DIODE(_342_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_342_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net104),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net104),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net104),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net104),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net98),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net3),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net99),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net99),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net99),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net1),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1313 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1341 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1369 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1565 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1593 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1621 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1649 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1677 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1733 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1789 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1957 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1985 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2013 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2069 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2085 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2097 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2125 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2153 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2181 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2209 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_221 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2237 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2265 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2293 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2321 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2349 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2377 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2405 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2433 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2461 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2489 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2517 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2545 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2573 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2601 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2629 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2657 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2685 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2713 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2741 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2769 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2797 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2825 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2853 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2881 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2909 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2937 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2965 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2993 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3021 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3049 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3077 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_333 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_361 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_389 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_417 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_445 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_473 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_501 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_529 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_557 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_585 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_613 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_641 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_669 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_697 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_725 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_753 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_781 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_809 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_837 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_865 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_893 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_921 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_949 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_0_977 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_0_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1509 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1533 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_1651 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1677 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1707 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1789 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1957 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_1987 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2069 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2149 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2267 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_10_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_307 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_10_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_475 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_10_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_10_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_10_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_11_10 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_11_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_14 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_1617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1623 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1649 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_11_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_1673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1679 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_11_18 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2041 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2071 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2085 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2097 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2121 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2127 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_22 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_11_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2911 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_335 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_34 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_385 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_11_46 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_11_54 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_11_6 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_11_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_11_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1509 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1533 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_1651 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1677 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1707 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1789 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1957 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_1987 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2069 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2149 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2267 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_12_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_307 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_12_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_475 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_12_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_12_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_13_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1425 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_1513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_1617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1623 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1649 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_13_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_1673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1679 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_1681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2041 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2071 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_2073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2077 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_2081 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2088 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2100 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2112 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_13_2124 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_13_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2893 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_13_2902 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_2910 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_13_317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_13_325 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_335 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_340 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_347 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_359 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_371 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_13_383 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_13_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_13_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_13_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_13_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_13_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1397 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_14_1509 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1534 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_1651 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1677 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1683 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_1704 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1789 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1957 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_1987 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_14_2069 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_2076 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_2083 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_14_2090 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_2098 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2149 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2267 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_14_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_14_2885 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_14_2894 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_14_2901 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_2908 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2915 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2927 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_307 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_14_309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_14_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_14_320 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_327 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_3289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_3295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_334 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_341 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_348 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_14_355 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_475 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_14_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_14_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_14_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_14_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_15_1089 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1096 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1108 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_15_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_1401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1408 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1420 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1432 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1444 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_1513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_15_1605 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_15_1621 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1628 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1640 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1652 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1664 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_1676 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_1681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2021 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2031 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2043 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_15_2055 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_2063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2068 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_2076 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2086 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2094 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_15_2125 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_15_2185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2196 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2208 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2220 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_15_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_15_2232 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2748 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2760 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2772 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2784 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_15_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2796 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_15_2869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2880 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2887 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2894 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2901 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_2908 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2916 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2928 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2940 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2952 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_15_2964 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_15_305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_15_309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_313 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_15_326 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_334 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_340 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_347 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_354 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_366 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_378 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_15_390 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_15_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_15_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_15_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_15_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1109 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1116 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1128 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_16_1140 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1244 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1248 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_1252 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1264 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1276 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1288 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1300 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1312 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_1397 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1405 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1409 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1416 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1423 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1509 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1534 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_1606 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1612 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_1619 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1630 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_16_1642 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_16_1650 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1677 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1683 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1704 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1745 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1752 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1759 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1768 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1780 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1792 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1804 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1816 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1913 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1920 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_1927 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1936 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1948 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1960 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1972 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_1984 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_2045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_2053 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2058 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_2073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_2095 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2110 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_16_2153 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_2181 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2188 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_2202 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_16_2210 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2216 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2228 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2240 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2252 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_2264 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2473 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_2482 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_2490 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_16_2585 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_2593 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_2598 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2608 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2622 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2634 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2646 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_16_2658 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_16_2729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2742 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2756 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_2768 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_16_2865 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2870 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_16_2885 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_2897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_16_2904 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_2908 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_2919 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_2932 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_304 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_16_330 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_355 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_425 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_436 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_443 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_450 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_462 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_16_474 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_592 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_598 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_602 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_614 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_626 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_638 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_822 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_16_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_834 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_16_865 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_928 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_935 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_943 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_950 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_962 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_16_974 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_16_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_16_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_1004 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_1080 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1087 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_1100 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1106 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_1110 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_1118 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_1228 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_1243 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_1254 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1268 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_17_1280 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_1396 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1405 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1415 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1423 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1430 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1442 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_17_1454 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_17_1581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_17_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1599 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1620 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1629 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_1633 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1639 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1650 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1662 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_17_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_1674 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1740 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1747 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1754 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1761 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1768 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1775 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_1782 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_1790 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_1909 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_1917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_1927 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_1940 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1947 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_17_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2041 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_2050 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_2064 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2117 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2124 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2196 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2200 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2210 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2223 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_17_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2235 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2474 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2487 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_2494 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2501 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2508 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2577 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_2585 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_2593 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2604 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_2611 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2618 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_17_2728 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_2732 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_2738 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2754 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2761 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2768 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2780 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_17_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_2792 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_17_281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2857 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2864 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2871 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2908 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_293 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2940 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2952 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_2964 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_306 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_330 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_346 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_364 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_371 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_17_383 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_17_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_408 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_415 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_428 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_437 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_444 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_565 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_574 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_594 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_600 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_604 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_611 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_17_818 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_836 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_844 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_856 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_868 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_880 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_17_892 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_17_897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_908 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_915 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_928 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_17_932 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_937 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_17_956 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_968 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_980 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_17_992 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_1061 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1068 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1075 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1088 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1112 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1126 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_18_1145 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_1220 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1227 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_1251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1270 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_18_1313 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_18_1373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1383 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1387 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_1411 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1424 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1432 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1444 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1456 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1468 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_1480 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1491 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1503 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1515 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1527 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_18_1539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1565 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1571 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_1578 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_18_1586 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1592 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_18_1597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_1603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1611 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1632 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1648 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_18_1653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1666 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1678 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1690 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1702 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_1730 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1745 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_1758 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_1786 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1794 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1806 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_18_1818 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_1889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_18_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1916 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1920 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_1933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_1955 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1962 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1974 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_18_1986 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_2040 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_18_2045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2058 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2082 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_2095 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_2124 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2138 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_2150 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_2169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2176 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_2191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_2202 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_18_2210 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_2257 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_18_2265 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2481 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2488 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2493 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2507 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2514 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2526 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_2538 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_2546 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_18_2573 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2579 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2592 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2599 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2605 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_2615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2621 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2638 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_18_2657 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_2685 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2698 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_2710 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2720 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2724 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2753 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_2766 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_277 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2776 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2783 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2795 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2807 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_18_281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_2819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2844 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_18_2856 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2860 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2880 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_2905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_291 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2929 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_2936 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2950 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2962 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_2974 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_2986 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_2994 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_304 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_353 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_360 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_368 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_375 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_381 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_386 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_394 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_409 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_416 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_434 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_458 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_466 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_474 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_18_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_577 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_584 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_594 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_607 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_614 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_633 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_18_641 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_18_808 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_826 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_18_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_18_852 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_858 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_862 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_893 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_910 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_916 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_920 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_936 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_949 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_956 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_963 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_18_970 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_978 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_18_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_19_1005 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1060 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1086 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_1110 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1118 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_1130 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1138 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1142 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1154 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_1166 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1174 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_19_1201 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1220 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1228 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1237 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_1250 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1274 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_1357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1368 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_1376 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1383 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1396 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1406 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1430 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1434 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1444 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1451 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1463 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1475 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1487 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1499 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_19_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_1537 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1548 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_1560 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_1578 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_1611 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1620 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1629 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1639 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1649 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1657 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1661 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1676 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1685 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1689 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_19_1693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_1709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1713 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1723 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1731 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_1737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1767 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1780 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1788 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1801 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1808 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1815 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1827 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_1839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_1885 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_1889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1893 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1900 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_1949 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1956 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_1964 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_1971 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1983 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1995 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_2007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_19_2029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2033 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2041 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_2049 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_19_2057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2068 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2082 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2109 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_2122 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_2138 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_2157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_2165 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2170 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2210 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_2234 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2244 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2256 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2268 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2280 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_2292 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_2445 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2453 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2460 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_2492 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2516 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2524 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2536 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2548 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_19_2560 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2565 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2572 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_19_2577 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2600 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_2624 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2633 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2641 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2649 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2656 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2668 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_2680 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_19_269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_2701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_2710 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2718 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2723 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_2736 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_274 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2778 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_19_2797 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_2825 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2831 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2836 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2844 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_285 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2852 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2860 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2891 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_2904 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_2946 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_2959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_308 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_3273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_3280 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_3292 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_3296 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_3300 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_332 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_370 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_377 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_383 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_388 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_397 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_410 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_416 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_437 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_444 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_452 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_465 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_471 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_475 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_487 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_499 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_19_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_556 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_566 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_579 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_611 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_19_617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_19_775 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_797 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_801 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_19_829 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_836 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_844 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_851 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_875 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_19_887 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_921 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_19_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_966 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_974 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_19_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_1617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1623 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1649 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_1673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1679 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2041 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2071 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2085 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2097 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2121 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2127 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_1_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_1_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2911 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_335 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_385 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_1_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_1_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_1_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1012 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1024 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1042 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_108 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1088 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1116 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_20_1173 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1180 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_1192 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1196 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1200 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1228 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_1256 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1284 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_1298 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_1329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1340 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1355 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1368 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_137 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1394 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1424 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_144 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_1469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_1476 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_20_1509 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1516 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1528 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1544 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_1556 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_156 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_20_1560 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1564 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1592 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1620 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1648 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1676 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1684 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_1691 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_1699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1704 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1732 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_174 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1802 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_1810 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_1818 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_1833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1843 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_186 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_1861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1872 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_1886 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_1894 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1900 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_194 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_1970 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_1977 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_1985 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_20 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2010 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2027 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2040 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_2045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2068 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_208 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_2096 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2124 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2137 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_2140 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2151 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_2157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2176 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_220 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_2250 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_2262 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_2305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2310 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_20_2322 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_20_2337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_20_237 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_2377 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2384 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_2396 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2412 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2418 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2428 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2437 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2444 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2450 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2460 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_249 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2524 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_2531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_2539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2544 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_2570 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_265 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_20_2673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2677 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_2685 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2689 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_2697 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_276 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2801 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2807 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2811 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_2823 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2829 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2837 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2852 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_2857 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2880 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_29 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2908 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_2972 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_2979 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_2991 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_2997 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_3005 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3011 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_20_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_3037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_304 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_3044 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_20_3077 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3084 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_20_309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3096 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_3112 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_3124 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_3137 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3144 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_3156 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_3165 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3173 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3178 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_20_3190 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_3193 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_3201 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3206 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_3211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_3233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_3244 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_20_3261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3266 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3270 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3274 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_3277 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3283 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3300 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_332 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_360 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_37 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_385 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_416 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_444 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_470 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_486 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_498 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_508 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_520 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 FILLER_20_53 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_533 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_538 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_551 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_584 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_612 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_648 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_660 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_676 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_20_688 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_20_69 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_708 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_20_720 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_74 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_742 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_20_754 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_2 FILLER_20_769 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_780 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_8 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_20_808 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_20_82 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_836 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_20_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_878 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_885 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_892 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_920 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_20_925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_948 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_20_97 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_20_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_20_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_20_981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_20_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1957 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_1987 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2069 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2149 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2267 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_2_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_307 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_2_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_475 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_2_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_2_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_3_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_3_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2911 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_335 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_385 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_3_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_3_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_3_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1957 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2149 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_4_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_307 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_4_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_475 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_4_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_4_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_5_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_5_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_5_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2911 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_335 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_385 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_5_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_5_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_5_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_5_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_5_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_5_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1957 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2149 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_6_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_307 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_6_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_475 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_6_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_6_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_6_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_7_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1649 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_7_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_1673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2041 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2071 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2085 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2097 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2121 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2127 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_7_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_7_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2911 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_3285 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_3300 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_335 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_385 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_7_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_7_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_7_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_7_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_7_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_133 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1565 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1589 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1609 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1621 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1645 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_1651 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1721 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1733 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1757 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1889 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_189 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1901 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1925 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1931 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1945 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1957 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1981 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_1987 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_1989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2001 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2013 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2037 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2043 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2057 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2069 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2093 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2099 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2149 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2155 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2205 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_2211 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2261 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2267 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2317 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2323 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2373 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2379 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2429 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2435 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_245 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2485 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2491 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_251 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2541 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2547 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2597 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2603 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2653 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2659 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_8_2709 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2715 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2765 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_2771 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2821 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2827 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2877 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2883 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_29 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2933 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2939 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_2977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_2989 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_2995 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_2997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_3021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_3045 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_3051 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_3053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_307 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_3077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_3101 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_3107 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_3109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_3157 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_3163 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_3165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_3213 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_3219 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_3221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_3269 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_3275 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_3277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_3289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_8 FILLER_8_3301 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_357 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_363 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_41 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_413 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_419 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_469 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_475 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_525 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_53 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_531 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_581 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_587 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_637 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_643 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_65 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_693 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_699 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_749 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_755 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_77 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_805 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_811 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_8_83 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_85 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_861 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_867 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_917 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_923 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_97 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_8_973 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_979 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_8_981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_8_993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_105 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_9_111 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_113 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_125 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1425 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1437 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1449 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1455 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_15 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1505 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1511 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1537 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1549 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1561 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1567 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1593 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1605 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_161 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_1617 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1623 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1649 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1661 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_1673 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1679 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_169 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1705 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1717 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1729 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1735 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1761 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1773 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1785 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1791 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1805 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_181 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1817 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1829 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1841 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1847 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1873 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1885 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1897 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1903 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1929 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1941 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1953 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_1959 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_1961 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1973 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1985 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1997 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2009 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2015 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2017 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2029 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2041 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2053 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2065 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2071 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2073 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2085 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2097 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2109 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2121 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2127 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2129 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2141 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2153 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2165 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_217 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_2177 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2183 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2185 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2197 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2209 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2221 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_9_223 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_2233 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2239 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2241 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_225 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2253 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2265 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2277 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2289 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2295 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2297 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2309 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2321 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2333 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2345 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2351 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2353 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2365 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_237 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2377 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2389 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2401 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2407 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2409 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2421 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2433 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2445 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2457 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2463 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2465 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2477 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2489 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2501 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2513 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2519 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2521 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2533 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2545 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2557 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2569 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2575 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2577 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2589 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2601 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2613 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2625 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2631 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2633 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2645 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2657 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2669 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2681 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2687 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2689 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_27 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2701 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2713 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2725 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_273 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_2737 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2743 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2745 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2757 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2769 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2781 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_9_279 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_2793 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2799 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2801 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_281 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2813 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2825 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2837 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2849 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2855 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2857 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2869 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2881 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2893 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2905 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2911 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2913 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2925 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_293 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2937 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2949 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_2961 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_2967 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_2969 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2981 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_2993 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3005 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_3017 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_3023 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_3025 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3037 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3049 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_305 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3061 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_3073 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_3079 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_3081 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3093 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3105 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3117 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_3129 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_3135 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_3137 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3149 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3161 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_317 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3173 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_3185 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_3191 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_3193 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3205 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3217 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3229 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_3241 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_3247 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_3249 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3261 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3273 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_3285 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_329 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_3297 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_3303 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_3305 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_335 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_337 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_349 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_361 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_373 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_385 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_39 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_9_391 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_393 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_405 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_417 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_429 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_441 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_447 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_449 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_461 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_473 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_485 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_497 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_503 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_505 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_4 FILLER_9_51 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_517 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_529 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_541 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_553 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_559 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_561 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_57 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_573 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_585 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_597 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_609 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_615 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_617 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_629 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_641 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_653 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_665 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_671 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_673 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_685 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_69 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_697 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_709 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_721 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_727 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_729 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_741 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_753 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_765 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_777 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_783 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_785 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_797 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_809 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_81 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_821 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_833 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_839 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_841 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_853 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_865 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_877 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_889 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_895 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_897 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_909 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_921 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_93 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_933 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_6 FILLER_9_945 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_951 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_9_953 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_965 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_977 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_ef_sc_hd__decap_12 FILLER_9_989 (.VGND(GND),
    .VPWR(VDD),
    .VPB(VDD),
    .VNB(GND));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 (.VGND(GND),
    .VPWR(VDD));
 sky130_fd_sc_hd__buf_4 _348_ (.A(net2),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_2 _349_ (.A(_200_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_201_));
 sky130_fd_sc_hd__mux2_1 _350_ (.A0(net16),
    .A1(net14),
    .S(_201_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_202_));
 sky130_fd_sc_hd__clkbuf_1 _351_ (.A(_202_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_199_));
 sky130_fd_sc_hd__mux2_1 _352_ (.A0(net14),
    .A1(net13),
    .S(_201_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _353_ (.A(_203_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_198_));
 sky130_fd_sc_hd__mux2_1 _354_ (.A0(net13),
    .A1(net12),
    .S(_201_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_204_));
 sky130_fd_sc_hd__clkbuf_1 _355_ (.A(_204_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_197_));
 sky130_fd_sc_hd__mux2_1 _356_ (.A0(net12),
    .A1(net11),
    .S(_201_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_205_));
 sky130_fd_sc_hd__clkbuf_1 _357_ (.A(_205_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_196_));
 sky130_fd_sc_hd__mux2_1 _358_ (.A0(net11),
    .A1(net10),
    .S(_201_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_206_));
 sky130_fd_sc_hd__clkbuf_1 _359_ (.A(_206_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_195_));
 sky130_fd_sc_hd__clkbuf_2 _360_ (.A(_200_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_207_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(net10),
    .A1(net9),
    .S(_207_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_208_));
 sky130_fd_sc_hd__clkbuf_1 _362_ (.A(_208_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_194_));
 sky130_fd_sc_hd__mux2_1 _363_ (.A0(net9),
    .A1(net8),
    .S(_207_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_209_));
 sky130_fd_sc_hd__clkbuf_1 _364_ (.A(_209_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_193_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(net8),
    .A1(net7),
    .S(_207_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_210_));
 sky130_fd_sc_hd__clkbuf_1 _366_ (.A(_210_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_192_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(net7),
    .A1(net6),
    .S(_207_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_1 _368_ (.A(_211_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_191_));
 sky130_fd_sc_hd__mux2_1 _369_ (.A0(net6),
    .A1(net5),
    .S(_207_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_212_));
 sky130_fd_sc_hd__clkbuf_1 _370_ (.A(_212_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_190_));
 sky130_fd_sc_hd__clkbuf_2 _371_ (.A(_200_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_213_));
 sky130_fd_sc_hd__mux2_1 _372_ (.A0(net5),
    .A1(net103),
    .S(_213_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_214_));
 sky130_fd_sc_hd__clkbuf_1 _373_ (.A(_214_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_189_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(net103),
    .A1(net92),
    .S(_213_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_215_));
 sky130_fd_sc_hd__clkbuf_1 _375_ (.A(_215_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_188_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(net92),
    .A1(net81),
    .S(_213_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_216_));
 sky130_fd_sc_hd__clkbuf_1 _377_ (.A(_216_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_187_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(net81),
    .A1(net70),
    .S(_213_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_217_));
 sky130_fd_sc_hd__clkbuf_1 _379_ (.A(_217_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_186_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(net70),
    .A1(net59),
    .S(_213_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_218_));
 sky130_fd_sc_hd__clkbuf_1 _381_ (.A(_218_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_185_));
 sky130_fd_sc_hd__clkbuf_2 _382_ (.A(_200_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_219_));
 sky130_fd_sc_hd__mux2_1 _383_ (.A0(net59),
    .A1(net48),
    .S(_219_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_220_));
 sky130_fd_sc_hd__clkbuf_1 _384_ (.A(_220_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_184_));
 sky130_fd_sc_hd__mux2_1 _385_ (.A0(net48),
    .A1(net37),
    .S(_219_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_221_));
 sky130_fd_sc_hd__clkbuf_1 _386_ (.A(_221_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_183_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(net37),
    .A1(net26),
    .S(_219_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_222_));
 sky130_fd_sc_hd__clkbuf_1 _388_ (.A(_222_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_182_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(net26),
    .A1(net15),
    .S(_219_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_223_));
 sky130_fd_sc_hd__clkbuf_1 _390_ (.A(_223_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_181_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(net15),
    .A1(net4),
    .S(_219_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_224_));
 sky130_fd_sc_hd__clkbuf_1 _392_ (.A(_224_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_180_));
 sky130_fd_sc_hd__clkbuf_4 _393_ (.A(_200_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_225_));
 sky130_fd_sc_hd__mux2_1 _394_ (.A0(net4),
    .A1(net1),
    .S(_225_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_226_));
 sky130_fd_sc_hd__clkbuf_1 _395_ (.A(_226_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_179_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(net102),
    .A1(net101),
    .S(_225_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_227_));
 sky130_fd_sc_hd__clkbuf_1 _397_ (.A(_227_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_178_));
 sky130_fd_sc_hd__mux2_1 _398_ (.A0(net101),
    .A1(net100),
    .S(_225_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_228_));
 sky130_fd_sc_hd__clkbuf_1 _399_ (.A(_228_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_177_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(net100),
    .A1(net99),
    .S(_225_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_229_));
 sky130_fd_sc_hd__clkbuf_1 _401_ (.A(_229_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_176_));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(net99),
    .A1(net98),
    .S(_225_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_230_));
 sky130_fd_sc_hd__clkbuf_1 _403_ (.A(_230_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_175_));
 sky130_fd_sc_hd__clkbuf_2 _404_ (.A(net2),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_231_));
 sky130_fd_sc_hd__clkbuf_2 _405_ (.A(_231_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_232_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(net98),
    .A1(net97),
    .S(_232_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_233_));
 sky130_fd_sc_hd__clkbuf_1 _407_ (.A(_233_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_174_));
 sky130_fd_sc_hd__mux2_1 _408_ (.A0(net97),
    .A1(net96),
    .S(_232_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_234_));
 sky130_fd_sc_hd__clkbuf_1 _409_ (.A(_234_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_173_));
 sky130_fd_sc_hd__mux2_1 _410_ (.A0(net96),
    .A1(net95),
    .S(_232_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_235_));
 sky130_fd_sc_hd__clkbuf_1 _411_ (.A(_235_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_172_));
 sky130_fd_sc_hd__mux2_1 _412_ (.A0(net95),
    .A1(net94),
    .S(_232_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_236_));
 sky130_fd_sc_hd__clkbuf_1 _413_ (.A(_236_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_171_));
 sky130_fd_sc_hd__mux2_1 _414_ (.A0(net94),
    .A1(net93),
    .S(_232_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_237_));
 sky130_fd_sc_hd__clkbuf_1 _415_ (.A(_237_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_170_));
 sky130_fd_sc_hd__clkbuf_2 _416_ (.A(_231_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_238_));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(net93),
    .A1(net91),
    .S(_238_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_1 _418_ (.A(_239_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_169_));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(net91),
    .A1(net90),
    .S(_238_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_240_));
 sky130_fd_sc_hd__clkbuf_1 _420_ (.A(_240_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_168_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(net90),
    .A1(net89),
    .S(_238_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_241_));
 sky130_fd_sc_hd__clkbuf_1 _422_ (.A(_241_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_167_));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(net89),
    .A1(net88),
    .S(_238_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_242_));
 sky130_fd_sc_hd__clkbuf_1 _424_ (.A(_242_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_166_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(net88),
    .A1(net87),
    .S(_238_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_243_));
 sky130_fd_sc_hd__clkbuf_1 _426_ (.A(_243_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_165_));
 sky130_fd_sc_hd__clkbuf_2 _427_ (.A(_231_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_244_));
 sky130_fd_sc_hd__mux2_1 _428_ (.A0(net87),
    .A1(net86),
    .S(_244_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_245_));
 sky130_fd_sc_hd__clkbuf_1 _429_ (.A(_245_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_164_));
 sky130_fd_sc_hd__mux2_1 _430_ (.A0(net86),
    .A1(net85),
    .S(_244_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_246_));
 sky130_fd_sc_hd__clkbuf_1 _431_ (.A(_246_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_163_));
 sky130_fd_sc_hd__mux2_1 _432_ (.A0(net85),
    .A1(net84),
    .S(_244_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_247_));
 sky130_fd_sc_hd__clkbuf_1 _433_ (.A(_247_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _434_ (.A0(net84),
    .A1(net83),
    .S(_244_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_248_));
 sky130_fd_sc_hd__clkbuf_1 _435_ (.A(_248_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_161_));
 sky130_fd_sc_hd__mux2_1 _436_ (.A0(net83),
    .A1(net82),
    .S(_244_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_249_));
 sky130_fd_sc_hd__clkbuf_1 _437_ (.A(_249_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_160_));
 sky130_fd_sc_hd__clkbuf_2 _438_ (.A(_231_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_250_));
 sky130_fd_sc_hd__mux2_1 _439_ (.A0(net82),
    .A1(net80),
    .S(_250_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_251_));
 sky130_fd_sc_hd__clkbuf_1 _440_ (.A(_251_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_159_));
 sky130_fd_sc_hd__mux2_1 _441_ (.A0(net80),
    .A1(net79),
    .S(_250_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_252_));
 sky130_fd_sc_hd__clkbuf_1 _442_ (.A(_252_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(net79),
    .A1(net78),
    .S(_250_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_253_));
 sky130_fd_sc_hd__clkbuf_1 _444_ (.A(_253_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(net78),
    .A1(net77),
    .S(_250_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_254_));
 sky130_fd_sc_hd__clkbuf_1 _446_ (.A(_254_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(net77),
    .A1(net76),
    .S(_250_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_255_));
 sky130_fd_sc_hd__clkbuf_1 _448_ (.A(_255_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_155_));
 sky130_fd_sc_hd__clkbuf_2 _449_ (.A(_231_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_256_));
 sky130_fd_sc_hd__mux2_1 _450_ (.A0(net76),
    .A1(net75),
    .S(_256_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_257_));
 sky130_fd_sc_hd__clkbuf_1 _451_ (.A(_257_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_154_));
 sky130_fd_sc_hd__mux2_1 _452_ (.A0(net75),
    .A1(net74),
    .S(_256_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_258_));
 sky130_fd_sc_hd__clkbuf_1 _453_ (.A(_258_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _454_ (.A0(net74),
    .A1(net73),
    .S(_256_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_259_));
 sky130_fd_sc_hd__clkbuf_1 _455_ (.A(_259_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _456_ (.A0(net73),
    .A1(net72),
    .S(_256_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_260_));
 sky130_fd_sc_hd__clkbuf_1 _457_ (.A(_260_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_151_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(net72),
    .A1(net71),
    .S(_256_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_261_));
 sky130_fd_sc_hd__clkbuf_1 _459_ (.A(_261_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_150_));
 sky130_fd_sc_hd__clkbuf_2 _460_ (.A(net2),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_262_));
 sky130_fd_sc_hd__clkbuf_2 _461_ (.A(_262_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_263_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(net71),
    .A1(net69),
    .S(_263_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_264_));
 sky130_fd_sc_hd__clkbuf_1 _463_ (.A(_264_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _464_ (.A0(net69),
    .A1(net68),
    .S(_263_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_265_));
 sky130_fd_sc_hd__clkbuf_1 _465_ (.A(_265_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _466_ (.A0(net68),
    .A1(net67),
    .S(_263_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_266_));
 sky130_fd_sc_hd__clkbuf_1 _467_ (.A(_266_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(net67),
    .A1(net66),
    .S(_263_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_267_));
 sky130_fd_sc_hd__clkbuf_1 _469_ (.A(_267_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(net66),
    .A1(net65),
    .S(_263_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_268_));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(_268_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_145_));
 sky130_fd_sc_hd__clkbuf_2 _472_ (.A(_262_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_269_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(net65),
    .A1(net64),
    .S(_269_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_270_));
 sky130_fd_sc_hd__clkbuf_1 _474_ (.A(_270_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(net64),
    .A1(net63),
    .S(_269_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_271_));
 sky130_fd_sc_hd__clkbuf_1 _476_ (.A(_271_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(net63),
    .A1(net62),
    .S(_269_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_272_));
 sky130_fd_sc_hd__clkbuf_1 _478_ (.A(_272_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _479_ (.A0(net62),
    .A1(net61),
    .S(_269_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_273_));
 sky130_fd_sc_hd__clkbuf_1 _480_ (.A(_273_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_141_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(net61),
    .A1(net60),
    .S(_269_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_274_));
 sky130_fd_sc_hd__clkbuf_1 _482_ (.A(_274_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_140_));
 sky130_fd_sc_hd__clkbuf_2 _483_ (.A(_262_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_275_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(net60),
    .A1(net58),
    .S(_275_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_276_));
 sky130_fd_sc_hd__clkbuf_1 _485_ (.A(_276_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _486_ (.A0(net58),
    .A1(net57),
    .S(_275_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_277_));
 sky130_fd_sc_hd__clkbuf_1 _487_ (.A(_277_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _488_ (.A0(net57),
    .A1(net56),
    .S(_275_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_278_));
 sky130_fd_sc_hd__clkbuf_1 _489_ (.A(_278_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_137_));
 sky130_fd_sc_hd__mux2_1 _490_ (.A0(net56),
    .A1(net55),
    .S(_275_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_279_));
 sky130_fd_sc_hd__clkbuf_1 _491_ (.A(_279_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _492_ (.A0(net55),
    .A1(net54),
    .S(_275_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_280_));
 sky130_fd_sc_hd__clkbuf_1 _493_ (.A(_280_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_135_));
 sky130_fd_sc_hd__clkbuf_2 _494_ (.A(_262_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_281_));
 sky130_fd_sc_hd__mux2_1 _495_ (.A0(net54),
    .A1(net53),
    .S(_281_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_282_));
 sky130_fd_sc_hd__clkbuf_1 _496_ (.A(_282_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _497_ (.A0(net53),
    .A1(net52),
    .S(_281_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_283_));
 sky130_fd_sc_hd__clkbuf_1 _498_ (.A(_283_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(net52),
    .A1(net51),
    .S(_281_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_284_));
 sky130_fd_sc_hd__clkbuf_1 _500_ (.A(_284_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _501_ (.A0(net51),
    .A1(net50),
    .S(_281_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_285_));
 sky130_fd_sc_hd__clkbuf_1 _502_ (.A(_285_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _503_ (.A0(net50),
    .A1(net49),
    .S(_281_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_286_));
 sky130_fd_sc_hd__clkbuf_1 _504_ (.A(_286_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_130_));
 sky130_fd_sc_hd__clkbuf_2 _505_ (.A(_262_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_287_));
 sky130_fd_sc_hd__mux2_1 _506_ (.A0(net49),
    .A1(net47),
    .S(_287_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_288_));
 sky130_fd_sc_hd__clkbuf_1 _507_ (.A(_288_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _508_ (.A0(net47),
    .A1(net46),
    .S(_287_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_289_));
 sky130_fd_sc_hd__clkbuf_1 _509_ (.A(_289_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _510_ (.A0(net46),
    .A1(net45),
    .S(_287_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_290_));
 sky130_fd_sc_hd__clkbuf_1 _511_ (.A(_290_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _512_ (.A0(net45),
    .A1(net44),
    .S(_287_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_291_));
 sky130_fd_sc_hd__clkbuf_1 _513_ (.A(_291_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _514_ (.A0(net44),
    .A1(net43),
    .S(_287_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_292_));
 sky130_fd_sc_hd__clkbuf_1 _515_ (.A(_292_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_125_));
 sky130_fd_sc_hd__buf_2 _516_ (.A(net2),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_293_));
 sky130_fd_sc_hd__clkbuf_2 _517_ (.A(_293_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_294_));
 sky130_fd_sc_hd__mux2_1 _518_ (.A0(net43),
    .A1(net42),
    .S(_294_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_295_));
 sky130_fd_sc_hd__clkbuf_1 _519_ (.A(_295_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _520_ (.A0(net42),
    .A1(net41),
    .S(_294_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_296_));
 sky130_fd_sc_hd__clkbuf_1 _521_ (.A(_296_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _522_ (.A0(net41),
    .A1(net40),
    .S(_294_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_297_));
 sky130_fd_sc_hd__clkbuf_1 _523_ (.A(_297_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _524_ (.A0(net40),
    .A1(net39),
    .S(_294_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_298_));
 sky130_fd_sc_hd__clkbuf_1 _525_ (.A(_298_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _526_ (.A0(net39),
    .A1(net38),
    .S(_294_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_299_));
 sky130_fd_sc_hd__clkbuf_1 _527_ (.A(_299_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_120_));
 sky130_fd_sc_hd__clkbuf_2 _528_ (.A(_293_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_300_));
 sky130_fd_sc_hd__mux2_1 _529_ (.A0(net38),
    .A1(net36),
    .S(_300_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_301_));
 sky130_fd_sc_hd__clkbuf_1 _530_ (.A(_301_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _531_ (.A0(net36),
    .A1(net35),
    .S(_300_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_302_));
 sky130_fd_sc_hd__clkbuf_1 _532_ (.A(_302_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _533_ (.A0(net35),
    .A1(net34),
    .S(_300_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_303_));
 sky130_fd_sc_hd__clkbuf_1 _534_ (.A(_303_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _535_ (.A0(net34),
    .A1(net33),
    .S(_300_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_304_));
 sky130_fd_sc_hd__clkbuf_1 _536_ (.A(_304_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _537_ (.A0(net33),
    .A1(net32),
    .S(_300_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_305_));
 sky130_fd_sc_hd__clkbuf_1 _538_ (.A(_305_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_115_));
 sky130_fd_sc_hd__clkbuf_2 _539_ (.A(_293_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_306_));
 sky130_fd_sc_hd__mux2_1 _540_ (.A0(net32),
    .A1(net31),
    .S(_306_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_307_));
 sky130_fd_sc_hd__clkbuf_1 _541_ (.A(_307_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _542_ (.A0(net31),
    .A1(net30),
    .S(_306_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_308_));
 sky130_fd_sc_hd__clkbuf_1 _543_ (.A(_308_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _544_ (.A0(net30),
    .A1(net29),
    .S(_306_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_309_));
 sky130_fd_sc_hd__clkbuf_1 _545_ (.A(_309_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_112_));
 sky130_fd_sc_hd__mux2_1 _546_ (.A0(net29),
    .A1(net28),
    .S(_306_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_310_));
 sky130_fd_sc_hd__clkbuf_1 _547_ (.A(_310_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _548_ (.A0(net28),
    .A1(net27),
    .S(_306_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_311_));
 sky130_fd_sc_hd__clkbuf_1 _549_ (.A(_311_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_110_));
 sky130_fd_sc_hd__clkbuf_2 _550_ (.A(_293_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_312_));
 sky130_fd_sc_hd__mux2_1 _551_ (.A0(net27),
    .A1(net25),
    .S(_312_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_313_));
 sky130_fd_sc_hd__clkbuf_1 _552_ (.A(_313_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_109_));
 sky130_fd_sc_hd__mux2_1 _553_ (.A0(net25),
    .A1(net24),
    .S(_312_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_314_));
 sky130_fd_sc_hd__clkbuf_1 _554_ (.A(_314_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _555_ (.A0(net24),
    .A1(net23),
    .S(_312_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_315_));
 sky130_fd_sc_hd__clkbuf_1 _556_ (.A(_315_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _557_ (.A0(net23),
    .A1(net22),
    .S(_312_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_316_));
 sky130_fd_sc_hd__clkbuf_1 _558_ (.A(_316_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _559_ (.A0(net22),
    .A1(net21),
    .S(_312_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_317_));
 sky130_fd_sc_hd__clkbuf_1 _560_ (.A(_317_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_105_));
 sky130_fd_sc_hd__clkbuf_2 _561_ (.A(_293_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_318_));
 sky130_fd_sc_hd__mux2_1 _562_ (.A0(net21),
    .A1(net20),
    .S(_318_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_319_));
 sky130_fd_sc_hd__clkbuf_1 _563_ (.A(_319_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _564_ (.A0(net20),
    .A1(net19),
    .S(_318_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_320_));
 sky130_fd_sc_hd__clkbuf_1 _565_ (.A(_320_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _566_ (.A0(net19),
    .A1(net18),
    .S(_318_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_321_));
 sky130_fd_sc_hd__clkbuf_1 _567_ (.A(_321_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _568_ (.A0(net18),
    .A1(net17),
    .S(_318_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_322_));
 sky130_fd_sc_hd__clkbuf_1 _569_ (.A(_322_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _570_ (.A0(net17),
    .A1(net16),
    .S(_318_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_323_));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(_323_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_100_));
 sky130_fd_sc_hd__buf_2 _572_ (.A(net3),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_324_));
 sky130_fd_sc_hd__buf_2 _573_ (.A(_324_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_325_));
 sky130_fd_sc_hd__inv_2 _574_ (.A(_325_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _575_ (.A(_325_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _576_ (.A(_325_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _577_ (.A(_325_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _578_ (.A(_325_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_004_));
 sky130_fd_sc_hd__clkbuf_2 _579_ (.A(_324_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_326_));
 sky130_fd_sc_hd__inv_2 _580_ (.A(_326_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _581_ (.A(_326_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _582_ (.A(_326_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(_326_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _584_ (.A(_326_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_009_));
 sky130_fd_sc_hd__clkbuf_2 _585_ (.A(_324_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_327_));
 sky130_fd_sc_hd__inv_2 _586_ (.A(_327_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _587_ (.A(_327_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _588_ (.A(_327_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _589_ (.A(_327_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _590_ (.A(_327_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_014_));
 sky130_fd_sc_hd__clkbuf_2 _591_ (.A(_324_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_328_));
 sky130_fd_sc_hd__inv_2 _592_ (.A(_328_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _593_ (.A(_328_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _594_ (.A(_328_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _595_ (.A(_328_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _596_ (.A(_328_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_019_));
 sky130_fd_sc_hd__clkbuf_2 _597_ (.A(_324_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_329_));
 sky130_fd_sc_hd__inv_2 _598_ (.A(_329_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _599_ (.A(_329_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _600_ (.A(_329_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _601_ (.A(_329_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _602_ (.A(_329_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_024_));
 sky130_fd_sc_hd__clkbuf_2 _603_ (.A(net3),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_330_));
 sky130_fd_sc_hd__buf_2 _604_ (.A(_330_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_331_));
 sky130_fd_sc_hd__inv_2 _605_ (.A(_331_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _606_ (.A(_331_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _607_ (.A(_331_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _608_ (.A(_331_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _609_ (.A(_331_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_029_));
 sky130_fd_sc_hd__clkbuf_2 _610_ (.A(_330_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_332_));
 sky130_fd_sc_hd__inv_2 _611_ (.A(_332_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _612_ (.A(_332_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _613_ (.A(_332_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _614_ (.A(_332_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _615_ (.A(_332_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_034_));
 sky130_fd_sc_hd__clkbuf_2 _616_ (.A(_330_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_333_));
 sky130_fd_sc_hd__inv_2 _617_ (.A(_333_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _618_ (.A(_333_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _619_ (.A(_333_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _620_ (.A(_333_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _621_ (.A(_333_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_039_));
 sky130_fd_sc_hd__clkbuf_2 _622_ (.A(_330_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_334_));
 sky130_fd_sc_hd__inv_2 _623_ (.A(_334_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _624_ (.A(_334_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _625_ (.A(_334_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _626_ (.A(_334_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _627_ (.A(_334_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_044_));
 sky130_fd_sc_hd__buf_2 _628_ (.A(_330_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_335_));
 sky130_fd_sc_hd__inv_2 _629_ (.A(_335_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _630_ (.A(_335_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _631_ (.A(_335_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _632_ (.A(_335_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _633_ (.A(_335_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_049_));
 sky130_fd_sc_hd__clkbuf_2 _634_ (.A(net3),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_336_));
 sky130_fd_sc_hd__buf_2 _635_ (.A(_336_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_337_));
 sky130_fd_sc_hd__inv_2 _636_ (.A(_337_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _637_ (.A(_337_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _638_ (.A(_337_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _639_ (.A(_337_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _640_ (.A(_337_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_054_));
 sky130_fd_sc_hd__clkbuf_2 _641_ (.A(_336_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_338_));
 sky130_fd_sc_hd__inv_2 _642_ (.A(_338_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _643_ (.A(_338_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _644_ (.A(_338_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _645_ (.A(_338_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _646_ (.A(_338_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_059_));
 sky130_fd_sc_hd__clkbuf_2 _647_ (.A(_336_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_339_));
 sky130_fd_sc_hd__inv_2 _648_ (.A(_339_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _649_ (.A(_339_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _650_ (.A(_339_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _651_ (.A(_339_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _652_ (.A(_339_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_064_));
 sky130_fd_sc_hd__clkbuf_2 _653_ (.A(_336_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_340_));
 sky130_fd_sc_hd__inv_2 _654_ (.A(_340_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _655_ (.A(_340_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _656_ (.A(_340_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _657_ (.A(_340_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _658_ (.A(_340_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_069_));
 sky130_fd_sc_hd__clkbuf_2 _659_ (.A(_336_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_341_));
 sky130_fd_sc_hd__inv_2 _660_ (.A(_341_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _661_ (.A(_341_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _662_ (.A(_341_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _663_ (.A(_341_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _664_ (.A(_341_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_074_));
 sky130_fd_sc_hd__buf_4 _665_ (.A(net3),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_342_));
 sky130_fd_sc_hd__clkbuf_4 _666_ (.A(_342_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_343_));
 sky130_fd_sc_hd__inv_2 _667_ (.A(_343_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _668_ (.A(_343_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _669_ (.A(_343_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _670_ (.A(_343_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _671_ (.A(_343_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_079_));
 sky130_fd_sc_hd__clkbuf_2 _672_ (.A(_342_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_344_));
 sky130_fd_sc_hd__inv_2 _673_ (.A(_344_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _674_ (.A(_344_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _675_ (.A(_344_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _676_ (.A(_344_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _677_ (.A(_344_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_084_));
 sky130_fd_sc_hd__clkbuf_2 _678_ (.A(_342_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_345_));
 sky130_fd_sc_hd__inv_2 _679_ (.A(_345_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _680_ (.A(_345_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _681_ (.A(_345_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _682_ (.A(_345_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _683_ (.A(_345_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_089_));
 sky130_fd_sc_hd__clkbuf_2 _684_ (.A(_342_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_346_));
 sky130_fd_sc_hd__inv_2 _685_ (.A(_346_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _686_ (.A(_346_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _687_ (.A(_346_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _688_ (.A(_346_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _689_ (.A(_346_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_094_));
 sky130_fd_sc_hd__clkbuf_2 _690_ (.A(_342_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(_347_));
 sky130_fd_sc_hd__inv_2 _691_ (.A(_347_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _692_ (.A(_347_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _693_ (.A(_347_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _694_ (.A(_347_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _695_ (.A(_347_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(_099_));
 sky130_fd_sc_hd__dfrtp_1 _696_ (.CLK(clknet_3_2__leaf_clk),
    .D(_100_),
    .RESET_B(_000_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _697_ (.CLK(clknet_3_3__leaf_clk),
    .D(_101_),
    .RESET_B(_001_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _698_ (.CLK(clknet_3_1__leaf_clk),
    .D(_102_),
    .RESET_B(_002_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _699_ (.CLK(clknet_3_2__leaf_clk),
    .D(_103_),
    .RESET_B(_003_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _700_ (.CLK(clknet_3_3__leaf_clk),
    .D(_104_),
    .RESET_B(_004_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _701_ (.CLK(clknet_3_1__leaf_clk),
    .D(_105_),
    .RESET_B(_005_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _702_ (.CLK(clknet_3_3__leaf_clk),
    .D(_106_),
    .RESET_B(_006_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _703_ (.CLK(clknet_3_1__leaf_clk),
    .D(_107_),
    .RESET_B(_007_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _704_ (.CLK(clknet_3_3__leaf_clk),
    .D(_108_),
    .RESET_B(_008_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _705_ (.CLK(clknet_3_3__leaf_clk),
    .D(_109_),
    .RESET_B(_009_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _706_ (.CLK(clknet_3_3__leaf_clk),
    .D(_110_),
    .RESET_B(_010_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _707_ (.CLK(clknet_3_3__leaf_clk),
    .D(_111_),
    .RESET_B(_011_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _708_ (.CLK(clknet_3_3__leaf_clk),
    .D(_112_),
    .RESET_B(_012_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _709_ (.CLK(clknet_3_3__leaf_clk),
    .D(_113_),
    .RESET_B(_013_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _710_ (.CLK(clknet_3_3__leaf_clk),
    .D(_114_),
    .RESET_B(_014_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _711_ (.CLK(clknet_3_2__leaf_clk),
    .D(_115_),
    .RESET_B(_015_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _712_ (.CLK(clknet_3_0__leaf_clk),
    .D(_116_),
    .RESET_B(_016_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _713_ (.CLK(clknet_3_2__leaf_clk),
    .D(_117_),
    .RESET_B(_017_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _714_ (.CLK(clknet_3_2__leaf_clk),
    .D(_118_),
    .RESET_B(_018_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_1 _715_ (.CLK(clknet_3_1__leaf_clk),
    .D(_119_),
    .RESET_B(_019_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _716_ (.CLK(clknet_3_2__leaf_clk),
    .D(_120_),
    .RESET_B(_020_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _717_ (.CLK(clknet_3_0__leaf_clk),
    .D(_121_),
    .RESET_B(_021_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _718_ (.CLK(clknet_3_2__leaf_clk),
    .D(_122_),
    .RESET_B(_022_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _719_ (.CLK(clknet_3_2__leaf_clk),
    .D(_123_),
    .RESET_B(_023_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _720_ (.CLK(clknet_3_2__leaf_clk),
    .D(_124_),
    .RESET_B(_024_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _721_ (.CLK(clknet_3_2__leaf_clk),
    .D(_125_),
    .RESET_B(_025_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _722_ (.CLK(clknet_3_2__leaf_clk),
    .D(_126_),
    .RESET_B(_026_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _723_ (.CLK(clknet_3_3__leaf_clk),
    .D(_127_),
    .RESET_B(_027_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_1 _724_ (.CLK(clknet_3_6__leaf_clk),
    .D(_128_),
    .RESET_B(_028_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _725_ (.CLK(clknet_3_7__leaf_clk),
    .D(_129_),
    .RESET_B(_029_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _726_ (.CLK(clknet_3_7__leaf_clk),
    .D(_130_),
    .RESET_B(_030_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _727_ (.CLK(clknet_3_6__leaf_clk),
    .D(_131_),
    .RESET_B(_031_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _728_ (.CLK(clknet_3_7__leaf_clk),
    .D(_132_),
    .RESET_B(_032_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _729_ (.CLK(clknet_3_7__leaf_clk),
    .D(_133_),
    .RESET_B(_033_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _730_ (.CLK(clknet_3_5__leaf_clk),
    .D(_134_),
    .RESET_B(_034_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _731_ (.CLK(clknet_3_7__leaf_clk),
    .D(_135_),
    .RESET_B(_035_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _732_ (.CLK(clknet_3_7__leaf_clk),
    .D(_136_),
    .RESET_B(_036_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _733_ (.CLK(clknet_3_6__leaf_clk),
    .D(_137_),
    .RESET_B(_037_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _734_ (.CLK(clknet_3_7__leaf_clk),
    .D(_138_),
    .RESET_B(_038_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _735_ (.CLK(clknet_3_4__leaf_clk),
    .D(_139_),
    .RESET_B(_039_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _736_ (.CLK(clknet_3_7__leaf_clk),
    .D(_140_),
    .RESET_B(_040_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _737_ (.CLK(clknet_3_4__leaf_clk),
    .D(_141_),
    .RESET_B(_041_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _738_ (.CLK(clknet_3_4__leaf_clk),
    .D(_142_),
    .RESET_B(_042_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _739_ (.CLK(clknet_3_4__leaf_clk),
    .D(_143_),
    .RESET_B(_043_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _740_ (.CLK(clknet_3_4__leaf_clk),
    .D(_144_),
    .RESET_B(_044_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 _741_ (.CLK(clknet_3_5__leaf_clk),
    .D(_145_),
    .RESET_B(_045_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _742_ (.CLK(clknet_3_5__leaf_clk),
    .D(_146_),
    .RESET_B(_046_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _743_ (.CLK(clknet_3_5__leaf_clk),
    .D(_147_),
    .RESET_B(_047_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _744_ (.CLK(clknet_3_7__leaf_clk),
    .D(_148_),
    .RESET_B(_048_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _745_ (.CLK(clknet_3_4__leaf_clk),
    .D(_149_),
    .RESET_B(_049_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _746_ (.CLK(clknet_3_7__leaf_clk),
    .D(_150_),
    .RESET_B(_050_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _747_ (.CLK(clknet_3_7__leaf_clk),
    .D(_151_),
    .RESET_B(_051_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _748_ (.CLK(clknet_3_4__leaf_clk),
    .D(_152_),
    .RESET_B(_052_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _749_ (.CLK(clknet_3_5__leaf_clk),
    .D(_153_),
    .RESET_B(_053_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _750_ (.CLK(clknet_3_6__leaf_clk),
    .D(_154_),
    .RESET_B(_054_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _751_ (.CLK(clknet_3_6__leaf_clk),
    .D(_155_),
    .RESET_B(_055_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _752_ (.CLK(clknet_3_6__leaf_clk),
    .D(_156_),
    .RESET_B(_056_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _753_ (.CLK(clknet_3_5__leaf_clk),
    .D(_157_),
    .RESET_B(_057_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _754_ (.CLK(clknet_3_6__leaf_clk),
    .D(_158_),
    .RESET_B(_058_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _755_ (.CLK(clknet_3_5__leaf_clk),
    .D(_159_),
    .RESET_B(_059_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _756_ (.CLK(clknet_3_6__leaf_clk),
    .D(_160_),
    .RESET_B(_060_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _757_ (.CLK(clknet_3_7__leaf_clk),
    .D(_161_),
    .RESET_B(_061_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _758_ (.CLK(clknet_3_4__leaf_clk),
    .D(_162_),
    .RESET_B(_062_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _759_ (.CLK(clknet_3_7__leaf_clk),
    .D(_163_),
    .RESET_B(_063_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _760_ (.CLK(clknet_3_7__leaf_clk),
    .D(_164_),
    .RESET_B(_064_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _761_ (.CLK(clknet_3_6__leaf_clk),
    .D(_165_),
    .RESET_B(_065_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _762_ (.CLK(clknet_3_7__leaf_clk),
    .D(_166_),
    .RESET_B(_066_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _763_ (.CLK(clknet_3_4__leaf_clk),
    .D(_167_),
    .RESET_B(_067_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _764_ (.CLK(clknet_3_4__leaf_clk),
    .D(_168_),
    .RESET_B(_068_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _765_ (.CLK(clknet_3_6__leaf_clk),
    .D(_169_),
    .RESET_B(_069_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _766_ (.CLK(clknet_3_7__leaf_clk),
    .D(_170_),
    .RESET_B(_070_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _767_ (.CLK(clknet_3_4__leaf_clk),
    .D(_171_),
    .RESET_B(_071_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _768_ (.CLK(clknet_3_6__leaf_clk),
    .D(_172_),
    .RESET_B(_072_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _769_ (.CLK(clknet_3_4__leaf_clk),
    .D(_173_),
    .RESET_B(_073_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_4 _770_ (.CLK(clknet_3_6__leaf_clk),
    .D(_174_),
    .RESET_B(_074_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_4 _771_ (.CLK(clknet_3_4__leaf_clk),
    .D(_175_),
    .RESET_B(_075_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_4 _772_ (.CLK(clknet_3_7__leaf_clk),
    .D(_176_),
    .RESET_B(_076_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _773_ (.CLK(clknet_3_7__leaf_clk),
    .D(_177_),
    .RESET_B(_077_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_4 _774_ (.CLK(clknet_3_5__leaf_clk),
    .D(_178_),
    .RESET_B(_078_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _775_ (.CLK(clknet_3_6__leaf_clk),
    .D(_179_),
    .RESET_B(_079_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _776_ (.CLK(clknet_3_0__leaf_clk),
    .D(_180_),
    .RESET_B(_080_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _777_ (.CLK(clknet_3_3__leaf_clk),
    .D(_181_),
    .RESET_B(_081_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _778_ (.CLK(clknet_3_0__leaf_clk),
    .D(_182_),
    .RESET_B(_082_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _779_ (.CLK(clknet_3_0__leaf_clk),
    .D(_183_),
    .RESET_B(_083_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _780_ (.CLK(clknet_3_1__leaf_clk),
    .D(_184_),
    .RESET_B(_084_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _781_ (.CLK(clknet_3_1__leaf_clk),
    .D(_185_),
    .RESET_B(_085_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _782_ (.CLK(clknet_3_0__leaf_clk),
    .D(_186_),
    .RESET_B(_086_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _783_ (.CLK(clknet_3_1__leaf_clk),
    .D(_187_),
    .RESET_B(_087_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _784_ (.CLK(clknet_3_1__leaf_clk),
    .D(_188_),
    .RESET_B(_088_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _785_ (.CLK(clknet_3_3__leaf_clk),
    .D(_189_),
    .RESET_B(_089_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net5));
 sky130_fd_sc_hd__dfrtp_1 _786_ (.CLK(clknet_3_2__leaf_clk),
    .D(_190_),
    .RESET_B(_090_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net6));
 sky130_fd_sc_hd__dfrtp_1 _787_ (.CLK(clknet_3_1__leaf_clk),
    .D(_191_),
    .RESET_B(_091_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _788_ (.CLK(clknet_3_3__leaf_clk),
    .D(_192_),
    .RESET_B(_092_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net8));
 sky130_fd_sc_hd__dfrtp_1 _789_ (.CLK(clknet_3_0__leaf_clk),
    .D(_193_),
    .RESET_B(_093_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net9));
 sky130_fd_sc_hd__dfrtp_1 _790_ (.CLK(clknet_3_3__leaf_clk),
    .D(_194_),
    .RESET_B(_094_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net10));
 sky130_fd_sc_hd__dfrtp_1 _791_ (.CLK(clknet_3_0__leaf_clk),
    .D(_195_),
    .RESET_B(_095_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_1 _792_ (.CLK(clknet_3_3__leaf_clk),
    .D(_196_),
    .RESET_B(_096_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _793_ (.CLK(clknet_3_1__leaf_clk),
    .D(_197_),
    .RESET_B(_097_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _794_ (.CLK(clknet_3_1__leaf_clk),
    .D(_198_),
    .RESET_B(_098_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _795_ (.CLK(clknet_3_1__leaf_clk),
    .D(_199_),
    .RESET_B(_099_),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .Q(net16));
 sky130_fd_sc_hd__buf_6 _796_ (.A(net102),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(data_in),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(ena),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(rst),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[15]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net100),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[97]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net101),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[98]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net102),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[99]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net103),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[9]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net104),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(data_out));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[16]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net12),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[17]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[18]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[19]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[1]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[20]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[21]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[22]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[23]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[24]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[25]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[26]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[27]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[28]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[29]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[2]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[30]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[31]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[32]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[33]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[34]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[35]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[36]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[37]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[38]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[39]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[3]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[40]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[41]));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net4),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[0]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[42]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net41),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[43]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[44]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net43),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[45]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[46]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[47]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[48]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net47),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[49]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[4]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[50]));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net5),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[10]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[51]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[52]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[53]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[54]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[55]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[56]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[57]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[58]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[59]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[5]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net6),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[11]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[60]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[61]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[62]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[63]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[64]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[65]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[66]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[67]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[68]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[69]));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net7),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[12]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[6]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[70]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[71]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[72]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[73]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[74]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[75]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[76]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[77]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[78]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net8),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[13]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[79]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[7]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[80]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[81]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[82]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[83]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[84]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[85]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[86]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[87]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net9),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[14]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[88]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[89]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[8]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[90]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[91]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[92]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[93]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[94]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[95]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .VGND(GND),
    .VNB(GND),
    .VPB(VDD),
    .VPWR(VDD),
    .X(ROW_SEL[96]));
endmodule
