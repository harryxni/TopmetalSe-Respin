magic
tech sky130A
timestamp 1758079492
<< metal5 >>
rect 20600 40800 22300 41300
rect 31000 41100 31639 41600
rect 32200 41100 33100 41300
rect 29000 40800 29400 41100
rect 20600 40500 21000 40800
rect 20600 40000 20900 40500
rect 21200 37700 21700 40800
rect 21860 40500 22300 40800
rect 22000 40300 22300 40500
rect 22100 40000 22300 40300
rect 22800 40000 23200 40300
rect 24500 40000 24700 40300
rect 26000 40000 26300 40300
rect 26800 40000 27100 40300
rect 28100 40000 28300 40300
rect 28900 40020 29400 40800
rect 28860 40000 29400 40020
rect 30200 40000 30600 40300
rect 22600 39820 23400 40000
rect 22600 39800 23500 39820
rect 22400 39660 23500 39800
rect 23660 39800 25000 40000
rect 25200 39800 27200 40000
rect 27800 39820 28643 40000
rect 28860 39860 29740 40000
rect 27800 39800 28640 39820
rect 23660 39660 25040 39800
rect 22400 39500 23440 39660
rect 23760 39500 25040 39660
rect 25200 39500 27400 39800
rect 27700 39660 28640 39800
rect 27700 39587 28643 39660
rect 27700 39500 28691 39587
rect 28862 39500 29740 39860
rect 29900 39500 30800 40000
rect 22300 39200 22800 39500
rect 22300 37900 22700 39200
rect 23200 39000 23600 39500
rect 23300 38200 23600 39000
rect 22300 37700 22800 37900
rect 23200 37700 23600 38200
rect 23900 39200 24400 39500
rect 24600 39340 25040 39500
rect 24600 39200 25100 39340
rect 25400 39200 25900 39500
rect 26200 39200 26600 39500
rect 23900 37700 24200 39200
rect 24700 37900 25200 39200
rect 24700 37700 25100 37900
rect 25400 37700 25800 39200
rect 26200 37700 26500 39200
rect 26900 39000 27400 39500
rect 27000 37700 27400 39000
rect 27600 39200 28100 39500
rect 28300 39200 28691 39500
rect 27600 39000 28000 39200
rect 28400 39000 28691 39200
rect 27600 38400 28691 39000
rect 27600 38200 28000 38400
rect 28524 38200 28691 38202
rect 27600 37860 28100 38200
rect 28524 37900 28693 38200
rect 27660 37700 28100 37860
rect 28400 37700 28693 37900
rect 28900 37700 29400 39500
rect 29900 39000 30200 39500
rect 30500 39000 30800 39500
rect 30360 38840 30800 39000
rect 30200 38700 30800 38840
rect 29900 38400 30800 38700
rect 29800 38200 30400 38400
rect 29800 37700 30200 38200
rect 30560 38040 30800 38400
rect 30500 37700 30800 38040
rect 31200 38815 31639 41100
rect 32000 40800 33100 41100
rect 31900 40500 32400 40800
rect 32600 40500 33100 40800
rect 31900 40000 32300 40500
rect 32800 40300 33100 40500
rect 31900 39800 32500 40000
rect 32900 39800 33100 40300
rect 33800 40000 34100 40300
rect 33500 39800 34300 40000
rect 31900 39640 32740 39800
rect 31900 39500 32800 39640
rect 33500 39500 34400 39800
rect 32000 39200 33000 39500
rect 33400 39200 33800 39500
rect 32200 39000 33100 39200
rect 33400 39000 33700 39200
rect 34100 39000 34600 39500
rect 31200 37700 31640 38815
rect 32400 38700 34600 39000
rect 31800 38200 32200 38700
rect 32600 38400 34600 38700
rect 32800 38200 33700 38400
rect 31800 37700 32300 38200
rect 32900 37900 33200 38200
rect 32800 37700 33200 37900
rect 33400 37900 33700 38200
rect 34300 37900 34600 38200
rect 33400 37700 33800 37900
rect 34200 37700 34600 37900
rect 21000 37100 22000 37700
rect 22400 37400 22900 37700
rect 23060 37400 23500 37700
rect 23900 37400 24440 37700
rect 24600 37560 25100 37700
rect 24600 37400 25040 37560
rect 25300 37400 25900 37700
rect 26060 37400 26600 37700
rect 26900 37400 27500 37700
rect 27700 37560 28693 37700
rect 22600 37100 23400 37400
rect 23900 37100 25000 37400
rect 25200 37100 27600 37400
rect 27760 37100 28693 37560
rect 29000 37400 32500 37700
rect 32660 37400 33100 37700
rect 33400 37400 34600 37700
rect 29000 37100 29740 37400
rect 29900 37100 31740 37400
rect 31900 37100 33100 37400
rect 33500 37100 34400 37400
rect 22700 36900 23200 37100
rect 23900 36900 24700 37100
rect 28100 36900 28400 37100
rect 29200 36900 29600 37100
rect 30000 36900 30400 37100
rect 30700 36900 31000 37100
rect 31900 36900 32060 37100
rect 32300 36900 32900 37100
rect 33700 36900 34200 37100
rect 23900 36400 24200 36900
rect 23600 35800 24500 36400
rect 23500 34300 24800 34500
rect 23500 34000 25100 34300
rect 23800 32700 24200 34000
rect 24500 33800 25100 34000
rect 24600 33500 25100 33800
rect 29400 33567 29900 33873
rect 24600 33200 25200 33500
rect 25900 33200 26200 33500
rect 27000 33200 27400 33500
rect 28600 33200 28800 33500
rect 30800 33200 31200 33500
rect 24600 32700 25100 33200
rect 25700 33000 26500 33200
rect 25600 32700 26500 33000
rect 26800 32701 27559 33200
rect 27888 33000 29000 33200
rect 26800 32700 27405 32701
rect 27888 32700 29140 33000
rect 29300 32700 29900 33200
rect 30100 33000 31300 33200
rect 30100 32700 31400 33000
rect 23800 32400 25000 32700
rect 25400 32400 25900 32700
rect 26200 32400 26501 32700
rect 23800 31900 24800 32400
rect 25400 32200 25800 32400
rect 26300 32200 26501 32400
rect 26690 32400 27000 32700
rect 28000 32400 28400 32700
rect 28700 32540 29140 32700
rect 28700 32400 29200 32540
rect 26690 32200 27200 32400
rect 25400 31992 26501 32200
rect 26800 32040 27340 32200
rect 23800 30900 24200 31900
rect 24400 31700 25000 31900
rect 25400 31700 26508 31992
rect 26800 31900 27500 32040
rect 26800 31700 27700 31900
rect 24500 31400 25100 31700
rect 24600 31100 25100 31400
rect 25400 31400 25800 31700
rect 27000 31400 27700 31700
rect 24600 31060 25101 31100
rect 24660 30900 25101 31060
rect 25400 30900 25900 31400
rect 26742 31100 26902 31159
rect 27200 31100 27700 31400
rect 26300 30900 26472 31087
rect 23600 30600 24500 30900
rect 24700 30600 25101 30900
rect 25600 30600 26472 30900
rect 23500 30400 24500 30600
rect 24800 30400 25101 30600
rect 25591 30400 26472 30600
rect 26742 30900 27000 31100
rect 27400 30900 27700 31100
rect 26742 30600 27700 30900
rect 28000 30900 28300 32400
rect 28800 31100 29300 32400
rect 28800 30900 29200 31100
rect 29500 30900 29900 32700
rect 30200 32400 30700 32700
rect 31000 32400 31400 32700
rect 30200 30900 30600 32400
rect 31100 30900 31400 32400
rect 28000 30600 28540 30900
rect 28700 30760 29200 30900
rect 28700 30600 29140 30760
rect 29400 30600 30000 30900
rect 30160 30600 30800 30900
rect 31000 30600 31600 30900
rect 26742 30549 27600 30600
rect 26923 30400 27600 30549
rect 28000 30400 29000 30600
rect 29300 30400 31700 30600
rect 25900 30100 26300 30400
rect 27000 30100 27500 30400
rect 28000 30100 28800 30400
rect 28000 29600 28300 30100
rect 27700 29100 28600 29600
rect 27200 27800 27600 28000
rect 17400 27200 18400 27800
rect 18600 27200 19400 27800
rect 25000 27500 25700 27800
rect 25000 27200 25800 27500
rect 26200 27200 26988 27800
rect 27155 27200 27600 27800
rect 28900 27500 30100 27800
rect 30600 27500 31800 27800
rect 28800 27200 30100 27500
rect 30500 27200 31800 27500
rect 17600 25900 18100 27200
rect 18700 27000 19300 27200
rect 25100 27000 25800 27200
rect 26400 27000 26900 27200
rect 27200 27000 27600 27200
rect 28700 27000 29200 27200
rect 29500 27000 30100 27200
rect 30400 27000 31000 27200
rect 31300 27000 31800 27200
rect 18800 25900 19200 27000
rect 25200 26700 25900 27000
rect 20000 26400 20400 26700
rect 19800 26200 20600 26400
rect 17600 25400 19200 25900
rect 19700 25900 20600 26200
rect 20900 26399 21549 26400
rect 23396 26399 23600 26400
rect 20900 25900 22015 26399
rect 22191 25902 22995 26399
rect 22191 25900 22996 25902
rect 19700 25400 20000 25900
rect 20300 25740 20740 25900
rect 20300 25400 20800 25740
rect 17600 24100 18100 25400
rect 18800 24400 19200 25400
rect 20160 25240 20800 25400
rect 20000 25100 20800 25240
rect 19800 24900 20800 25100
rect 19700 24600 20200 24900
rect 18800 24100 19300 24400
rect 19600 24100 20000 24600
rect 20360 24440 20800 24900
rect 20300 24100 20800 24440
rect 21100 25700 22000 25900
rect 21100 24100 21500 25700
rect 21700 25400 22000 25700
rect 22200 25854 22996 25900
rect 22200 25700 23000 25854
rect 22200 24100 22600 25700
rect 22800 25400 23000 25700
rect 23200 25400 23600 26399
rect 23900 25900 24500 26400
rect 25300 26200 26000 26700
rect 25300 25900 26200 26200
rect 24000 25700 24200 25900
rect 23300 25100 23600 25400
rect 23900 25400 24200 25700
rect 23900 25100 24100 25400
rect 23300 24600 24100 25100
rect 23400 24100 24000 24600
rect 25300 24400 25600 25900
rect 25760 25700 26300 25900
rect 26500 25860 26800 27000
rect 28600 26400 29000 27000
rect 29600 26700 30100 27000
rect 27000 25900 27600 26400
rect 25800 25400 26400 25700
rect 25900 25100 26400 25400
rect 26560 25100 26800 25860
rect 25900 24900 26800 25100
rect 26000 24600 26800 24900
rect 26200 24400 26800 24600
rect 25200 24100 25600 24400
rect 17500 23800 18400 24100
rect 17400 23600 18400 23800
rect 18600 23600 19400 24100
rect 19600 23800 20840 24100
rect 21000 23800 21600 24100
rect 22100 23800 22700 24100
rect 19700 23600 21700 23800
rect 22000 23600 22800 23800
rect 23500 23600 23900 24100
rect 25000 23600 25900 24100
rect 26300 23800 26800 24400
rect 27200 24100 27600 25900
rect 28400 24900 28900 26400
rect 29800 26200 30100 26700
rect 30260 26400 30700 27000
rect 31400 26560 31800 27000
rect 32400 26700 32600 27000
rect 35400 26700 35600 27000
rect 36800 26700 37200 27000
rect 30260 26200 30600 26400
rect 31400 26200 31740 26560
rect 32000 26400 33000 26700
rect 29900 25900 30600 26200
rect 31579 26073 31740 26200
rect 31900 26200 33100 26400
rect 30100 25100 30600 25900
rect 31900 25400 32300 26200
rect 32600 25100 33100 26200
rect 33500 25900 34600 26700
rect 35000 26400 36000 26700
rect 36600 26400 37400 26700
rect 34900 26200 36100 26400
rect 36500 26200 37600 26400
rect 33500 25400 33700 25900
rect 34800 25700 35300 26200
rect 35600 25900 36100 26200
rect 33500 25100 34200 25400
rect 34800 25220 35200 25700
rect 30200 25060 30600 25100
rect 30260 24900 30600 25060
rect 32500 24900 33000 25100
rect 33400 24900 34400 25100
rect 34700 25060 35200 25220
rect 34760 24900 35200 25060
rect 28400 24600 29000 24900
rect 29900 24600 30100 24900
rect 28600 24400 29000 24600
rect 29800 24400 30100 24600
rect 30260 24400 30700 24900
rect 31600 24560 31800 24900
rect 32300 24600 32900 24900
rect 33400 24600 34600 24900
rect 31580 24400 31760 24560
rect 32000 24400 32600 24600
rect 33400 24400 33700 24600
rect 34100 24400 34600 24600
rect 28600 24100 29200 24400
rect 29600 24100 30100 24400
rect 30400 24100 31000 24400
rect 31400 24100 31740 24400
rect 31920 24241 33200 24400
rect 27100 23800 27700 24100
rect 28700 23800 30000 24100
rect 30400 23800 31700 24100
rect 31900 23800 33200 24241
rect 34200 24100 34600 24400
rect 34800 24600 35200 24900
rect 34800 24100 35300 24600
rect 35800 24400 36200 25900
rect 36400 25700 36800 26200
rect 37200 25700 37700 26200
rect 36400 25100 36700 25700
rect 36400 24600 36800 25100
rect 37300 24900 37700 25700
rect 37200 24600 37700 24900
rect 35800 24100 36100 24400
rect 36500 24100 37700 24600
rect 34200 23800 34634 24100
rect 34900 23800 35400 24100
rect 35600 23800 36100 24100
rect 36700 24098 37100 24100
rect 36700 23800 36941 24098
rect 37260 23938 37700 24100
rect 37200 23800 37700 23938
rect 26400 23600 26800 23800
rect 27000 23600 27800 23800
rect 28800 23600 29900 23800
rect 30500 23600 31600 23800
rect 31900 23600 33700 23800
rect 34200 23600 34600 23800
rect 35000 23600 36000 23800
rect 37110 23776 37600 23800
rect 37100 23600 37600 23776
rect 19800 23300 20200 23600
rect 20500 23300 20900 23600
rect 23500 23300 23800 23600
rect 26500 23300 26800 23600
rect 29000 23300 29600 23600
rect 30800 23300 31300 23600
rect 23400 23100 23800 23300
rect 33200 23100 33700 23600
rect 34100 23100 34600 23600
rect 35200 23300 35800 23600
rect 37000 23300 37600 23600
rect 36800 23100 37400 23300
rect 22900 22500 23600 23100
rect 33400 22800 34400 23100
rect 36600 22800 37300 23100
rect 33500 22500 34300 22800
rect 36600 22500 37100 22800
rect 23000 22300 23500 22500
<< properties >>
<< end >>
