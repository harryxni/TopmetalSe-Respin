magic
tech sky130A
timestamp 1757709129
<< viali >>
rect 796 6740 813 6757
rect 2314 6740 2331 6757
rect 3832 6740 3849 6757
rect 5396 6740 5413 6757
rect 7052 6740 7069 6757
rect 8432 6740 8449 6757
rect 9996 6740 10013 6757
rect 11514 6740 11531 6757
rect 12848 6740 12865 6757
rect 14504 6740 14521 6757
rect 15792 6740 15809 6757
rect 23796 6740 23813 6757
rect 25176 6740 25193 6757
rect 25498 6740 25515 6757
rect 71452 6740 71469 6757
rect 72372 6740 72389 6757
rect 74160 6740 74177 6757
rect 78812 6740 78829 6757
rect 91370 6740 91387 6757
rect 92888 6740 92905 6757
rect 105170 6740 105187 6757
rect 106688 6740 106705 6757
rect 134696 6740 134713 6757
rect 137140 6740 137157 6757
rect 137462 6740 137479 6757
rect 138934 6740 138951 6757
rect 140452 6740 140469 6757
rect 142292 6740 142309 6757
rect 143580 6740 143597 6757
rect 145052 6740 145069 6757
rect 146616 6740 146633 6757
rect 148134 6740 148151 6757
rect 149652 6740 149669 6757
rect 150710 6740 150727 6757
rect 150894 6740 150911 6757
rect 151078 6740 151095 6757
rect 151492 6740 151509 6757
rect 151676 6740 151693 6757
rect 22140 6706 22157 6723
rect 30236 6706 30253 6723
rect 31524 6706 31541 6723
rect 37688 6706 37705 6723
rect 46980 6706 46997 6723
rect 50568 6706 50585 6723
rect 54708 6706 54725 6723
rect 55628 6706 55645 6723
rect 60642 6706 60659 6723
rect 62068 6706 62085 6723
rect 68324 6706 68341 6723
rect 70164 6706 70181 6723
rect 77892 6706 77909 6723
rect 85206 6706 85223 6723
rect 86540 6706 86557 6723
rect 86908 6706 86925 6723
rect 87920 6706 87937 6723
rect 89070 6706 89087 6723
rect 90772 6706 90789 6723
rect 99926 6706 99943 6723
rect 101950 6706 101967 6723
rect 108206 6706 108223 6723
rect 110092 6706 110109 6723
rect 113312 6706 113329 6723
rect 114830 6706 114847 6723
rect 119982 6706 119999 6723
rect 123570 6706 123587 6723
rect 124766 6706 124783 6723
rect 126422 6706 126439 6723
rect 127710 6706 127727 6723
rect 129734 6706 129751 6723
rect 131344 6706 131361 6723
rect 133000 6706 133017 6723
rect 13170 6672 13187 6689
rect 13630 6672 13647 6689
rect 17356 6672 17373 6689
rect 18782 6672 18799 6689
rect 22784 6672 22801 6689
rect 25820 6672 25837 6689
rect 36354 6672 36371 6689
rect 36814 6672 36831 6689
rect 39252 6672 39269 6689
rect 40126 6672 40143 6689
rect 40770 6672 40787 6689
rect 40816 6672 40833 6689
rect 49004 6672 49021 6689
rect 49096 6672 49113 6689
rect 56134 6672 56151 6689
rect 60136 6672 60153 6689
rect 62850 6672 62867 6689
rect 63356 6672 63373 6689
rect 65150 6672 65167 6689
rect 66300 6672 66317 6689
rect 74028 6672 74045 6689
rect 75454 6672 75471 6689
rect 76742 6672 76759 6689
rect 80468 6672 80485 6689
rect 83320 6672 83337 6689
rect 83780 6672 83797 6689
rect 87138 6672 87155 6689
rect 87184 6672 87201 6689
rect 89484 6672 89501 6689
rect 91048 6672 91065 6689
rect 94268 6672 94285 6689
rect 94912 6672 94929 6689
rect 99374 6672 99391 6689
rect 100570 6672 100587 6689
rect 102364 6672 102381 6689
rect 103928 6672 103945 6689
rect 112162 6672 112179 6689
rect 113542 6672 113559 6689
rect 113588 6672 113605 6689
rect 115244 6672 115261 6689
rect 116118 6672 116135 6689
rect 118602 6672 118619 6689
rect 118648 6672 118665 6689
rect 120396 6672 120413 6689
rect 121684 6672 121701 6689
rect 122558 6672 122575 6689
rect 125088 6672 125105 6689
rect 131022 6672 131039 6689
rect 131620 6672 131637 6689
rect 133276 6672 133293 6689
rect 134564 6672 134581 6689
rect 135852 6672 135869 6689
rect 152228 6672 152245 6689
rect 152458 6672 152475 6689
rect 152688 6672 152705 6689
rect 888 6638 905 6655
rect 2406 6638 2423 6655
rect 3924 6638 3941 6655
rect 5488 6638 5505 6655
rect 7144 6638 7161 6655
rect 8524 6638 8541 6655
rect 10088 6638 10105 6655
rect 11606 6638 11623 6655
rect 13032 6638 13049 6655
rect 14918 6638 14935 6655
rect 16206 6638 16223 6655
rect 20070 6638 20087 6655
rect 21266 6638 21283 6655
rect 23888 6638 23905 6655
rect 25268 6638 25285 6655
rect 25682 6638 25699 6655
rect 26510 6638 26527 6655
rect 27798 6638 27815 6655
rect 28948 6638 28965 6655
rect 30328 6638 30345 6655
rect 31616 6638 31633 6655
rect 33088 6638 33105 6655
rect 34652 6638 34669 6655
rect 36262 6638 36279 6655
rect 38102 6638 38119 6655
rect 41230 6638 41247 6655
rect 41552 6638 41569 6655
rect 41966 6638 41983 6655
rect 43254 6638 43271 6655
rect 44404 6638 44421 6655
rect 47072 6638 47089 6655
rect 48452 6638 48469 6655
rect 49694 6638 49711 6655
rect 50982 6638 50999 6655
rect 52132 6638 52149 6655
rect 54800 6638 54817 6655
rect 55720 6638 55737 6655
rect 57422 6638 57439 6655
rect 58710 6638 58727 6655
rect 60090 6638 60107 6655
rect 60734 6638 60751 6655
rect 62160 6638 62177 6655
rect 63310 6638 63327 6655
rect 63770 6638 63787 6655
rect 68416 6638 68433 6655
rect 70256 6638 70273 6655
rect 71544 6638 71561 6655
rect 72464 6638 72481 6655
rect 72878 6638 72895 6655
rect 77984 6638 78001 6655
rect 78214 6638 78231 6655
rect 78904 6638 78921 6655
rect 79318 6638 79335 6655
rect 81756 6638 81773 6655
rect 85298 6638 85315 6655
rect 86632 6638 86649 6655
rect 87092 6638 87109 6655
rect 87828 6638 87845 6655
rect 88196 6638 88213 6655
rect 91002 6638 91019 6655
rect 91462 6638 91479 6655
rect 92980 6638 92997 6655
rect 93670 6638 93687 6655
rect 94222 6638 94239 6655
rect 94774 6638 94791 6655
rect 95924 6638 95941 6655
rect 97212 6638 97229 6655
rect 100018 6638 100035 6655
rect 101076 6638 101093 6655
rect 103836 6638 103853 6655
rect 105262 6638 105279 6655
rect 106780 6638 106797 6655
rect 108298 6638 108315 6655
rect 110184 6638 110201 6655
rect 111472 6638 111489 6655
rect 112944 6638 112961 6655
rect 113956 6638 113973 6655
rect 116532 6638 116549 6655
rect 116946 6638 116963 6655
rect 117544 6638 117561 6655
rect 118556 6638 118573 6655
rect 119108 6638 119125 6655
rect 123662 6638 123679 6655
rect 124996 6638 125013 6655
rect 125548 6638 125565 6655
rect 126836 6638 126853 6655
rect 128124 6638 128141 6655
rect 129826 6638 129843 6655
rect 132126 6638 132143 6655
rect 134288 6638 134305 6655
rect 137232 6638 137249 6655
rect 137554 6638 137571 6655
rect 139026 6638 139043 6655
rect 140544 6638 140561 6655
rect 142384 6638 142401 6655
rect 143672 6638 143689 6655
rect 145144 6638 145161 6655
rect 146708 6638 146725 6655
rect 148226 6638 148243 6655
rect 149744 6638 149761 6655
rect 151860 6638 151877 6655
rect 13768 6604 13785 6621
rect 15056 6604 15073 6621
rect 16344 6604 16361 6621
rect 17494 6604 17511 6621
rect 18920 6604 18937 6621
rect 20208 6604 20225 6621
rect 21404 6604 21421 6621
rect 22738 6604 22755 6621
rect 26648 6604 26665 6621
rect 27936 6604 27953 6621
rect 29086 6604 29103 6621
rect 36952 6604 36969 6621
rect 38240 6604 38257 6621
rect 39390 6604 39407 6621
rect 42104 6604 42121 6621
rect 43392 6604 43409 6621
rect 44542 6604 44559 6621
rect 45922 6604 45939 6621
rect 46014 6604 46031 6621
rect 49832 6604 49849 6621
rect 51120 6604 51137 6621
rect 52270 6604 52287 6621
rect 56272 6604 56289 6621
rect 57560 6604 57577 6621
rect 58848 6604 58865 6621
rect 60044 6604 60061 6621
rect 62758 6604 62775 6621
rect 63908 6604 63925 6621
rect 65288 6604 65305 6621
rect 66438 6604 66455 6621
rect 73016 6604 73033 6621
rect 75040 6604 75057 6621
rect 75592 6604 75609 6621
rect 76880 6604 76897 6621
rect 78260 6604 78277 6621
rect 79456 6604 79473 6621
rect 80606 6604 80623 6621
rect 81894 6604 81911 6621
rect 83274 6604 83291 6621
rect 83688 6604 83705 6621
rect 88334 6604 88351 6621
rect 89622 6604 89639 6621
rect 90956 6604 90973 6621
rect 93716 6604 93733 6621
rect 96062 6604 96079 6621
rect 96936 6604 96953 6621
rect 97350 6604 97367 6621
rect 98224 6604 98241 6621
rect 98914 6604 98931 6621
rect 99328 6604 99345 6621
rect 101214 6604 101231 6621
rect 102502 6604 102519 6621
rect 114094 6604 114111 6621
rect 115382 6604 115399 6621
rect 119246 6604 119263 6621
rect 120534 6604 120551 6621
rect 121822 6604 121839 6621
rect 125686 6604 125703 6621
rect 126974 6604 126991 6621
rect 128262 6604 128279 6621
rect 130930 6604 130947 6621
rect 131528 6604 131545 6621
rect 132264 6604 132281 6621
rect 133414 6604 133431 6621
rect 135990 6604 136007 6621
rect 13078 6570 13095 6587
rect 17080 6570 17097 6587
rect 18230 6570 18247 6587
rect 19656 6570 19673 6587
rect 20944 6570 20961 6587
rect 22508 6570 22525 6587
rect 22692 6570 22709 6587
rect 25728 6570 25745 6587
rect 27384 6570 27401 6587
rect 28672 6570 28689 6587
rect 29822 6570 29839 6587
rect 32996 6570 33013 6587
rect 34560 6570 34577 6587
rect 36032 6570 36049 6587
rect 36216 6570 36233 6587
rect 38976 6570 38993 6587
rect 40540 6570 40557 6587
rect 40724 6570 40741 6587
rect 41138 6570 41155 6587
rect 41460 6570 41477 6587
rect 42840 6570 42857 6587
rect 44128 6570 44145 6587
rect 45278 6570 45295 6587
rect 48360 6570 48377 6587
rect 48774 6570 48791 6587
rect 48958 6570 48975 6587
rect 51856 6570 51873 6587
rect 53006 6570 53023 6587
rect 57008 6570 57025 6587
rect 58296 6570 58313 6587
rect 59584 6570 59601 6587
rect 59860 6570 59877 6587
rect 63080 6570 63097 6587
rect 63264 6570 63281 6587
rect 64644 6570 64661 6587
rect 66024 6570 66041 6587
rect 67174 6570 67191 6587
rect 73752 6570 73769 6587
rect 76328 6570 76345 6587
rect 77616 6570 77633 6587
rect 80192 6570 80209 6587
rect 81342 6570 81359 6587
rect 82630 6570 82647 6587
rect 83044 6570 83061 6587
rect 83228 6570 83245 6587
rect 90358 6570 90375 6587
rect 93992 6570 94009 6587
rect 94176 6570 94193 6587
rect 95648 6570 95665 6587
rect 99098 6570 99115 6587
rect 99282 6570 99299 6587
rect 100248 6570 100265 6587
rect 100432 6570 100449 6587
rect 100478 6570 100495 6587
rect 103238 6570 103255 6587
rect 103652 6570 103669 6587
rect 103882 6570 103899 6587
rect 111380 6570 111397 6587
rect 111840 6570 111857 6587
rect 112024 6570 112041 6587
rect 112070 6570 112087 6587
rect 112852 6570 112869 6587
rect 113496 6570 113513 6587
rect 116578 6570 116595 6587
rect 116854 6570 116871 6587
rect 117452 6570 117469 6587
rect 118372 6570 118389 6587
rect 121270 6570 121287 6587
rect 124950 6570 124967 6587
rect 128998 6570 129015 6587
rect 131574 6570 131591 6587
rect 135438 6570 135455 6587
rect 136726 6570 136743 6587
rect 147950 6570 147967 6587
rect 13032 6468 13049 6485
rect 13722 6468 13739 6485
rect 16942 6468 16959 6485
rect 17402 6468 17419 6485
rect 17770 6468 17787 6485
rect 18322 6468 18339 6485
rect 21266 6468 21283 6485
rect 21726 6468 21743 6485
rect 22278 6468 22295 6485
rect 26004 6468 26021 6485
rect 26786 6468 26803 6485
rect 26970 6468 26987 6485
rect 29270 6468 29287 6485
rect 36078 6468 36095 6485
rect 44772 6468 44789 6485
rect 45554 6468 45571 6485
rect 56134 6468 56151 6485
rect 59124 6468 59141 6485
rect 59354 6468 59371 6485
rect 63356 6468 63373 6485
rect 64046 6468 64063 6485
rect 64368 6468 64385 6485
rect 64598 6468 64615 6485
rect 65150 6468 65167 6485
rect 66760 6468 66777 6485
rect 67174 6468 67191 6485
rect 72740 6468 72757 6485
rect 75730 6468 75747 6485
rect 76374 6468 76391 6485
rect 76558 6468 76575 6485
rect 76742 6468 76759 6485
rect 76926 6468 76943 6485
rect 77110 6468 77127 6485
rect 77478 6468 77495 6485
rect 78030 6468 78047 6485
rect 78214 6468 78231 6485
rect 78398 6468 78415 6485
rect 78582 6468 78599 6485
rect 81802 6468 81819 6485
rect 82216 6468 82233 6485
rect 83918 6468 83935 6485
rect 87506 6468 87523 6485
rect 87828 6468 87845 6485
rect 90404 6468 90421 6485
rect 96154 6468 96171 6485
rect 97994 6468 98011 6485
rect 103284 6468 103301 6485
rect 126192 6468 126209 6485
rect 132310 6468 132327 6485
rect 151308 6468 151325 6485
rect 152228 6468 152245 6485
rect 14504 6434 14521 6451
rect 18276 6434 18293 6451
rect 18690 6434 18707 6451
rect 19242 6434 19259 6451
rect 19886 6434 19903 6451
rect 29316 6434 29333 6451
rect 38930 6434 38947 6451
rect 39298 6434 39315 6451
rect 49740 6434 49757 6451
rect 52316 6434 52333 6451
rect 52362 6434 52379 6451
rect 56180 6434 56197 6451
rect 57008 6434 57025 6451
rect 57836 6434 57853 6451
rect 66806 6434 66823 6451
rect 72970 6434 72987 6451
rect 79640 6434 79657 6451
rect 82262 6434 82279 6451
rect 90818 6434 90835 6451
rect 94774 6434 94791 6451
rect 95464 6434 95481 6451
rect 96660 6434 96677 6451
rect 97948 6434 97965 6451
rect 115520 6434 115537 6451
rect 119384 6434 119401 6451
rect 120488 6434 120505 6451
rect 122650 6434 122667 6451
rect 125686 6434 125703 6451
rect 126238 6434 126255 6451
rect 130884 6434 130901 6451
rect 131620 6434 131637 6451
rect 131712 6434 131729 6451
rect 132770 6434 132787 6451
rect 135898 6434 135915 6451
rect 136450 6434 136467 6451
rect 152504 6434 152521 6451
rect 152734 6434 152751 6451
rect 13124 6400 13141 6417
rect 13906 6400 13923 6417
rect 17356 6400 17373 6417
rect 17862 6400 17879 6417
rect 19196 6400 19213 6417
rect 20852 6400 20869 6417
rect 21220 6400 21237 6417
rect 22370 6400 22387 6417
rect 26096 6400 26113 6417
rect 26464 6400 26481 6417
rect 27016 6400 27033 6417
rect 27384 6400 27401 6417
rect 28534 6400 28551 6417
rect 36170 6400 36187 6417
rect 37550 6400 37567 6417
rect 37780 6400 37797 6417
rect 38884 6400 38901 6417
rect 39252 6400 39269 6417
rect 39666 6400 39683 6417
rect 39896 6400 39913 6417
rect 43116 6400 43133 6417
rect 45232 6400 45249 6417
rect 45646 6400 45663 6417
rect 49280 6400 49297 6417
rect 53052 6400 53069 6417
rect 56548 6400 56565 6417
rect 56916 6400 56933 6417
rect 57330 6400 57347 6417
rect 59446 6400 59463 6417
rect 63448 6400 63465 6417
rect 63724 6400 63741 6417
rect 64138 6400 64155 6417
rect 64552 6400 64569 6417
rect 65104 6400 65121 6417
rect 65426 6400 65443 6417
rect 67266 6400 67283 6417
rect 67680 6400 67697 6417
rect 71498 6400 71515 6417
rect 72924 6400 72941 6417
rect 73522 6400 73539 6417
rect 74948 6400 74965 6417
rect 77432 6400 77449 6417
rect 79594 6400 79611 6417
rect 80008 6400 80025 6417
rect 80606 6400 80623 6417
rect 80928 6400 80945 6417
rect 82676 6400 82693 6417
rect 83274 6400 83291 6417
rect 83688 6400 83705 6417
rect 84010 6400 84027 6417
rect 87598 6400 87615 6417
rect 87920 6400 87937 6417
rect 88196 6400 88213 6417
rect 89300 6400 89317 6417
rect 90496 6400 90513 6417
rect 90772 6400 90789 6417
rect 91094 6400 91111 6417
rect 94038 6400 94055 6417
rect 94314 6400 94331 6417
rect 94682 6400 94699 6417
rect 95510 6400 95527 6417
rect 96108 6400 96125 6417
rect 97534 6400 97551 6417
rect 98684 6400 98701 6417
rect 98730 6400 98747 6417
rect 99190 6400 99207 6417
rect 100248 6400 100265 6417
rect 100662 6400 100679 6417
rect 102410 6400 102427 6417
rect 103744 6400 103761 6417
rect 113358 6400 113375 6417
rect 113680 6400 113697 6417
rect 113956 6400 113973 6417
rect 115152 6400 115169 6417
rect 115382 6400 115399 6417
rect 116532 6400 116549 6417
rect 118510 6400 118527 6417
rect 118832 6400 118849 6417
rect 119246 6400 119263 6417
rect 120350 6400 120367 6417
rect 121914 6400 121931 6417
rect 122282 6400 122299 6417
rect 122374 6400 122391 6417
rect 122604 6400 122621 6417
rect 125180 6400 125197 6417
rect 125778 6400 125795 6417
rect 128124 6400 128141 6417
rect 128538 6400 128555 6417
rect 131252 6400 131269 6417
rect 132080 6400 132097 6417
rect 132402 6400 132419 6417
rect 132632 6400 132649 6417
rect 133920 6400 133937 6417
rect 134564 6400 134581 6417
rect 135852 6400 135869 6417
rect 151400 6400 151417 6417
rect 152320 6400 152337 6417
rect 13952 6366 13969 6383
rect 14044 6366 14061 6383
rect 14550 6366 14567 6383
rect 14642 6366 14659 6383
rect 14918 6366 14935 6383
rect 15056 6366 15073 6383
rect 16068 6366 16085 6383
rect 16206 6366 16223 6383
rect 17448 6366 17465 6383
rect 18782 6366 18799 6383
rect 19288 6366 19305 6383
rect 19748 6366 19765 6383
rect 21772 6366 21789 6383
rect 21864 6366 21881 6383
rect 27062 6366 27079 6383
rect 27522 6366 27539 6383
rect 29362 6366 29379 6383
rect 37918 6366 37935 6383
rect 40034 6366 40051 6383
rect 42012 6366 42029 6383
rect 42150 6366 42167 6383
rect 43254 6366 43271 6383
rect 44818 6366 44835 6383
rect 44910 6366 44927 6383
rect 49602 6366 49619 6383
rect 50706 6366 50723 6383
rect 50844 6366 50861 6383
rect 52408 6366 52425 6383
rect 56272 6366 56289 6383
rect 56594 6366 56611 6383
rect 57882 6366 57899 6383
rect 57928 6366 57945 6383
rect 58250 6366 58267 6383
rect 58388 6366 58405 6383
rect 64690 6366 64707 6383
rect 65564 6366 65581 6383
rect 66300 6366 66317 6383
rect 66898 6366 66915 6383
rect 71636 6366 71653 6383
rect 73062 6366 73079 6383
rect 73752 6366 73769 6383
rect 73890 6366 73907 6383
rect 74626 6366 74643 6383
rect 75776 6366 75793 6383
rect 75868 6366 75885 6383
rect 77524 6366 77541 6383
rect 79732 6366 79749 6383
rect 81066 6366 81083 6383
rect 82308 6366 82325 6383
rect 88334 6366 88351 6383
rect 89438 6366 89455 6383
rect 95602 6366 95619 6383
rect 96200 6366 96217 6383
rect 96522 6366 96539 6383
rect 98086 6366 98103 6383
rect 98822 6366 98839 6383
rect 99052 6366 99069 6383
rect 100294 6366 100311 6383
rect 101306 6366 101323 6383
rect 101444 6366 101461 6383
rect 102548 6366 102565 6383
rect 114094 6366 114111 6383
rect 116578 6366 116595 6383
rect 126284 6366 126301 6383
rect 126836 6366 126853 6383
rect 126974 6366 126991 6383
rect 127710 6366 127727 6383
rect 128170 6366 128187 6383
rect 128216 6366 128233 6383
rect 133966 6366 133983 6383
rect 134012 6366 134029 6383
rect 134702 6366 134719 6383
rect 135990 6366 136007 6383
rect 136496 6366 136513 6383
rect 136542 6366 136559 6383
rect 37458 6332 37475 6349
rect 39574 6332 39591 6349
rect 40770 6332 40787 6349
rect 50476 6332 50493 6349
rect 52960 6332 52977 6349
rect 67772 6332 67789 6349
rect 76190 6332 76207 6349
rect 77248 6332 77265 6349
rect 79410 6332 79427 6349
rect 80100 6332 80117 6349
rect 83596 6332 83613 6349
rect 93946 6332 93963 6349
rect 103652 6332 103669 6349
rect 113588 6332 113605 6349
rect 118740 6332 118757 6349
rect 125088 6332 125105 6349
rect 127940 6332 127957 6349
rect 131344 6332 131361 6349
rect 14320 6298 14337 6315
rect 15792 6298 15809 6315
rect 17172 6298 17189 6315
rect 19012 6298 19029 6315
rect 20622 6298 20639 6315
rect 20898 6298 20915 6315
rect 21542 6298 21559 6315
rect 26510 6298 26527 6315
rect 28258 6298 28275 6315
rect 28580 6298 28597 6315
rect 29086 6298 29103 6315
rect 38654 6298 38671 6315
rect 42886 6298 42903 6315
rect 43990 6298 44007 6315
rect 44588 6298 44605 6315
rect 45278 6298 45295 6315
rect 49188 6298 49205 6315
rect 51580 6298 51597 6315
rect 52132 6298 52149 6315
rect 55950 6298 55967 6315
rect 57376 6298 57393 6315
rect 57652 6298 57669 6315
rect 63770 6298 63787 6315
rect 66576 6298 66593 6315
rect 73430 6298 73447 6315
rect 74994 6298 75011 6315
rect 75546 6298 75563 6315
rect 80652 6298 80669 6315
rect 82032 6298 82049 6315
rect 82722 6298 82739 6315
rect 83320 6298 83337 6315
rect 89070 6298 89087 6315
rect 90174 6298 90191 6315
rect 91140 6298 91157 6315
rect 94360 6298 94377 6315
rect 95280 6298 95297 6315
rect 95924 6298 95941 6315
rect 97764 6298 97781 6315
rect 98500 6298 98517 6315
rect 99098 6298 99115 6315
rect 100570 6298 100587 6315
rect 102180 6298 102197 6315
rect 113266 6298 113283 6315
rect 114830 6298 114847 6315
rect 115060 6298 115077 6315
rect 116256 6298 116273 6315
rect 118418 6298 118435 6315
rect 120120 6298 120137 6315
rect 121224 6298 121241 6315
rect 121960 6298 121977 6315
rect 126008 6298 126025 6315
rect 128584 6298 128601 6315
rect 130930 6298 130947 6315
rect 131988 6298 132005 6315
rect 133506 6298 133523 6315
rect 133736 6298 133753 6315
rect 135438 6298 135455 6315
rect 135668 6298 135685 6315
rect 136266 6298 136283 6315
rect 15654 6196 15671 6213
rect 16988 6196 17005 6213
rect 17402 6196 17419 6213
rect 18598 6196 18615 6213
rect 19242 6196 19259 6213
rect 19610 6196 19627 6213
rect 21588 6196 21605 6213
rect 21910 6196 21927 6213
rect 27062 6196 27079 6213
rect 27338 6196 27355 6213
rect 28672 6196 28689 6213
rect 28994 6196 29011 6213
rect 37596 6196 37613 6213
rect 39666 6196 39683 6213
rect 40126 6196 40143 6213
rect 42794 6196 42811 6213
rect 43208 6196 43225 6213
rect 44450 6196 44467 6213
rect 45094 6196 45111 6213
rect 49556 6196 49573 6213
rect 49924 6196 49941 6213
rect 51948 6196 51965 6213
rect 52592 6196 52609 6213
rect 56548 6196 56565 6213
rect 56870 6196 56887 6213
rect 59216 6196 59233 6213
rect 63862 6196 63879 6213
rect 65426 6196 65443 6213
rect 66346 6196 66363 6213
rect 73660 6196 73677 6213
rect 76282 6196 76299 6213
rect 77064 6196 77081 6213
rect 82676 6196 82693 6213
rect 87966 6196 87983 6213
rect 90680 6196 90697 6213
rect 94268 6196 94285 6213
rect 95096 6196 95113 6213
rect 100846 6196 100863 6213
rect 103238 6196 103255 6213
rect 113904 6196 113921 6213
rect 116118 6196 116135 6213
rect 119982 6196 119999 6213
rect 121776 6196 121793 6213
rect 122098 6196 122115 6213
rect 125548 6196 125565 6213
rect 128446 6196 128463 6213
rect 131252 6196 131269 6213
rect 132310 6196 132327 6213
rect 135530 6196 135547 6213
rect 152734 6196 152751 6213
rect 38746 6162 38763 6179
rect 44726 6162 44743 6179
rect 74212 6162 74229 6179
rect 76650 6162 76667 6179
rect 80008 6162 80025 6179
rect 83044 6162 83061 6179
rect 90450 6162 90467 6179
rect 96292 6162 96309 6179
rect 100570 6162 100587 6179
rect 114876 6162 114893 6179
rect 119384 6162 119401 6179
rect 121178 6162 121195 6179
rect 126054 6162 126071 6179
rect 127158 6162 127175 6179
rect 128170 6162 128187 6179
rect 132034 6162 132051 6179
rect 135852 6162 135869 6179
rect 13860 6128 13877 6145
rect 14366 6128 14383 6145
rect 14458 6128 14475 6145
rect 14780 6128 14797 6145
rect 15884 6128 15901 6145
rect 20438 6128 20455 6145
rect 26188 6128 26205 6145
rect 27844 6128 27861 6145
rect 28350 6128 28367 6145
rect 38378 6128 38395 6145
rect 38470 6128 38487 6145
rect 39068 6128 39085 6145
rect 42242 6128 42259 6145
rect 42334 6128 42351 6145
rect 43530 6128 43547 6145
rect 44082 6128 44099 6145
rect 50476 6128 50493 6145
rect 51580 6128 51597 6145
rect 52270 6128 52287 6145
rect 57192 6128 57209 6145
rect 58894 6128 58911 6145
rect 65932 6128 65949 6145
rect 76052 6128 76069 6145
rect 76098 6128 76115 6145
rect 76972 6128 76989 6145
rect 80652 6128 80669 6145
rect 80744 6128 80761 6145
rect 81250 6128 81267 6145
rect 81342 6128 81359 6145
rect 81802 6128 81819 6145
rect 88518 6128 88535 6145
rect 88564 6128 88581 6145
rect 95418 6128 95435 6145
rect 96844 6128 96861 6145
rect 98776 6128 98793 6145
rect 101766 6128 101783 6145
rect 102364 6128 102381 6145
rect 115796 6128 115813 6145
rect 119660 6128 119677 6145
rect 120718 6128 120735 6145
rect 121408 6128 121425 6145
rect 121454 6128 121471 6145
rect 126284 6128 126301 6145
rect 127664 6128 127681 6145
rect 132862 6128 132879 6145
rect 132954 6128 132971 6145
rect 134380 6128 134397 6145
rect 136128 6128 136145 6145
rect 13722 6094 13739 6111
rect 14320 6094 14337 6111
rect 17080 6094 17097 6111
rect 17356 6094 17373 6111
rect 17678 6094 17695 6111
rect 18184 6094 18201 6111
rect 18552 6094 18569 6111
rect 19334 6094 19351 6111
rect 19564 6094 19581 6111
rect 20300 6094 20317 6111
rect 20714 6094 20731 6111
rect 21864 6094 21881 6111
rect 27292 6094 27309 6111
rect 28304 6094 28321 6111
rect 28764 6094 28781 6111
rect 29086 6094 29103 6111
rect 37688 6094 37705 6111
rect 38332 6094 38349 6111
rect 38976 6094 38993 6111
rect 39620 6094 39637 6111
rect 40080 6094 40097 6111
rect 42196 6094 42213 6111
rect 42748 6094 42765 6111
rect 43438 6094 43455 6111
rect 43990 6094 44007 6111
rect 44404 6094 44421 6111
rect 44818 6094 44835 6111
rect 45048 6094 45065 6111
rect 49648 6094 49665 6111
rect 49878 6094 49895 6111
rect 51488 6094 51505 6111
rect 51902 6094 51919 6111
rect 52224 6094 52241 6111
rect 52546 6094 52563 6111
rect 56640 6094 56657 6111
rect 56962 6094 56979 6111
rect 58802 6094 58819 6111
rect 59170 6094 59187 6111
rect 63954 6094 63971 6111
rect 64322 6094 64339 6111
rect 64552 6094 64569 6111
rect 65840 6094 65857 6111
rect 66300 6094 66317 6111
rect 68876 6094 68893 6111
rect 73752 6094 73769 6111
rect 74166 6094 74183 6111
rect 74718 6094 74735 6111
rect 76236 6094 76253 6111
rect 77156 6094 77173 6111
rect 80100 6094 80117 6111
rect 80606 6094 80623 6111
rect 88058 6094 88075 6111
rect 88472 6094 88489 6111
rect 89576 6094 89593 6111
rect 90772 6094 90789 6111
rect 94360 6094 94377 6111
rect 94774 6094 94791 6111
rect 95188 6094 95205 6111
rect 97212 6094 97229 6111
rect 98224 6094 98241 6111
rect 98362 6094 98379 6111
rect 98730 6094 98747 6111
rect 100524 6094 100541 6111
rect 100938 6094 100955 6111
rect 101628 6094 101645 6111
rect 113772 6094 113789 6111
rect 114968 6094 114985 6111
rect 116072 6094 116089 6111
rect 119016 6094 119033 6111
rect 119568 6094 119585 6111
rect 119614 6094 119631 6111
rect 120074 6094 120091 6111
rect 120626 6094 120643 6111
rect 121868 6094 121885 6111
rect 122190 6094 122207 6111
rect 125640 6094 125657 6111
rect 125962 6094 125979 6111
rect 127572 6094 127589 6111
rect 128124 6094 128141 6111
rect 128538 6094 128555 6111
rect 131344 6094 131361 6111
rect 131988 6094 132005 6111
rect 132402 6094 132419 6111
rect 133276 6094 133293 6111
rect 135484 6094 135501 6111
rect 136036 6094 136053 6111
rect 14918 6060 14935 6077
rect 16022 6060 16039 6077
rect 17724 6060 17741 6077
rect 20852 6060 20869 6077
rect 26326 6060 26343 6077
rect 27752 6060 27769 6077
rect 50384 6060 50401 6077
rect 50430 6060 50447 6077
rect 50982 6060 50999 6077
rect 51074 6060 51091 6077
rect 57330 6060 57347 6077
rect 58756 6060 58773 6077
rect 64690 6060 64707 6077
rect 69014 6060 69031 6077
rect 72924 6060 72941 6077
rect 73108 6060 73125 6077
rect 76834 6060 76851 6077
rect 81940 6060 81957 6077
rect 82952 6060 82969 6077
rect 88978 6060 88995 6077
rect 89714 6060 89731 6077
rect 95556 6060 95573 6077
rect 96706 6060 96723 6077
rect 97350 6060 97367 6077
rect 102502 6060 102519 6077
rect 124536 6060 124553 6077
rect 124628 6060 124645 6077
rect 126422 6060 126439 6077
rect 132816 6060 132833 6077
rect 133414 6060 133431 6077
rect 134518 6060 134535 6077
rect 13538 6026 13555 6043
rect 13768 6026 13785 6043
rect 14136 6026 14153 6043
rect 16758 6026 16775 6043
rect 18230 6026 18247 6043
rect 20116 6026 20133 6043
rect 20346 6026 20363 6043
rect 28028 6026 28045 6043
rect 28074 6026 28091 6043
rect 28258 6026 28275 6043
rect 38148 6026 38165 6043
rect 38930 6026 38947 6043
rect 42012 6026 42029 6043
rect 43392 6026 43409 6043
rect 43806 6026 43823 6043
rect 44036 6026 44053 6043
rect 50200 6026 50217 6043
rect 51304 6026 51321 6043
rect 51534 6026 51551 6043
rect 58066 6026 58083 6043
rect 58572 6026 58589 6043
rect 64230 6026 64247 6043
rect 65656 6026 65673 6043
rect 65886 6026 65903 6043
rect 75362 6026 75379 6043
rect 75822 6026 75839 6043
rect 76006 6026 76023 6043
rect 76880 6026 76897 6043
rect 80422 6026 80439 6043
rect 81020 6026 81037 6043
rect 81204 6026 81221 6043
rect 88288 6026 88305 6043
rect 89024 6026 89041 6043
rect 94820 6026 94837 6043
rect 96522 6026 96539 6043
rect 96752 6026 96769 6043
rect 98408 6026 98425 6043
rect 98500 6026 98517 6043
rect 98684 6026 98701 6043
rect 101444 6026 101461 6043
rect 101674 6026 101691 6043
rect 114646 6026 114663 6043
rect 115474 6026 115491 6043
rect 115658 6026 115675 6043
rect 115704 6026 115721 6043
rect 119108 6026 119125 6043
rect 120442 6026 120459 6043
rect 120672 6026 120689 6043
rect 121362 6026 121379 6043
rect 127388 6026 127405 6043
rect 127618 6026 127635 6043
rect 132632 6026 132649 6043
rect 134150 6026 134167 6043
rect 135254 6026 135271 6043
rect 136082 6026 136099 6043
rect 13906 5924 13923 5941
rect 16298 5924 16315 5941
rect 16896 5924 16913 5941
rect 17218 5924 17235 5941
rect 17494 5924 17511 5941
rect 19196 5924 19213 5941
rect 19518 5924 19535 5941
rect 19840 5924 19857 5941
rect 20070 5924 20087 5941
rect 20576 5924 20593 5941
rect 20852 5924 20869 5941
rect 26418 5924 26435 5941
rect 26832 5924 26849 5941
rect 27200 5924 27217 5941
rect 27660 5924 27677 5941
rect 28258 5924 28275 5941
rect 28580 5924 28597 5941
rect 37780 5924 37797 5941
rect 38010 5924 38027 5941
rect 38470 5924 38487 5941
rect 38930 5924 38947 5941
rect 39252 5924 39269 5941
rect 42196 5924 42213 5941
rect 43024 5924 43041 5941
rect 43576 5924 43593 5941
rect 43944 5924 43961 5941
rect 44450 5924 44467 5941
rect 50108 5924 50125 5941
rect 50476 5924 50493 5941
rect 50936 5924 50953 5941
rect 56916 5924 56933 5941
rect 57514 5924 57531 5941
rect 58112 5924 58129 5941
rect 58480 5924 58497 5941
rect 58802 5924 58819 5941
rect 64690 5924 64707 5941
rect 65242 5924 65259 5941
rect 65472 5924 65489 5941
rect 66208 5924 66225 5941
rect 75546 5924 75563 5941
rect 76006 5924 76023 5941
rect 76374 5924 76391 5941
rect 81158 5924 81175 5941
rect 81480 5924 81497 5941
rect 81756 5924 81773 5941
rect 82124 5924 82141 5941
rect 82446 5924 82463 5941
rect 88242 5924 88259 5941
rect 88794 5924 88811 5941
rect 89024 5924 89041 5941
rect 89576 5924 89593 5941
rect 90036 5924 90053 5941
rect 95418 5924 95435 5941
rect 98132 5924 98149 5941
rect 101444 5924 101461 5941
rect 102042 5924 102059 5941
rect 102594 5924 102611 5941
rect 114140 5924 114157 5941
rect 114738 5924 114755 5941
rect 115198 5924 115215 5941
rect 115796 5924 115813 5941
rect 119384 5924 119401 5941
rect 120166 5924 120183 5941
rect 120534 5924 120551 5941
rect 120902 5924 120919 5941
rect 125916 5924 125933 5941
rect 127066 5924 127083 5941
rect 127480 5924 127497 5941
rect 127802 5924 127819 5941
rect 132494 5924 132511 5941
rect 133690 5924 133707 5941
rect 134104 5924 134121 5941
rect 135714 5924 135731 5941
rect 14412 5890 14429 5907
rect 20024 5890 20041 5907
rect 101168 5890 101185 5907
rect 101996 5890 102013 5907
rect 102640 5890 102657 5907
rect 114186 5890 114203 5907
rect 114784 5890 114801 5907
rect 119338 5890 119355 5907
rect 127020 5890 127037 5907
rect 132218 5890 132235 5907
rect 13998 5856 14015 5873
rect 14826 5856 14843 5873
rect 16252 5856 16269 5873
rect 16850 5856 16867 5873
rect 17172 5856 17189 5873
rect 17586 5856 17603 5873
rect 19288 5856 19305 5873
rect 19610 5856 19627 5873
rect 20530 5856 20547 5873
rect 20944 5856 20961 5873
rect 21450 5856 21467 5873
rect 26510 5856 26527 5873
rect 26924 5856 26941 5873
rect 27154 5856 27171 5873
rect 28212 5856 28229 5873
rect 28534 5856 28551 5873
rect 37964 5856 37981 5873
rect 38562 5856 38579 5873
rect 38884 5856 38901 5873
rect 39344 5856 39361 5873
rect 42288 5856 42305 5873
rect 42610 5856 42627 5873
rect 43070 5856 43087 5873
rect 43484 5856 43501 5873
rect 43898 5856 43915 5873
rect 44404 5856 44421 5873
rect 50200 5856 50217 5873
rect 50430 5856 50447 5873
rect 51580 5856 51597 5873
rect 57008 5856 57025 5873
rect 57560 5856 57577 5873
rect 58204 5856 58221 5873
rect 58434 5856 58451 5873
rect 58756 5856 58773 5873
rect 64644 5856 64661 5873
rect 65426 5856 65443 5873
rect 65840 5856 65857 5873
rect 66300 5856 66317 5873
rect 73890 5856 73907 5873
rect 75638 5856 75655 5873
rect 76098 5856 76115 5873
rect 76328 5856 76345 5873
rect 80560 5856 80577 5873
rect 80882 5856 80899 5873
rect 81112 5856 81129 5873
rect 81434 5856 81451 5873
rect 81848 5856 81865 5873
rect 82078 5856 82095 5873
rect 82400 5856 82417 5873
rect 88334 5856 88351 5873
rect 88978 5856 88995 5873
rect 89622 5856 89639 5873
rect 89990 5856 90007 5873
rect 94820 5856 94837 5873
rect 95050 5856 95067 5873
rect 95372 5856 95389 5873
rect 95924 5856 95941 5873
rect 97028 5856 97045 5873
rect 98224 5856 98241 5873
rect 101122 5856 101139 5873
rect 101536 5856 101553 5873
rect 115152 5856 115169 5873
rect 115474 5856 115491 5873
rect 115520 5856 115537 5873
rect 115888 5856 115905 5873
rect 120120 5856 120137 5873
rect 120626 5856 120643 5873
rect 120856 5856 120873 5873
rect 121270 5856 121287 5873
rect 126008 5856 126025 5873
rect 126192 5856 126209 5873
rect 126376 5856 126393 5873
rect 127434 5856 127451 5873
rect 127756 5856 127773 5873
rect 132172 5856 132189 5873
rect 132586 5856 132603 5873
rect 132816 5856 132833 5873
rect 134564 5856 134581 5873
rect 135668 5856 135685 5873
rect 14458 5822 14475 5839
rect 14550 5822 14567 5839
rect 14964 5822 14981 5839
rect 16344 5822 16361 5839
rect 20116 5822 20133 5839
rect 21542 5822 21559 5839
rect 27706 5822 27723 5839
rect 27798 5822 27815 5839
rect 38102 5822 38119 5839
rect 43162 5822 43179 5839
rect 50982 5822 50999 5839
rect 51028 5822 51045 5839
rect 57652 5822 57669 5839
rect 65518 5822 65535 5839
rect 74166 5822 74183 5839
rect 74304 5822 74321 5839
rect 89070 5822 89087 5839
rect 89668 5822 89685 5839
rect 96062 5822 96079 5839
rect 97166 5822 97183 5839
rect 97902 5822 97919 5839
rect 102134 5822 102151 5839
rect 102732 5822 102749 5839
rect 114232 5822 114249 5839
rect 114876 5822 114893 5839
rect 120212 5822 120229 5839
rect 127112 5822 127129 5839
rect 132954 5822 132971 5839
rect 134150 5822 134167 5839
rect 134196 5822 134213 5839
rect 134702 5822 134719 5839
rect 135438 5822 135455 5839
rect 21726 5788 21743 5805
rect 73798 5788 73815 5805
rect 80468 5788 80485 5805
rect 80790 5788 80807 5805
rect 89392 5788 89409 5805
rect 95096 5788 95113 5805
rect 113956 5788 113973 5805
rect 119936 5788 119953 5805
rect 126468 5788 126485 5805
rect 14228 5754 14245 5771
rect 15700 5754 15717 5771
rect 16068 5754 16085 5771
rect 27476 5754 27493 5771
rect 42518 5754 42535 5771
rect 42840 5754 42857 5771
rect 50752 5754 50769 5771
rect 51488 5754 51505 5771
rect 57330 5754 57347 5771
rect 65932 5754 65949 5771
rect 75040 5754 75057 5771
rect 94728 5754 94745 5771
rect 96798 5754 96815 5771
rect 101812 5754 101829 5771
rect 102410 5754 102427 5771
rect 114554 5754 114571 5771
rect 121178 5754 121195 5771
rect 126836 5754 126853 5771
rect 133920 5754 133937 5771
rect 14412 5652 14429 5669
rect 16804 5652 16821 5669
rect 20162 5652 20179 5669
rect 20530 5652 20547 5669
rect 20806 5652 20823 5669
rect 27660 5652 27677 5669
rect 28120 5652 28137 5669
rect 38240 5652 38257 5669
rect 39114 5652 39131 5669
rect 43116 5652 43133 5669
rect 43484 5652 43501 5669
rect 44128 5652 44145 5669
rect 51442 5652 51459 5669
rect 58020 5652 58037 5669
rect 58572 5652 58589 5669
rect 65242 5652 65259 5669
rect 65610 5652 65627 5669
rect 65886 5652 65903 5669
rect 74028 5652 74045 5669
rect 75408 5652 75425 5669
rect 78674 5652 78691 5669
rect 81020 5652 81037 5669
rect 81342 5652 81359 5669
rect 81802 5652 81819 5669
rect 119982 5652 119999 5669
rect 120442 5652 120459 5669
rect 120718 5652 120735 5669
rect 121086 5652 121103 5669
rect 126284 5652 126301 5669
rect 126560 5652 126577 5669
rect 126882 5652 126899 5669
rect 132770 5652 132787 5669
rect 134012 5652 134029 5669
rect 21128 5618 21145 5635
rect 43806 5618 43823 5635
rect 51764 5618 51781 5635
rect 57698 5618 57715 5635
rect 74948 5618 74965 5635
rect 127204 5618 127221 5635
rect 133414 5618 133431 5635
rect 14826 5584 14843 5601
rect 16160 5584 16177 5601
rect 16252 5584 16269 5601
rect 51166 5584 51183 5601
rect 74258 5584 74275 5601
rect 74350 5584 74367 5601
rect 88794 5584 88811 5601
rect 89116 5584 89133 5601
rect 95142 5584 95159 5601
rect 96016 5584 96033 5601
rect 96890 5584 96907 5601
rect 97488 5584 97505 5601
rect 101444 5584 101461 5601
rect 132494 5584 132511 5601
rect 133736 5584 133753 5601
rect 134288 5584 134305 5601
rect 134702 5584 134719 5601
rect 135300 5584 135317 5601
rect 14504 5550 14521 5567
rect 16114 5550 16131 5567
rect 16758 5550 16775 5567
rect 20254 5550 20271 5567
rect 20484 5550 20501 5567
rect 20898 5550 20915 5567
rect 21220 5550 21237 5567
rect 27752 5550 27769 5567
rect 28212 5550 28229 5567
rect 38332 5550 38349 5567
rect 39206 5550 39223 5567
rect 43208 5550 43225 5567
rect 43438 5550 43455 5567
rect 43898 5550 43915 5567
rect 44220 5550 44237 5567
rect 51074 5550 51091 5567
rect 51534 5550 51551 5567
rect 51856 5550 51873 5567
rect 57652 5550 57669 5567
rect 58112 5550 58129 5567
rect 58664 5550 58681 5567
rect 65334 5550 65351 5567
rect 65564 5550 65581 5567
rect 65978 5550 65995 5567
rect 71038 5550 71055 5567
rect 75500 5550 75517 5567
rect 81112 5550 81129 5567
rect 81434 5550 81451 5567
rect 81756 5550 81773 5567
rect 88748 5550 88765 5567
rect 89070 5550 89087 5567
rect 89576 5550 89593 5567
rect 95096 5550 95113 5567
rect 95418 5550 95435 5567
rect 95464 5550 95481 5567
rect 97396 5550 97413 5567
rect 97902 5550 97919 5567
rect 101168 5550 101185 5567
rect 101398 5550 101415 5567
rect 101720 5550 101737 5567
rect 102456 5550 102473 5567
rect 114692 5550 114709 5567
rect 119936 5550 119953 5567
rect 120396 5550 120413 5567
rect 120810 5550 120827 5567
rect 121040 5550 121057 5567
rect 126238 5550 126255 5567
rect 126652 5550 126669 5567
rect 126974 5550 126991 5567
rect 127296 5550 127313 5567
rect 132448 5550 132465 5567
rect 132862 5550 132879 5567
rect 133598 5550 133615 5567
rect 134104 5550 134121 5567
rect 135208 5550 135225 5567
rect 135254 5550 135271 5567
rect 14964 5516 14981 5533
rect 70210 5516 70227 5533
rect 74810 5516 74827 5533
rect 78030 5516 78047 5533
rect 96154 5516 96171 5533
rect 133644 5516 133661 5533
rect 134610 5516 134627 5533
rect 134656 5516 134673 5533
rect 15700 5482 15717 5499
rect 15930 5482 15947 5499
rect 74212 5482 74229 5499
rect 89484 5482 89501 5499
rect 97212 5482 97229 5499
rect 97442 5482 97459 5499
rect 97810 5482 97827 5499
rect 101076 5482 101093 5499
rect 101766 5482 101783 5499
rect 102364 5482 102381 5499
rect 114600 5482 114617 5499
rect 134426 5482 134443 5499
rect 135024 5482 135041 5499
rect 14826 5380 14843 5397
rect 15332 5380 15349 5397
rect 15378 5380 15395 5397
rect 16068 5380 16085 5397
rect 16390 5380 16407 5397
rect 16712 5380 16729 5397
rect 50844 5380 50861 5397
rect 65242 5380 65259 5397
rect 70992 5380 71009 5397
rect 74442 5380 74459 5397
rect 75362 5380 75379 5397
rect 95924 5380 95941 5397
rect 97120 5380 97137 5397
rect 101444 5380 101461 5397
rect 126836 5380 126853 5397
rect 133276 5380 133293 5397
rect 133874 5380 133891 5397
rect 134196 5380 134213 5397
rect 70348 5346 70365 5363
rect 78076 5346 78093 5363
rect 96752 5346 96769 5363
rect 14918 5312 14935 5329
rect 16160 5312 16177 5329
rect 16482 5312 16499 5329
rect 16804 5312 16821 5329
rect 50936 5312 50953 5329
rect 65196 5312 65213 5329
rect 74534 5312 74551 5329
rect 75316 5312 75333 5329
rect 93624 5312 93641 5329
rect 95648 5312 95665 5329
rect 96016 5312 96033 5329
rect 96338 5312 96355 5329
rect 97074 5312 97091 5329
rect 101536 5312 101553 5329
rect 126928 5312 126945 5329
rect 133000 5312 133017 5329
rect 133230 5312 133247 5329
rect 133552 5312 133569 5329
rect 133966 5312 133983 5329
rect 134288 5312 134305 5329
rect 134564 5312 134581 5329
rect 134610 5312 134627 5329
rect 15424 5278 15441 5295
rect 93762 5278 93779 5295
rect 15148 5244 15165 5261
rect 95556 5244 95573 5261
rect 96430 5244 96447 5261
rect 96844 5244 96861 5261
rect 133598 5244 133615 5261
rect 78812 5210 78829 5227
rect 132908 5210 132925 5227
rect 15470 5108 15487 5125
rect 15838 5108 15855 5125
rect 16436 5108 16453 5125
rect 16804 5108 16821 5125
rect 95924 5108 95941 5125
rect 96568 5108 96585 5125
rect 133874 5108 133891 5125
rect 134518 5108 134535 5125
rect 15148 5074 15165 5091
rect 16160 5074 16177 5091
rect 133552 5074 133569 5091
rect 134242 5074 134259 5091
rect 78904 5040 78921 5057
rect 15240 5006 15257 5023
rect 15562 5006 15579 5023
rect 15792 5006 15809 5023
rect 16114 5006 16131 5023
rect 16528 5006 16545 5023
rect 16758 5006 16775 5023
rect 70210 5006 70227 5023
rect 78030 5006 78047 5023
rect 96016 5006 96033 5023
rect 96338 5006 96355 5023
rect 96660 5006 96677 5023
rect 133644 5006 133661 5023
rect 133966 5006 133983 5023
rect 134196 5006 134213 5023
rect 134610 5006 134627 5023
rect 152228 5006 152245 5023
rect 152412 4972 152429 4989
rect 70854 4938 70871 4955
rect 96246 4938 96263 4955
rect 16436 4802 16453 4819
rect 70348 4802 70365 4819
rect 78076 4802 78093 4819
rect 78950 4802 78967 4819
rect 96522 4802 96539 4819
rect 133966 4802 133983 4819
rect 15654 4768 15671 4785
rect 16068 4768 16085 4785
rect 16390 4768 16407 4785
rect 96246 4768 96263 4785
rect 96476 4768 96493 4785
rect 133920 4768 133937 4785
rect 16114 4734 16131 4751
rect 15562 4700 15579 4717
rect 96154 4700 96171 4717
rect 70992 4666 71009 4683
rect 796 4224 813 4241
rect 704 4156 721 4173
rect 980 4156 997 4173
rect 1164 4156 1181 4173
rect 1348 4156 1365 4173
rect 1532 4156 1549 4173
rect 151998 3136 152015 3153
rect 152136 3102 152153 3119
<< metal1 >>
rect 94951 6926 94954 6932
rect 36172 6912 37750 6926
rect 14497 6872 14500 6898
rect 14526 6892 14529 6898
rect 16475 6892 16478 6898
rect 14526 6878 16478 6892
rect 14526 6872 14529 6878
rect 16475 6872 16478 6878
rect 16504 6872 16507 6898
rect 23099 6872 23102 6898
rect 23128 6892 23131 6898
rect 31701 6892 31704 6898
rect 23128 6878 31704 6892
rect 23128 6872 23131 6878
rect 31701 6872 31704 6878
rect 31730 6872 31733 6898
rect 34645 6872 34648 6898
rect 34674 6892 34677 6898
rect 36172 6892 36186 6912
rect 37681 6892 37684 6898
rect 34674 6878 36186 6892
rect 36218 6878 37684 6892
rect 34674 6872 34677 6878
rect 36218 6864 36232 6878
rect 37681 6872 37684 6878
rect 37710 6872 37713 6898
rect 37736 6892 37750 6912
rect 94638 6912 94954 6926
rect 38003 6892 38006 6898
rect 37736 6878 38006 6892
rect 38003 6872 38006 6878
rect 38032 6872 38035 6898
rect 45317 6872 45320 6898
rect 45346 6892 45349 6898
rect 51205 6892 51208 6898
rect 45346 6878 51208 6892
rect 45346 6872 45349 6878
rect 51205 6872 51208 6878
rect 51234 6872 51237 6898
rect 56909 6872 56912 6898
rect 56938 6892 56941 6898
rect 62751 6892 62754 6898
rect 56938 6878 62754 6892
rect 56938 6872 56941 6878
rect 62751 6872 62754 6878
rect 62780 6892 62783 6898
rect 65925 6892 65928 6898
rect 62780 6878 65928 6892
rect 62780 6872 62783 6878
rect 65925 6872 65928 6878
rect 65954 6872 65957 6898
rect 80829 6872 80832 6898
rect 80858 6892 80861 6898
rect 83037 6892 83040 6898
rect 80858 6878 83040 6892
rect 80858 6872 80861 6878
rect 83037 6872 83040 6878
rect 83066 6892 83069 6898
rect 83681 6892 83684 6898
rect 83066 6878 83684 6892
rect 83066 6872 83069 6878
rect 83681 6872 83684 6878
rect 83710 6872 83713 6898
rect 87085 6872 87088 6898
rect 87114 6892 87117 6898
rect 88879 6892 88882 6898
rect 87114 6878 88882 6892
rect 87114 6872 87117 6878
rect 88879 6872 88882 6878
rect 88908 6872 88911 6898
rect 90949 6872 90952 6898
rect 90978 6892 90981 6898
rect 94638 6892 94652 6912
rect 94951 6906 94954 6912
rect 94980 6906 94983 6932
rect 90978 6878 94652 6892
rect 90978 6872 90981 6878
rect 94675 6872 94678 6898
rect 94704 6892 94707 6898
rect 96607 6892 96610 6898
rect 94704 6878 96610 6892
rect 94704 6872 94707 6878
rect 96607 6872 96610 6878
rect 96636 6872 96639 6898
rect 97987 6872 97990 6898
rect 98016 6892 98019 6898
rect 151393 6892 151396 6898
rect 98016 6878 151396 6892
rect 98016 6872 98019 6878
rect 151393 6872 151396 6878
rect 151422 6872 151425 6898
rect 13577 6838 13580 6864
rect 13606 6858 13609 6864
rect 18269 6858 18272 6864
rect 13606 6844 18272 6858
rect 13606 6838 13609 6844
rect 18269 6838 18272 6844
rect 18298 6838 18301 6864
rect 21259 6838 21262 6864
rect 21288 6858 21291 6864
rect 23927 6858 23930 6864
rect 21288 6844 23930 6858
rect 21288 6838 21291 6844
rect 23927 6838 23930 6844
rect 23956 6838 23959 6864
rect 25813 6838 25816 6864
rect 25842 6858 25845 6864
rect 27055 6858 27058 6864
rect 25842 6844 27058 6858
rect 25842 6838 25845 6844
rect 27055 6838 27058 6844
rect 27084 6838 27087 6864
rect 33081 6838 33084 6864
rect 33110 6858 33113 6864
rect 36209 6858 36212 6864
rect 33110 6844 36212 6858
rect 33110 6838 33113 6844
rect 36209 6838 36212 6844
rect 36238 6838 36241 6864
rect 36945 6838 36948 6864
rect 36974 6858 36977 6864
rect 38187 6858 38190 6864
rect 36974 6844 38190 6858
rect 36974 6838 36977 6844
rect 38187 6838 38190 6844
rect 38216 6838 38219 6864
rect 41545 6838 41548 6864
rect 41574 6858 41577 6864
rect 43201 6858 43204 6864
rect 41574 6844 43204 6858
rect 41574 6838 41577 6844
rect 43201 6838 43204 6844
rect 43230 6838 43233 6864
rect 45915 6838 45918 6864
rect 45944 6858 45947 6864
rect 50975 6858 50978 6864
rect 45944 6844 50978 6858
rect 45944 6838 45947 6844
rect 50975 6838 50978 6844
rect 51004 6838 51007 6864
rect 57323 6838 57326 6864
rect 57352 6858 57355 6864
rect 63717 6858 63720 6864
rect 57352 6844 63720 6858
rect 57352 6838 57355 6844
rect 63717 6838 63720 6844
rect 63746 6838 63749 6864
rect 63763 6838 63766 6864
rect 63792 6858 63795 6864
rect 64867 6858 64870 6864
rect 63792 6844 64870 6858
rect 63792 6838 63795 6844
rect 64867 6838 64870 6844
rect 64896 6838 64899 6864
rect 66799 6838 66802 6864
rect 66828 6858 66831 6864
rect 68409 6858 68412 6864
rect 66828 6844 68412 6858
rect 66828 6838 66831 6844
rect 68409 6838 68412 6844
rect 68438 6838 68441 6864
rect 74067 6838 74070 6864
rect 74096 6858 74099 6864
rect 75217 6858 75220 6864
rect 74096 6844 75220 6858
rect 74096 6838 74099 6844
rect 75217 6838 75220 6844
rect 75246 6838 75249 6864
rect 78575 6838 78578 6864
rect 78604 6858 78607 6864
rect 150703 6858 150706 6864
rect 78604 6844 150706 6858
rect 78604 6838 78607 6844
rect 150703 6838 150706 6844
rect 150732 6838 150735 6864
rect 552 6813 152904 6824
rect 552 6787 19524 6813
rect 19550 6787 19556 6813
rect 19582 6787 19588 6813
rect 19614 6787 19620 6813
rect 19646 6787 19652 6813
rect 19678 6787 57623 6813
rect 57649 6787 57655 6813
rect 57681 6787 57687 6813
rect 57713 6787 57719 6813
rect 57745 6787 57751 6813
rect 57777 6787 95722 6813
rect 95748 6787 95754 6813
rect 95780 6787 95786 6813
rect 95812 6787 95818 6813
rect 95844 6787 95850 6813
rect 95876 6787 133821 6813
rect 133847 6787 133853 6813
rect 133879 6787 133885 6813
rect 133911 6787 133917 6813
rect 133943 6787 133949 6813
rect 133975 6787 152904 6813
rect 552 6776 152904 6787
rect 789 6756 792 6762
rect 769 6742 792 6756
rect 789 6736 792 6742
rect 818 6736 821 6762
rect 2307 6756 2310 6762
rect 2287 6742 2310 6756
rect 2307 6736 2310 6742
rect 2336 6736 2339 6762
rect 3825 6756 3828 6762
rect 3805 6742 3828 6756
rect 3825 6736 3828 6742
rect 3854 6736 3857 6762
rect 5389 6756 5392 6762
rect 5369 6742 5392 6756
rect 5389 6736 5392 6742
rect 5418 6736 5421 6762
rect 6907 6736 6910 6762
rect 6936 6756 6939 6762
rect 7046 6757 7075 6760
rect 7046 6756 7052 6757
rect 6936 6742 7052 6756
rect 6936 6736 6939 6742
rect 7046 6740 7052 6742
rect 7069 6740 7075 6757
rect 8425 6756 8428 6762
rect 8405 6742 8428 6756
rect 7046 6737 7075 6740
rect 8425 6736 8428 6742
rect 8454 6736 8457 6762
rect 9989 6756 9992 6762
rect 9969 6742 9992 6756
rect 9989 6736 9992 6742
rect 10018 6736 10021 6762
rect 11507 6756 11510 6762
rect 11487 6742 11510 6756
rect 11507 6736 11510 6742
rect 11536 6736 11539 6762
rect 12842 6757 12871 6760
rect 12842 6740 12848 6757
rect 12865 6756 12871 6757
rect 13807 6756 13810 6762
rect 12865 6742 13810 6756
rect 12865 6740 12871 6742
rect 12842 6737 12871 6740
rect 13807 6736 13810 6742
rect 13836 6736 13839 6762
rect 13853 6736 13856 6762
rect 13882 6756 13885 6762
rect 14498 6757 14527 6760
rect 14498 6756 14504 6757
rect 13882 6742 14504 6756
rect 13882 6736 13885 6742
rect 14498 6740 14504 6742
rect 14521 6740 14527 6757
rect 14498 6737 14527 6740
rect 15233 6736 15236 6762
rect 15262 6756 15265 6762
rect 15786 6757 15815 6760
rect 15786 6756 15792 6757
rect 15262 6742 15792 6756
rect 15262 6736 15265 6742
rect 15786 6740 15792 6742
rect 15809 6740 15815 6757
rect 15786 6737 15815 6740
rect 18269 6736 18272 6762
rect 18298 6756 18301 6762
rect 23099 6756 23102 6762
rect 18298 6742 23102 6756
rect 18298 6736 18301 6742
rect 23099 6736 23102 6742
rect 23128 6736 23131 6762
rect 23789 6756 23792 6762
rect 23769 6742 23792 6756
rect 23789 6736 23792 6742
rect 23818 6736 23821 6762
rect 25170 6757 25199 6760
rect 25170 6740 25176 6757
rect 25193 6756 25199 6757
rect 25261 6756 25264 6762
rect 25193 6742 25264 6756
rect 25193 6740 25199 6742
rect 25170 6737 25199 6740
rect 25261 6736 25264 6742
rect 25290 6736 25293 6762
rect 25492 6757 25521 6760
rect 25492 6740 25498 6757
rect 25515 6756 25521 6757
rect 26503 6756 26506 6762
rect 25515 6742 26506 6756
rect 25515 6740 25521 6742
rect 25492 6737 25521 6740
rect 26503 6736 26506 6742
rect 26532 6736 26535 6762
rect 27791 6736 27794 6762
rect 27820 6756 27823 6762
rect 28941 6756 28944 6762
rect 27820 6742 28944 6756
rect 27820 6736 27823 6742
rect 28941 6736 28944 6742
rect 28970 6756 28973 6762
rect 30873 6756 30876 6762
rect 28970 6742 30876 6756
rect 28970 6736 28973 6742
rect 30873 6736 30876 6742
rect 30902 6736 30905 6762
rect 31701 6736 31704 6762
rect 31730 6756 31733 6762
rect 71445 6756 71448 6762
rect 31730 6742 71077 6756
rect 71425 6742 71448 6756
rect 31730 6736 31733 6742
rect 13577 6722 13580 6728
rect 3443 6708 13580 6722
rect 3443 6688 3457 6708
rect 13577 6702 13580 6708
rect 13606 6702 13609 6728
rect 22087 6702 22090 6728
rect 22116 6702 22119 6728
rect 22134 6723 22163 6726
rect 22134 6706 22140 6723
rect 22157 6706 22163 6723
rect 22134 6703 22163 6706
rect 13164 6689 13193 6692
rect 890 6674 3457 6688
rect 5490 6674 13048 6688
rect 890 6658 904 6674
rect 882 6655 911 6658
rect 882 6638 888 6655
rect 905 6638 911 6655
rect 2399 6654 2402 6660
rect 2379 6640 2402 6654
rect 882 6635 911 6638
rect 2399 6634 2402 6640
rect 2428 6634 2431 6660
rect 5490 6658 5504 6674
rect 3918 6655 3947 6658
rect 3918 6638 3924 6655
rect 3941 6638 3947 6655
rect 3918 6635 3947 6638
rect 5482 6655 5511 6658
rect 5482 6638 5488 6655
rect 5505 6638 5511 6655
rect 7137 6654 7140 6660
rect 7117 6640 7140 6654
rect 5482 6635 5511 6638
rect 3926 6620 3940 6635
rect 7137 6634 7140 6640
rect 7166 6634 7169 6660
rect 8517 6654 8520 6660
rect 8497 6640 8520 6654
rect 8517 6634 8520 6640
rect 8546 6634 8549 6660
rect 10081 6654 10084 6660
rect 10061 6640 10084 6654
rect 10081 6634 10084 6640
rect 10110 6634 10113 6660
rect 11599 6654 11602 6660
rect 11579 6640 11602 6654
rect 11599 6634 11602 6640
rect 11628 6634 11631 6660
rect 13034 6658 13048 6674
rect 13164 6672 13170 6689
rect 13187 6688 13193 6689
rect 13485 6688 13488 6694
rect 13187 6674 13488 6688
rect 13187 6672 13193 6674
rect 13164 6669 13193 6672
rect 13485 6668 13488 6674
rect 13514 6668 13517 6694
rect 13624 6689 13653 6692
rect 13624 6672 13630 6689
rect 13647 6688 13653 6689
rect 17350 6689 17379 6692
rect 17350 6688 17356 6689
rect 13647 6674 17356 6688
rect 13647 6672 13653 6674
rect 13624 6669 13653 6672
rect 17350 6672 17356 6674
rect 17373 6688 17379 6689
rect 18776 6689 18805 6692
rect 17373 6674 18522 6688
rect 17373 6672 17379 6674
rect 17350 6669 17379 6672
rect 13026 6655 13055 6658
rect 13026 6638 13032 6655
rect 13049 6638 13055 6655
rect 14911 6654 14914 6660
rect 14891 6640 14914 6654
rect 13026 6635 13055 6638
rect 13034 6620 13048 6635
rect 14911 6634 14914 6640
rect 14940 6634 14943 6660
rect 16199 6654 16202 6660
rect 16179 6640 16202 6654
rect 16199 6634 16202 6640
rect 16228 6634 16231 6660
rect 16889 6634 16892 6660
rect 16918 6634 16921 6660
rect 18508 6654 18522 6674
rect 18776 6672 18782 6689
rect 18799 6688 18805 6689
rect 22096 6688 22110 6702
rect 18799 6674 22110 6688
rect 18799 6672 18805 6674
rect 18776 6669 18805 6672
rect 22142 6660 22156 6703
rect 22179 6702 22182 6728
rect 22208 6722 22211 6728
rect 22208 6708 25928 6722
rect 22208 6702 22211 6708
rect 22777 6668 22780 6694
rect 22806 6688 22809 6694
rect 25813 6688 25816 6694
rect 22806 6674 22828 6688
rect 25793 6674 25816 6688
rect 22806 6668 22809 6674
rect 25813 6668 25816 6674
rect 25842 6668 25845 6694
rect 25914 6688 25928 6708
rect 29907 6702 29910 6728
rect 29936 6722 29939 6728
rect 30230 6723 30259 6726
rect 30230 6722 30236 6723
rect 29936 6708 30236 6722
rect 29936 6702 29939 6708
rect 30230 6706 30236 6708
rect 30253 6706 30259 6723
rect 31517 6722 31520 6728
rect 31497 6708 31520 6722
rect 30230 6703 30259 6706
rect 31517 6702 31520 6708
rect 31546 6702 31549 6728
rect 37681 6722 37684 6728
rect 31572 6708 36830 6722
rect 37661 6708 37684 6722
rect 31572 6688 31586 6708
rect 36347 6688 36350 6694
rect 25914 6674 31586 6688
rect 32423 6674 34714 6688
rect 36327 6674 36350 6688
rect 18508 6640 18798 6654
rect 13761 6620 13764 6626
rect 3926 6606 11047 6620
rect 13034 6606 13692 6620
rect 13741 6606 13764 6620
rect 11033 6586 11047 6606
rect 13072 6587 13101 6590
rect 13072 6586 13078 6587
rect 11033 6572 13078 6586
rect 13072 6570 13078 6572
rect 13095 6586 13101 6587
rect 13623 6586 13626 6592
rect 13095 6572 13626 6586
rect 13095 6570 13101 6572
rect 13072 6567 13101 6570
rect 13623 6566 13626 6572
rect 13652 6566 13655 6592
rect 13678 6586 13692 6606
rect 13761 6600 13764 6606
rect 13790 6600 13793 6626
rect 15050 6621 15079 6624
rect 14375 6606 14612 6620
rect 13853 6586 13856 6592
rect 13678 6572 13856 6586
rect 13853 6566 13856 6572
rect 13882 6566 13885 6592
rect 14598 6586 14612 6606
rect 15050 6604 15056 6621
rect 15073 6620 15079 6621
rect 15095 6620 15098 6626
rect 15073 6606 15098 6620
rect 15073 6604 15079 6606
rect 15050 6601 15079 6604
rect 15095 6600 15098 6606
rect 15124 6600 15127 6626
rect 16337 6620 16340 6626
rect 15663 6606 15877 6620
rect 16317 6606 16340 6620
rect 15233 6586 15236 6592
rect 14598 6572 15236 6586
rect 15233 6566 15236 6572
rect 15262 6566 15265 6592
rect 15863 6586 15877 6606
rect 16337 6600 16340 6606
rect 16366 6600 16369 6626
rect 17257 6600 17260 6626
rect 17286 6620 17289 6626
rect 17488 6621 17517 6624
rect 17488 6620 17494 6621
rect 17286 6606 17494 6620
rect 17286 6600 17289 6606
rect 17488 6604 17494 6606
rect 17511 6604 17517 6621
rect 17488 6601 17517 6604
rect 17993 6600 17996 6626
rect 18022 6600 18025 6626
rect 16797 6586 16800 6592
rect 15863 6572 16800 6586
rect 16797 6566 16800 6572
rect 16826 6566 16829 6592
rect 17073 6586 17076 6592
rect 17053 6572 17076 6586
rect 17073 6566 17076 6572
rect 17102 6566 17105 6592
rect 17165 6566 17168 6592
rect 17194 6586 17197 6592
rect 18224 6587 18253 6590
rect 18224 6586 18230 6587
rect 17194 6572 18230 6586
rect 17194 6566 17197 6572
rect 18224 6570 18230 6572
rect 18247 6586 18253 6587
rect 18729 6586 18732 6592
rect 18247 6572 18732 6586
rect 18247 6570 18253 6572
rect 18224 6567 18253 6570
rect 18729 6566 18732 6572
rect 18758 6566 18761 6592
rect 18784 6586 18798 6640
rect 19465 6634 19468 6660
rect 19494 6634 19497 6660
rect 20064 6655 20093 6658
rect 20064 6654 20070 6655
rect 19566 6640 20070 6654
rect 18913 6620 18916 6626
rect 18893 6606 18916 6620
rect 18913 6600 18916 6606
rect 18942 6600 18945 6626
rect 19566 6586 19580 6640
rect 20064 6638 20070 6640
rect 20087 6638 20093 6655
rect 21259 6654 21262 6660
rect 21239 6640 21262 6654
rect 20064 6635 20093 6638
rect 19649 6586 19652 6592
rect 18784 6572 19580 6586
rect 19629 6572 19652 6586
rect 19649 6566 19652 6572
rect 19678 6586 19681 6592
rect 19971 6586 19974 6592
rect 19678 6572 19974 6586
rect 19678 6566 19681 6572
rect 19971 6566 19974 6572
rect 20000 6566 20003 6592
rect 20072 6586 20086 6635
rect 21259 6634 21262 6640
rect 21288 6634 21291 6660
rect 22133 6634 22136 6660
rect 22162 6654 22165 6660
rect 23882 6655 23911 6658
rect 23882 6654 23888 6655
rect 22162 6640 23888 6654
rect 22162 6634 22165 6640
rect 23882 6638 23888 6640
rect 23905 6638 23911 6655
rect 23882 6635 23911 6638
rect 25262 6655 25291 6658
rect 25262 6638 25268 6655
rect 25285 6654 25291 6655
rect 25675 6654 25678 6660
rect 25285 6640 25678 6654
rect 25285 6638 25291 6640
rect 25262 6635 25291 6638
rect 20201 6620 20204 6626
rect 20181 6606 20204 6620
rect 20201 6600 20204 6606
rect 20230 6600 20233 6626
rect 20707 6600 20710 6626
rect 20736 6600 20739 6626
rect 21268 6620 21282 6634
rect 20900 6606 21282 6620
rect 21398 6621 21427 6624
rect 20900 6586 20914 6606
rect 21398 6604 21404 6621
rect 21421 6620 21427 6621
rect 21443 6620 21446 6626
rect 21421 6606 21446 6620
rect 21421 6604 21427 6606
rect 21398 6601 21427 6604
rect 21443 6600 21446 6606
rect 21472 6600 21475 6626
rect 21627 6600 21630 6626
rect 21656 6600 21659 6626
rect 22732 6621 22761 6624
rect 22732 6620 22738 6621
rect 22234 6606 22738 6620
rect 20072 6572 20914 6586
rect 20938 6587 20967 6590
rect 20938 6570 20944 6587
rect 20961 6586 20967 6587
rect 21213 6586 21216 6592
rect 20961 6572 21216 6586
rect 20961 6570 20967 6572
rect 20938 6567 20967 6570
rect 21213 6566 21216 6572
rect 21242 6586 21245 6592
rect 22234 6586 22248 6606
rect 22732 6604 22738 6606
rect 22755 6604 22761 6621
rect 22732 6601 22761 6604
rect 22501 6586 22504 6592
rect 21242 6572 22248 6586
rect 22481 6572 22504 6586
rect 21242 6566 21245 6572
rect 22501 6566 22504 6572
rect 22530 6566 22533 6592
rect 22685 6586 22688 6592
rect 22665 6572 22688 6586
rect 22685 6566 22688 6572
rect 22714 6566 22717 6592
rect 23890 6586 23904 6635
rect 25675 6634 25678 6640
rect 25704 6634 25707 6660
rect 26504 6655 26533 6658
rect 26504 6638 26510 6655
rect 26527 6638 26533 6655
rect 26504 6635 26533 6638
rect 23927 6600 23930 6626
rect 23956 6620 23959 6626
rect 26512 6620 26526 6635
rect 27193 6634 27196 6660
rect 27222 6634 27225 6660
rect 27377 6634 27380 6660
rect 27406 6654 27409 6660
rect 27791 6654 27794 6660
rect 27406 6640 27794 6654
rect 27406 6634 27409 6640
rect 27791 6634 27794 6640
rect 27820 6634 27823 6660
rect 28941 6654 28944 6660
rect 28921 6640 28944 6654
rect 28941 6634 28944 6640
rect 28970 6634 28973 6660
rect 30321 6654 30324 6660
rect 30301 6640 30324 6654
rect 30321 6634 30324 6640
rect 30350 6634 30353 6660
rect 31610 6655 31639 6658
rect 31610 6654 31616 6655
rect 30790 6640 31616 6654
rect 26641 6620 26644 6626
rect 23956 6606 26526 6620
rect 26621 6606 26644 6620
rect 23956 6600 23959 6606
rect 25722 6587 25751 6590
rect 25722 6586 25728 6587
rect 23890 6572 25728 6586
rect 25722 6570 25728 6572
rect 25745 6570 25751 6587
rect 26512 6586 26526 6606
rect 26641 6600 26644 6606
rect 26670 6600 26673 6626
rect 27929 6620 27932 6626
rect 27294 6606 27492 6620
rect 27909 6606 27932 6620
rect 27294 6586 27308 6606
rect 26512 6572 27308 6586
rect 25722 6567 25751 6570
rect 27331 6566 27334 6592
rect 27360 6586 27363 6592
rect 27378 6587 27407 6590
rect 27378 6586 27384 6587
rect 27360 6572 27384 6586
rect 27360 6566 27363 6572
rect 27378 6570 27384 6572
rect 27401 6570 27407 6587
rect 27478 6586 27492 6606
rect 27929 6600 27932 6606
rect 27958 6600 27961 6626
rect 28297 6600 28300 6626
rect 28326 6600 28329 6626
rect 28582 6606 28734 6620
rect 28582 6586 28596 6606
rect 28665 6586 28668 6592
rect 27478 6572 28596 6586
rect 28645 6572 28668 6586
rect 27378 6567 27407 6570
rect 28665 6566 28668 6572
rect 28694 6566 28697 6592
rect 28720 6586 28734 6606
rect 28849 6600 28852 6626
rect 28878 6620 28881 6626
rect 29080 6621 29109 6624
rect 29080 6620 29086 6621
rect 28878 6606 29086 6620
rect 28878 6600 28881 6606
rect 29080 6604 29086 6606
rect 29103 6604 29109 6621
rect 29080 6601 29109 6604
rect 29309 6600 29312 6626
rect 29338 6600 29341 6626
rect 30735 6620 30738 6626
rect 29732 6606 30738 6620
rect 29732 6586 29746 6606
rect 30735 6600 30738 6606
rect 30764 6600 30767 6626
rect 29815 6586 29818 6592
rect 28720 6572 29746 6586
rect 29795 6572 29818 6586
rect 29815 6566 29818 6572
rect 29844 6586 29847 6592
rect 30790 6586 30804 6640
rect 31610 6638 31616 6640
rect 31633 6654 31639 6655
rect 32423 6654 32437 6674
rect 33081 6654 33084 6660
rect 31633 6652 31678 6654
rect 31710 6652 32437 6654
rect 31633 6640 32437 6652
rect 33061 6640 33084 6654
rect 31633 6638 31639 6640
rect 31610 6635 31639 6638
rect 31664 6638 31724 6640
rect 33081 6634 33084 6640
rect 33110 6634 33113 6660
rect 34645 6654 34648 6660
rect 34625 6640 34648 6654
rect 34645 6634 34648 6640
rect 34674 6634 34677 6660
rect 34700 6654 34714 6674
rect 36347 6668 36350 6674
rect 36376 6668 36379 6694
rect 36816 6692 36830 6708
rect 37681 6702 37684 6708
rect 37710 6722 37713 6728
rect 37819 6722 37822 6728
rect 37710 6708 37822 6722
rect 37710 6702 37713 6708
rect 37819 6702 37822 6708
rect 37848 6702 37851 6728
rect 40013 6708 41246 6722
rect 36808 6689 36837 6692
rect 36808 6672 36814 6689
rect 36831 6688 36837 6689
rect 39246 6689 39275 6692
rect 39246 6688 39252 6689
rect 36831 6674 39252 6688
rect 36831 6672 36837 6674
rect 36808 6669 36837 6672
rect 39246 6672 39252 6674
rect 39269 6688 39275 6689
rect 40013 6688 40027 6708
rect 40119 6688 40122 6694
rect 39269 6674 40027 6688
rect 40075 6674 40122 6688
rect 39269 6672 39275 6674
rect 39246 6669 39275 6672
rect 40119 6668 40122 6674
rect 40148 6688 40151 6694
rect 40764 6689 40793 6692
rect 40764 6688 40770 6689
rect 40148 6674 40770 6688
rect 40148 6668 40151 6674
rect 40764 6672 40770 6674
rect 40787 6672 40793 6689
rect 40764 6669 40793 6672
rect 40809 6668 40812 6694
rect 40838 6688 40841 6694
rect 41232 6688 41246 6708
rect 46927 6702 46930 6728
rect 46956 6722 46959 6728
rect 46974 6723 47003 6726
rect 46974 6722 46980 6723
rect 46956 6708 46980 6722
rect 46956 6702 46959 6708
rect 46974 6706 46980 6708
rect 46997 6706 47003 6723
rect 46974 6703 47003 6706
rect 47258 6708 49687 6722
rect 47258 6688 47272 6708
rect 48998 6689 49027 6692
rect 48998 6688 49004 6689
rect 40838 6674 40860 6688
rect 41232 6674 47272 6688
rect 47304 6674 49004 6688
rect 40838 6668 40841 6674
rect 36256 6655 36285 6658
rect 36256 6654 36262 6655
rect 34700 6640 36262 6654
rect 36256 6638 36262 6640
rect 36279 6638 36285 6655
rect 36256 6635 36285 6638
rect 38096 6655 38125 6658
rect 38096 6638 38102 6655
rect 38119 6638 38125 6655
rect 39199 6654 39202 6660
rect 38801 6640 39202 6654
rect 38096 6635 38125 6638
rect 30873 6600 30876 6626
rect 30902 6620 30905 6626
rect 30902 6606 36922 6620
rect 30902 6600 30905 6606
rect 29844 6572 30804 6586
rect 29844 6566 29847 6572
rect 30827 6566 30830 6592
rect 30856 6586 30859 6592
rect 32943 6586 32946 6592
rect 30856 6572 32946 6586
rect 30856 6566 30859 6572
rect 32943 6566 32946 6572
rect 32972 6566 32975 6592
rect 32989 6566 32992 6592
rect 33018 6586 33021 6592
rect 34553 6586 34556 6592
rect 33018 6572 33040 6586
rect 34533 6572 34556 6586
rect 33018 6566 33021 6572
rect 34553 6566 34556 6572
rect 34582 6566 34585 6592
rect 36026 6587 36055 6590
rect 36026 6570 36032 6587
rect 36049 6586 36055 6587
rect 36163 6586 36166 6592
rect 36049 6572 36166 6586
rect 36049 6570 36055 6572
rect 36026 6567 36055 6570
rect 36163 6566 36166 6572
rect 36192 6566 36195 6592
rect 36209 6566 36212 6592
rect 36238 6586 36241 6592
rect 36908 6586 36922 6606
rect 36945 6600 36948 6626
rect 36974 6620 36977 6626
rect 37589 6620 37592 6626
rect 36974 6606 36996 6620
rect 37559 6606 37592 6620
rect 36974 6600 36977 6606
rect 37589 6600 37592 6606
rect 37618 6600 37621 6626
rect 38104 6586 38118 6635
rect 39199 6634 39202 6640
rect 39228 6634 39231 6660
rect 40717 6634 40720 6660
rect 40746 6634 40749 6660
rect 41224 6655 41253 6658
rect 41224 6638 41230 6655
rect 41247 6638 41253 6655
rect 41545 6654 41548 6660
rect 41525 6640 41548 6654
rect 41224 6635 41253 6638
rect 38233 6620 38236 6626
rect 38213 6606 38236 6620
rect 38233 6600 38236 6606
rect 38262 6600 38265 6626
rect 39383 6620 39386 6626
rect 38932 6606 39084 6620
rect 39363 6606 39386 6620
rect 38932 6586 38946 6606
rect 36238 6572 36260 6586
rect 36908 6572 38946 6586
rect 36238 6566 36241 6572
rect 38969 6566 38972 6592
rect 38998 6586 39001 6592
rect 39070 6586 39084 6606
rect 39383 6600 39386 6606
rect 39412 6600 39415 6626
rect 39659 6600 39662 6626
rect 39688 6600 39691 6626
rect 40027 6600 40030 6626
rect 40056 6620 40059 6626
rect 40726 6620 40740 6634
rect 41232 6620 41246 6635
rect 41545 6634 41548 6640
rect 41574 6634 41577 6660
rect 41959 6654 41962 6660
rect 41939 6640 41962 6654
rect 41959 6634 41962 6640
rect 41988 6634 41991 6660
rect 43248 6655 43277 6658
rect 43248 6654 43254 6655
rect 42796 6640 43254 6654
rect 41913 6620 41916 6626
rect 40056 6606 40556 6620
rect 40726 6606 41154 6620
rect 41232 6606 41916 6620
rect 40056 6600 40059 6606
rect 40395 6586 40398 6592
rect 38998 6572 39020 6586
rect 39070 6572 40398 6586
rect 38998 6566 39001 6572
rect 40395 6566 40398 6572
rect 40424 6566 40427 6592
rect 40542 6590 40556 6606
rect 40534 6587 40563 6590
rect 40534 6570 40540 6587
rect 40557 6570 40563 6587
rect 40717 6586 40720 6592
rect 40697 6572 40720 6586
rect 40534 6567 40563 6570
rect 40717 6566 40720 6572
rect 40746 6566 40749 6592
rect 41140 6590 41154 6606
rect 41913 6600 41916 6606
rect 41942 6600 41945 6626
rect 42098 6621 42127 6624
rect 42098 6604 42104 6621
rect 42121 6620 42127 6621
rect 42235 6620 42238 6626
rect 42121 6606 42238 6620
rect 42121 6604 42127 6606
rect 42098 6601 42127 6604
rect 42235 6600 42238 6606
rect 42264 6600 42267 6626
rect 42741 6620 42744 6626
rect 42711 6606 42744 6620
rect 42741 6600 42744 6606
rect 42770 6600 42773 6626
rect 41132 6587 41161 6590
rect 41132 6570 41138 6587
rect 41155 6570 41161 6587
rect 41453 6586 41456 6592
rect 41433 6572 41456 6586
rect 41132 6567 41161 6570
rect 41453 6566 41456 6572
rect 41482 6566 41485 6592
rect 41959 6566 41962 6592
rect 41988 6586 41991 6592
rect 42796 6586 42810 6640
rect 43248 6638 43254 6640
rect 43271 6638 43277 6655
rect 43248 6635 43277 6638
rect 41988 6572 42810 6586
rect 42834 6587 42863 6590
rect 41988 6566 41991 6572
rect 42834 6570 42840 6587
rect 42857 6586 42863 6587
rect 43017 6586 43020 6592
rect 42857 6572 43020 6586
rect 42857 6570 42863 6572
rect 42834 6567 42863 6570
rect 43017 6566 43020 6572
rect 43046 6566 43049 6592
rect 43256 6586 43270 6635
rect 43937 6634 43940 6660
rect 43966 6634 43969 6660
rect 44398 6655 44427 6658
rect 44398 6654 44404 6655
rect 44038 6640 44404 6654
rect 43385 6620 43388 6626
rect 43365 6606 43388 6620
rect 43385 6600 43388 6606
rect 43414 6600 43417 6626
rect 44038 6586 44052 6640
rect 44398 6638 44404 6640
rect 44421 6638 44427 6655
rect 47066 6655 47095 6658
rect 47066 6654 47072 6655
rect 44398 6635 44427 6638
rect 46568 6640 47072 6654
rect 44121 6586 44124 6592
rect 43256 6572 44052 6586
rect 44101 6572 44124 6586
rect 44121 6566 44124 6572
rect 44150 6566 44153 6592
rect 44406 6586 44420 6635
rect 44535 6620 44538 6626
rect 44515 6606 44538 6620
rect 44535 6600 44538 6606
rect 44564 6600 44567 6626
rect 44765 6600 44768 6626
rect 44794 6600 44797 6626
rect 45823 6620 45826 6626
rect 45234 6606 45826 6620
rect 45234 6586 45248 6606
rect 45823 6600 45826 6606
rect 45852 6600 45855 6626
rect 45915 6620 45918 6626
rect 45895 6606 45918 6620
rect 45915 6600 45918 6606
rect 45944 6600 45947 6626
rect 46007 6620 46010 6626
rect 45987 6606 46010 6620
rect 46007 6600 46010 6606
rect 46036 6600 46039 6626
rect 44406 6572 45248 6586
rect 45271 6566 45274 6592
rect 45300 6586 45303 6592
rect 46568 6586 46582 6640
rect 47066 6638 47072 6640
rect 47089 6654 47095 6655
rect 47304 6654 47318 6674
rect 48998 6672 49004 6674
rect 49021 6672 49027 6689
rect 48998 6669 49027 6672
rect 49090 6689 49119 6692
rect 49090 6672 49096 6689
rect 49113 6688 49119 6689
rect 49549 6688 49552 6694
rect 49113 6674 49552 6688
rect 49113 6672 49119 6674
rect 49090 6669 49119 6672
rect 49549 6668 49552 6674
rect 49578 6668 49581 6694
rect 49673 6688 49687 6708
rect 50377 6702 50380 6728
rect 50406 6722 50409 6728
rect 50562 6723 50591 6726
rect 50562 6722 50568 6723
rect 50406 6708 50568 6722
rect 50406 6702 50409 6708
rect 50562 6706 50568 6708
rect 50585 6706 50591 6723
rect 50562 6703 50591 6706
rect 54517 6702 54520 6728
rect 54546 6722 54549 6728
rect 54702 6723 54731 6726
rect 54702 6722 54708 6723
rect 54546 6708 54708 6722
rect 54546 6702 54549 6708
rect 54702 6706 54708 6708
rect 54725 6706 54731 6723
rect 54702 6703 54731 6706
rect 55622 6723 55651 6726
rect 55622 6706 55628 6723
rect 55645 6722 55651 6723
rect 55851 6722 55854 6728
rect 55645 6708 55854 6722
rect 55645 6706 55651 6708
rect 55622 6703 55651 6706
rect 55851 6702 55854 6708
rect 55880 6702 55883 6728
rect 59439 6702 59442 6728
rect 59468 6722 59471 6728
rect 60635 6722 60638 6728
rect 59468 6708 60152 6722
rect 60615 6708 60638 6722
rect 59468 6702 59471 6708
rect 56128 6689 56157 6692
rect 56128 6688 56134 6689
rect 49673 6674 56134 6688
rect 56128 6672 56134 6674
rect 56151 6688 56157 6689
rect 56151 6674 57438 6688
rect 56151 6672 56157 6674
rect 56128 6669 56157 6672
rect 57424 6660 57438 6674
rect 59117 6668 59120 6694
rect 59146 6688 59149 6694
rect 60138 6692 60152 6708
rect 60635 6702 60638 6708
rect 60664 6702 60667 6728
rect 62061 6722 62064 6728
rect 62041 6708 62064 6722
rect 62061 6702 62064 6708
rect 62090 6702 62093 6728
rect 63763 6722 63766 6728
rect 63358 6708 63766 6722
rect 63358 6692 63372 6708
rect 63763 6702 63766 6708
rect 63792 6702 63795 6728
rect 68317 6722 68320 6728
rect 68297 6708 68320 6722
rect 68317 6702 68320 6708
rect 68346 6702 68349 6728
rect 69789 6702 69792 6728
rect 69818 6722 69821 6728
rect 70158 6723 70187 6726
rect 70158 6722 70164 6723
rect 69818 6708 70164 6722
rect 69818 6702 69821 6708
rect 70158 6706 70164 6708
rect 70181 6706 70187 6723
rect 71063 6722 71077 6742
rect 71445 6736 71448 6742
rect 71474 6736 71477 6762
rect 72366 6757 72395 6760
rect 72366 6740 72372 6757
rect 72389 6756 72395 6757
rect 72871 6756 72874 6762
rect 72389 6742 72874 6756
rect 72389 6740 72395 6742
rect 72366 6737 72395 6740
rect 72871 6736 72874 6742
rect 72900 6736 72903 6762
rect 74067 6756 74070 6762
rect 72926 6742 74070 6756
rect 72926 6722 72940 6742
rect 74067 6736 74070 6742
rect 74096 6736 74099 6762
rect 74154 6757 74183 6760
rect 74154 6740 74160 6757
rect 74177 6756 74183 6757
rect 75401 6756 75404 6762
rect 74177 6742 75404 6756
rect 74177 6740 74183 6742
rect 74154 6737 74183 6740
rect 75401 6736 75404 6742
rect 75430 6736 75433 6762
rect 78621 6756 78624 6762
rect 76100 6742 78624 6756
rect 71063 6708 72940 6722
rect 70158 6703 70187 6706
rect 60130 6689 60159 6692
rect 59146 6674 60106 6688
rect 59146 6668 59149 6674
rect 47089 6640 47318 6654
rect 48446 6655 48475 6658
rect 47089 6638 47095 6640
rect 47066 6635 47095 6638
rect 48446 6638 48452 6655
rect 48469 6654 48475 6655
rect 49688 6655 49717 6658
rect 48469 6640 48974 6654
rect 48469 6638 48475 6640
rect 48446 6635 48475 6638
rect 48353 6586 48356 6592
rect 45300 6572 46582 6586
rect 48333 6572 48356 6586
rect 45300 6566 45303 6572
rect 48353 6566 48356 6572
rect 48382 6566 48385 6592
rect 48767 6586 48770 6592
rect 48747 6572 48770 6586
rect 48767 6566 48770 6572
rect 48796 6566 48799 6592
rect 48960 6590 48974 6640
rect 49688 6638 49694 6655
rect 49711 6638 49717 6655
rect 49688 6635 49717 6638
rect 48997 6600 49000 6626
rect 49026 6620 49029 6626
rect 49595 6620 49598 6626
rect 49026 6606 49598 6620
rect 49026 6600 49029 6606
rect 49595 6600 49598 6606
rect 49624 6620 49627 6626
rect 49696 6620 49710 6635
rect 50699 6634 50702 6660
rect 50728 6654 50731 6660
rect 50976 6655 51005 6658
rect 50976 6654 50982 6655
rect 50728 6640 50982 6654
rect 50728 6634 50731 6640
rect 50976 6638 50982 6640
rect 50999 6638 51005 6655
rect 50976 6635 51005 6638
rect 49825 6620 49828 6626
rect 49624 6606 49710 6620
rect 49805 6606 49828 6620
rect 49624 6600 49627 6606
rect 49825 6600 49828 6606
rect 49854 6600 49857 6626
rect 50469 6620 50472 6626
rect 50439 6606 50472 6620
rect 50469 6600 50472 6606
rect 50498 6600 50501 6626
rect 48952 6587 48981 6590
rect 48952 6570 48958 6587
rect 48975 6586 48981 6587
rect 50515 6586 50518 6592
rect 48975 6572 50518 6586
rect 48975 6570 48981 6572
rect 48952 6567 48981 6570
rect 50515 6566 50518 6572
rect 50544 6566 50547 6592
rect 50984 6586 50998 6635
rect 51665 6634 51668 6660
rect 51694 6634 51697 6660
rect 52125 6654 52128 6660
rect 51766 6640 52128 6654
rect 51113 6620 51116 6626
rect 51093 6606 51116 6620
rect 51113 6600 51116 6606
rect 51142 6600 51145 6626
rect 51766 6586 51780 6640
rect 52125 6634 52128 6640
rect 52154 6634 52157 6660
rect 54793 6654 54796 6660
rect 54773 6640 54796 6654
rect 54793 6634 54796 6640
rect 54822 6634 54825 6660
rect 55713 6654 55716 6660
rect 55693 6640 55716 6654
rect 55713 6634 55716 6640
rect 55742 6634 55745 6660
rect 57415 6654 57418 6660
rect 57395 6640 57418 6654
rect 57415 6634 57418 6640
rect 57444 6634 57447 6660
rect 58703 6654 58706 6660
rect 58683 6640 58706 6654
rect 58703 6634 58706 6640
rect 58732 6634 58735 6660
rect 59393 6634 59396 6660
rect 59422 6634 59425 6660
rect 60092 6658 60106 6674
rect 60130 6672 60136 6689
rect 60153 6672 60159 6689
rect 60130 6669 60159 6672
rect 62844 6689 62873 6692
rect 62844 6672 62850 6689
rect 62867 6688 62873 6689
rect 63350 6689 63379 6692
rect 63350 6688 63356 6689
rect 62867 6674 63356 6688
rect 62867 6672 62873 6674
rect 62844 6669 62873 6672
rect 63350 6672 63356 6674
rect 63373 6672 63379 6689
rect 65143 6688 65146 6694
rect 63350 6669 63379 6672
rect 63772 6674 65146 6688
rect 63772 6660 63786 6674
rect 65143 6668 65146 6674
rect 65172 6688 65175 6694
rect 66294 6689 66323 6692
rect 66294 6688 66300 6689
rect 65172 6674 66300 6688
rect 65172 6668 65175 6674
rect 66294 6672 66300 6674
rect 66317 6688 66323 6689
rect 71031 6688 71034 6694
rect 66317 6674 71034 6688
rect 66317 6672 66323 6674
rect 66294 6669 66323 6672
rect 71031 6668 71034 6674
rect 71060 6668 71063 6694
rect 74022 6689 74051 6692
rect 72466 6674 73837 6688
rect 60084 6655 60113 6658
rect 60084 6638 60090 6655
rect 60107 6654 60113 6655
rect 60728 6655 60757 6658
rect 60728 6654 60734 6655
rect 60107 6640 60734 6654
rect 60107 6638 60113 6640
rect 60084 6635 60113 6638
rect 60728 6638 60734 6640
rect 60751 6638 60757 6655
rect 62154 6655 62183 6658
rect 62154 6654 62160 6655
rect 60728 6635 60757 6638
rect 61403 6640 62160 6654
rect 52033 6600 52036 6626
rect 52062 6620 52065 6626
rect 52264 6621 52293 6624
rect 52264 6620 52270 6621
rect 52062 6606 52270 6620
rect 52062 6600 52065 6606
rect 52264 6604 52270 6606
rect 52287 6604 52293 6621
rect 52264 6601 52293 6604
rect 52493 6600 52496 6626
rect 52522 6600 52525 6626
rect 56265 6620 56268 6626
rect 56245 6606 56268 6620
rect 56265 6600 56268 6606
rect 56294 6600 56297 6626
rect 57093 6620 57096 6626
rect 56879 6606 57096 6620
rect 57093 6600 57096 6606
rect 57122 6600 57125 6626
rect 57553 6620 57556 6626
rect 57533 6606 57556 6620
rect 57553 6600 57556 6606
rect 57582 6600 57585 6626
rect 58473 6620 58476 6626
rect 58167 6606 58476 6620
rect 58473 6600 58476 6606
rect 58502 6600 58505 6626
rect 58841 6620 58844 6626
rect 58821 6606 58844 6620
rect 58841 6600 58844 6606
rect 58870 6600 58873 6626
rect 60038 6621 60067 6624
rect 60038 6620 60044 6621
rect 59586 6606 60044 6620
rect 50984 6572 51780 6586
rect 51849 6566 51852 6592
rect 51878 6586 51881 6592
rect 52217 6586 52220 6592
rect 51878 6572 52220 6586
rect 51878 6566 51881 6572
rect 52217 6566 52220 6572
rect 52246 6566 52249 6592
rect 52309 6566 52312 6592
rect 52338 6586 52341 6592
rect 53000 6587 53029 6590
rect 53000 6586 53006 6587
rect 52338 6572 53006 6586
rect 52338 6566 52341 6572
rect 53000 6570 53006 6572
rect 53023 6586 53029 6587
rect 54793 6586 54796 6592
rect 53023 6572 54796 6586
rect 53023 6570 53029 6572
rect 53000 6567 53029 6570
rect 54793 6566 54796 6572
rect 54822 6566 54825 6592
rect 57002 6587 57031 6590
rect 57002 6570 57008 6587
rect 57025 6586 57031 6587
rect 57277 6586 57280 6592
rect 57025 6572 57280 6586
rect 57025 6570 57031 6572
rect 57002 6567 57031 6570
rect 57277 6566 57280 6572
rect 57306 6586 57309 6592
rect 57461 6586 57464 6592
rect 57306 6572 57464 6586
rect 57306 6566 57309 6572
rect 57461 6566 57464 6572
rect 57490 6566 57493 6592
rect 57875 6566 57878 6592
rect 57904 6586 57907 6592
rect 58290 6587 58319 6590
rect 58290 6586 58296 6587
rect 57904 6572 58296 6586
rect 57904 6566 57907 6572
rect 58290 6570 58296 6572
rect 58313 6586 58319 6587
rect 59025 6586 59028 6592
rect 58313 6572 59028 6586
rect 58313 6570 58319 6572
rect 58290 6567 58319 6570
rect 59025 6566 59028 6572
rect 59054 6566 59057 6592
rect 59586 6590 59600 6606
rect 60038 6604 60044 6606
rect 60061 6620 60067 6621
rect 61403 6620 61417 6640
rect 62154 6638 62160 6640
rect 62177 6654 62183 6655
rect 63304 6655 63333 6658
rect 63304 6654 63310 6655
rect 62177 6640 63310 6654
rect 62177 6638 62183 6640
rect 62154 6635 62183 6638
rect 63304 6638 63310 6640
rect 63327 6638 63333 6655
rect 63763 6654 63766 6660
rect 63743 6640 63766 6654
rect 63304 6635 63333 6638
rect 63763 6634 63766 6640
rect 63792 6634 63795 6660
rect 64683 6654 64686 6660
rect 64469 6640 64686 6654
rect 64683 6634 64686 6640
rect 64712 6634 64715 6660
rect 68409 6654 68412 6660
rect 68389 6640 68412 6654
rect 68409 6634 68412 6640
rect 68438 6634 68441 6660
rect 70250 6655 70279 6658
rect 70250 6638 70256 6655
rect 70273 6638 70279 6655
rect 71537 6654 71540 6660
rect 71517 6640 71540 6654
rect 70250 6635 70279 6638
rect 62751 6620 62754 6626
rect 60061 6606 61417 6620
rect 62731 6606 62754 6620
rect 60061 6604 60067 6606
rect 60038 6601 60067 6604
rect 62751 6600 62754 6606
rect 62780 6600 62783 6626
rect 63901 6620 63904 6626
rect 63881 6606 63904 6620
rect 63901 6600 63904 6606
rect 63930 6600 63933 6626
rect 65282 6621 65311 6624
rect 65282 6620 65288 6621
rect 64554 6606 65288 6620
rect 59578 6587 59607 6590
rect 59578 6570 59584 6587
rect 59601 6570 59607 6587
rect 59853 6586 59856 6592
rect 59833 6572 59856 6586
rect 59578 6567 59607 6570
rect 59853 6566 59856 6572
rect 59882 6566 59885 6592
rect 63073 6586 63076 6592
rect 63053 6572 63076 6586
rect 63073 6566 63076 6572
rect 63102 6566 63105 6592
rect 63257 6586 63260 6592
rect 63237 6572 63260 6586
rect 63257 6566 63260 6572
rect 63286 6566 63289 6592
rect 64039 6566 64042 6592
rect 64068 6586 64071 6592
rect 64554 6586 64568 6606
rect 65282 6604 65288 6606
rect 65305 6604 65311 6621
rect 65282 6601 65311 6604
rect 65603 6600 65606 6626
rect 65632 6600 65635 6626
rect 66431 6620 66434 6626
rect 66411 6606 66434 6620
rect 66431 6600 66434 6606
rect 66460 6600 66463 6626
rect 66661 6600 66664 6626
rect 66690 6600 66693 6626
rect 70258 6620 70272 6635
rect 71537 6634 71540 6640
rect 71566 6634 71569 6660
rect 72466 6658 72480 6674
rect 72458 6655 72487 6658
rect 72458 6638 72464 6655
rect 72481 6638 72487 6655
rect 72871 6654 72874 6660
rect 72851 6640 72874 6654
rect 72458 6635 72487 6638
rect 72871 6634 72874 6640
rect 72900 6634 72903 6660
rect 73823 6654 73837 6674
rect 74022 6672 74028 6689
rect 74045 6688 74051 6689
rect 75448 6689 75477 6692
rect 75448 6688 75454 6689
rect 74045 6674 75454 6688
rect 74045 6672 74051 6674
rect 74022 6669 74051 6672
rect 75448 6672 75454 6674
rect 75471 6688 75477 6689
rect 76100 6688 76114 6742
rect 78621 6736 78624 6742
rect 78650 6736 78653 6762
rect 78806 6757 78835 6760
rect 78806 6740 78812 6757
rect 78829 6756 78835 6757
rect 78989 6756 78992 6762
rect 78829 6742 78992 6756
rect 78829 6740 78835 6742
rect 78806 6737 78835 6740
rect 78989 6736 78992 6742
rect 79018 6736 79021 6762
rect 79725 6736 79728 6762
rect 79754 6756 79757 6762
rect 80783 6756 80786 6762
rect 79754 6742 80786 6756
rect 79754 6736 79757 6742
rect 80783 6736 80786 6742
rect 80812 6756 80815 6762
rect 81335 6756 81338 6762
rect 80812 6742 81338 6756
rect 80812 6736 80815 6742
rect 81335 6736 81338 6742
rect 81364 6736 81367 6762
rect 81749 6736 81752 6762
rect 81778 6756 81781 6762
rect 88189 6756 88192 6762
rect 81778 6742 88192 6756
rect 81778 6736 81781 6742
rect 88189 6736 88192 6742
rect 88218 6736 88221 6762
rect 91363 6756 91366 6762
rect 88244 6742 91294 6756
rect 91343 6742 91366 6756
rect 77471 6702 77474 6728
rect 77500 6722 77503 6728
rect 77886 6723 77915 6726
rect 77886 6722 77892 6723
rect 77500 6708 77892 6722
rect 77500 6702 77503 6708
rect 77886 6706 77892 6708
rect 77909 6706 77915 6723
rect 77886 6703 77915 6706
rect 83221 6702 83224 6728
rect 83250 6722 83253 6728
rect 85199 6722 85202 6728
rect 83250 6708 85130 6722
rect 85179 6708 85202 6722
rect 83250 6702 83253 6708
rect 75471 6674 76114 6688
rect 76736 6689 76765 6692
rect 75471 6672 75477 6674
rect 75448 6669 75477 6672
rect 76736 6672 76742 6689
rect 76759 6688 76765 6689
rect 80461 6688 80464 6694
rect 76759 6674 79334 6688
rect 80417 6674 80464 6688
rect 76759 6672 76765 6674
rect 76736 6669 76765 6672
rect 79320 6660 79334 6674
rect 80461 6668 80464 6674
rect 80490 6688 80493 6694
rect 80490 6674 82554 6688
rect 80490 6668 80493 6674
rect 82540 6662 82554 6674
rect 82623 6668 82626 6694
rect 82652 6688 82655 6694
rect 83314 6689 83343 6692
rect 83314 6688 83320 6689
rect 82652 6674 83320 6688
rect 82652 6668 82655 6674
rect 83314 6672 83320 6674
rect 83337 6688 83343 6689
rect 83774 6689 83803 6692
rect 83774 6688 83780 6689
rect 83337 6674 83780 6688
rect 83337 6672 83343 6674
rect 83314 6669 83343 6672
rect 83774 6672 83780 6674
rect 83797 6672 83803 6689
rect 83774 6669 83803 6672
rect 73823 6640 74044 6654
rect 72963 6620 72966 6626
rect 67176 6606 72966 6620
rect 64068 6572 64568 6586
rect 64068 6566 64071 6572
rect 64591 6566 64594 6592
rect 64620 6586 64623 6592
rect 64638 6587 64667 6590
rect 64638 6586 64644 6587
rect 64620 6572 64644 6586
rect 64620 6566 64623 6572
rect 64638 6570 64644 6572
rect 64661 6570 64667 6587
rect 64638 6567 64667 6570
rect 65787 6566 65790 6592
rect 65816 6586 65819 6592
rect 66018 6587 66047 6590
rect 66018 6586 66024 6587
rect 65816 6572 66024 6586
rect 65816 6566 65819 6572
rect 66018 6570 66024 6572
rect 66041 6586 66047 6587
rect 66845 6586 66848 6592
rect 66041 6572 66848 6586
rect 66041 6570 66047 6572
rect 66018 6567 66047 6570
rect 66845 6566 66848 6572
rect 66874 6566 66877 6592
rect 67075 6566 67078 6592
rect 67104 6586 67107 6592
rect 67176 6590 67190 6606
rect 72963 6600 72966 6606
rect 72992 6600 72995 6626
rect 73009 6600 73012 6626
rect 73038 6620 73041 6626
rect 73791 6620 73794 6626
rect 73038 6606 73060 6620
rect 73623 6606 73794 6620
rect 73038 6600 73041 6606
rect 73791 6600 73794 6606
rect 73820 6600 73823 6626
rect 67168 6587 67197 6590
rect 67168 6586 67174 6587
rect 67104 6572 67174 6586
rect 67104 6566 67107 6572
rect 67168 6570 67174 6572
rect 67191 6570 67197 6587
rect 67168 6567 67197 6570
rect 72917 6566 72920 6592
rect 72946 6586 72949 6592
rect 73745 6586 73748 6592
rect 72946 6572 73748 6586
rect 72946 6566 72949 6572
rect 73745 6566 73748 6572
rect 73774 6566 73777 6592
rect 74030 6586 74044 6640
rect 77609 6634 77612 6660
rect 77638 6654 77641 6660
rect 77931 6654 77934 6660
rect 77638 6640 77934 6654
rect 77638 6634 77641 6640
rect 77931 6634 77934 6640
rect 77960 6654 77963 6660
rect 77978 6655 78007 6658
rect 77978 6654 77984 6655
rect 77960 6640 77984 6654
rect 77960 6634 77963 6640
rect 77978 6638 77984 6640
rect 78001 6638 78007 6655
rect 78207 6654 78210 6660
rect 78187 6640 78210 6654
rect 77978 6635 78007 6638
rect 78207 6634 78210 6640
rect 78236 6634 78239 6660
rect 78897 6654 78900 6660
rect 78877 6640 78900 6654
rect 78897 6634 78900 6640
rect 78926 6634 78929 6660
rect 79311 6654 79314 6660
rect 79291 6640 79314 6654
rect 79311 6634 79314 6640
rect 79340 6634 79343 6660
rect 81335 6634 81338 6660
rect 81364 6654 81367 6660
rect 81749 6654 81752 6660
rect 81364 6640 81680 6654
rect 81729 6640 81752 6654
rect 81364 6634 81367 6640
rect 75034 6621 75063 6624
rect 74773 6606 75010 6620
rect 74619 6586 74622 6592
rect 74030 6572 74622 6586
rect 74619 6566 74622 6572
rect 74648 6566 74651 6592
rect 74996 6586 75010 6606
rect 75034 6604 75040 6621
rect 75057 6620 75063 6621
rect 75217 6620 75220 6626
rect 75057 6606 75220 6620
rect 75057 6604 75063 6606
rect 75034 6601 75063 6604
rect 75217 6600 75220 6606
rect 75246 6600 75249 6626
rect 75539 6600 75542 6626
rect 75568 6620 75571 6626
rect 75586 6621 75615 6624
rect 75586 6620 75592 6621
rect 75568 6606 75592 6620
rect 75568 6600 75571 6606
rect 75586 6604 75592 6606
rect 75609 6604 75615 6621
rect 76229 6620 76232 6626
rect 76199 6606 76232 6620
rect 75586 6601 75615 6604
rect 76229 6600 76232 6606
rect 76258 6600 76261 6626
rect 76873 6620 76876 6626
rect 76284 6606 76436 6620
rect 76853 6606 76876 6620
rect 76284 6586 76298 6606
rect 74996 6572 76298 6586
rect 76321 6566 76324 6592
rect 76350 6586 76353 6592
rect 76422 6586 76436 6606
rect 76873 6600 76876 6606
rect 76902 6600 76905 6626
rect 77103 6600 77106 6626
rect 77132 6600 77135 6626
rect 78254 6621 78283 6624
rect 78254 6620 78260 6621
rect 77526 6606 78260 6620
rect 77526 6586 77540 6606
rect 78254 6604 78260 6606
rect 78277 6604 78283 6621
rect 78254 6601 78283 6604
rect 78299 6600 78302 6626
rect 78328 6620 78331 6626
rect 79449 6620 79452 6626
rect 78328 6606 78667 6620
rect 79429 6606 79452 6620
rect 78328 6600 78331 6606
rect 77609 6586 77612 6592
rect 76350 6572 76372 6586
rect 76422 6572 77540 6586
rect 77589 6572 77612 6586
rect 76350 6566 76353 6572
rect 77609 6566 77612 6572
rect 77638 6566 77641 6592
rect 78653 6586 78667 6606
rect 79449 6600 79452 6606
rect 79478 6600 79481 6626
rect 80599 6620 80602 6626
rect 80063 6606 80346 6620
rect 80579 6606 80602 6620
rect 79771 6586 79774 6592
rect 78653 6572 79774 6586
rect 79771 6566 79774 6572
rect 79800 6566 79803 6592
rect 80185 6586 80188 6592
rect 80165 6572 80188 6586
rect 80185 6566 80188 6572
rect 80214 6566 80217 6592
rect 80332 6586 80346 6606
rect 80599 6600 80602 6606
rect 80628 6600 80631 6626
rect 81381 6620 81384 6626
rect 81213 6606 81384 6620
rect 81381 6600 81384 6606
rect 81410 6600 81413 6626
rect 81013 6586 81016 6592
rect 80332 6572 81016 6586
rect 81013 6566 81016 6572
rect 81042 6566 81045 6592
rect 81243 6566 81246 6592
rect 81272 6586 81275 6592
rect 81336 6587 81365 6590
rect 81336 6586 81342 6587
rect 81272 6572 81342 6586
rect 81272 6566 81275 6572
rect 81336 6570 81342 6572
rect 81359 6570 81365 6587
rect 81666 6586 81680 6640
rect 81749 6634 81752 6640
rect 81778 6634 81781 6660
rect 82439 6634 82442 6660
rect 82468 6634 82471 6660
rect 82540 6654 82600 6662
rect 85116 6654 85130 6708
rect 85199 6702 85202 6708
rect 85228 6702 85231 6728
rect 86533 6722 86536 6728
rect 86513 6708 86536 6722
rect 86533 6702 86536 6708
rect 86562 6702 86565 6728
rect 86901 6722 86904 6728
rect 86881 6708 86904 6722
rect 86901 6702 86904 6708
rect 86930 6702 86933 6728
rect 87914 6723 87943 6726
rect 87914 6722 87920 6723
rect 87186 6708 87920 6722
rect 87186 6692 87200 6708
rect 87914 6706 87920 6708
rect 87937 6722 87943 6723
rect 87959 6722 87962 6728
rect 87937 6708 87962 6722
rect 87937 6706 87943 6708
rect 87914 6703 87943 6706
rect 87959 6702 87962 6708
rect 87988 6702 87991 6728
rect 88005 6702 88008 6728
rect 88034 6722 88037 6728
rect 88244 6722 88258 6742
rect 88034 6708 88258 6722
rect 88034 6702 88037 6708
rect 88879 6702 88882 6728
rect 88908 6722 88911 6728
rect 89064 6723 89093 6726
rect 89064 6722 89070 6723
rect 88908 6708 89070 6722
rect 88908 6702 88911 6708
rect 89064 6706 89070 6708
rect 89087 6706 89093 6723
rect 89064 6703 89093 6706
rect 90213 6702 90216 6728
rect 90242 6722 90245 6728
rect 90766 6723 90795 6726
rect 90766 6722 90772 6723
rect 90242 6708 90772 6722
rect 90242 6702 90245 6708
rect 90766 6706 90772 6708
rect 90789 6706 90795 6723
rect 90766 6703 90795 6706
rect 87132 6689 87161 6692
rect 87132 6688 87138 6689
rect 85300 6674 87138 6688
rect 85300 6658 85314 6674
rect 87132 6672 87138 6674
rect 87155 6672 87161 6689
rect 87132 6669 87161 6672
rect 87178 6689 87207 6692
rect 87178 6672 87184 6689
rect 87201 6672 87207 6689
rect 89478 6689 89507 6692
rect 89478 6688 89484 6689
rect 87178 6669 87207 6672
rect 87232 6674 87982 6688
rect 85292 6655 85321 6658
rect 85292 6654 85298 6655
rect 82540 6648 85084 6654
rect 82586 6640 85084 6648
rect 85116 6640 85298 6654
rect 81887 6620 81890 6626
rect 81867 6606 81890 6620
rect 81887 6600 81890 6606
rect 81916 6600 81919 6626
rect 82577 6620 82580 6626
rect 82540 6606 82580 6620
rect 82301 6586 82304 6592
rect 81666 6572 82304 6586
rect 81336 6567 81365 6570
rect 82301 6566 82304 6572
rect 82330 6586 82333 6592
rect 82540 6586 82554 6606
rect 82577 6600 82580 6606
rect 82606 6600 82609 6626
rect 83268 6621 83297 6624
rect 83268 6620 83274 6621
rect 82632 6606 83274 6620
rect 82632 6592 82646 6606
rect 83268 6604 83274 6606
rect 83291 6604 83297 6621
rect 83681 6620 83684 6626
rect 83637 6606 83684 6620
rect 83268 6601 83297 6604
rect 83681 6600 83684 6606
rect 83710 6600 83713 6626
rect 85070 6620 85084 6640
rect 85292 6638 85298 6640
rect 85315 6638 85321 6655
rect 85292 6635 85321 6638
rect 86626 6655 86655 6658
rect 86626 6638 86632 6655
rect 86649 6654 86655 6655
rect 87085 6654 87088 6660
rect 86649 6640 87088 6654
rect 86649 6638 86655 6640
rect 86626 6635 86655 6638
rect 87085 6634 87088 6640
rect 87114 6634 87117 6660
rect 87232 6620 87246 6674
rect 87822 6655 87851 6658
rect 87822 6654 87828 6655
rect 85070 6606 87246 6620
rect 87278 6640 87828 6654
rect 82623 6586 82626 6592
rect 82330 6572 82554 6586
rect 82603 6572 82626 6586
rect 82330 6566 82333 6572
rect 82623 6566 82626 6572
rect 82652 6566 82655 6592
rect 82669 6566 82672 6592
rect 82698 6586 82701 6592
rect 83038 6587 83067 6590
rect 83038 6586 83044 6587
rect 82698 6572 83044 6586
rect 82698 6566 82701 6572
rect 83038 6570 83044 6572
rect 83061 6570 83067 6587
rect 83221 6586 83224 6592
rect 83201 6572 83224 6586
rect 83038 6567 83067 6570
rect 83221 6566 83224 6572
rect 83250 6566 83253 6592
rect 83690 6586 83704 6600
rect 87278 6586 87292 6640
rect 87822 6638 87828 6640
rect 87845 6654 87851 6655
rect 87913 6654 87916 6660
rect 87845 6640 87916 6654
rect 87845 6638 87851 6640
rect 87822 6635 87851 6638
rect 87913 6634 87916 6640
rect 87942 6634 87945 6660
rect 87968 6652 87982 6674
rect 88060 6674 89484 6688
rect 88060 6652 88074 6674
rect 89478 6672 89484 6674
rect 89501 6688 89507 6689
rect 90949 6688 90952 6694
rect 89501 6674 90952 6688
rect 89501 6672 89507 6674
rect 89478 6669 89507 6672
rect 90949 6668 90952 6674
rect 90978 6668 90981 6694
rect 91041 6668 91044 6694
rect 91070 6688 91073 6694
rect 91280 6688 91294 6742
rect 91363 6736 91366 6742
rect 91392 6736 91395 6762
rect 92881 6756 92884 6762
rect 92861 6742 92884 6756
rect 92881 6736 92884 6742
rect 92910 6736 92913 6762
rect 94675 6756 94678 6762
rect 92936 6742 94678 6756
rect 92936 6688 92950 6742
rect 94675 6736 94678 6742
rect 94704 6736 94707 6762
rect 94730 6742 95434 6756
rect 94399 6702 94402 6728
rect 94428 6722 94431 6728
rect 94730 6722 94744 6742
rect 94428 6708 94744 6722
rect 94428 6702 94431 6708
rect 94767 6702 94770 6728
rect 94796 6722 94799 6728
rect 95420 6722 95434 6742
rect 95457 6736 95460 6762
rect 95486 6756 95489 6762
rect 96745 6756 96748 6762
rect 95486 6742 96748 6756
rect 95486 6736 95489 6742
rect 96745 6736 96748 6742
rect 96774 6736 96777 6762
rect 103553 6756 103556 6762
rect 98686 6742 103556 6756
rect 95917 6722 95920 6728
rect 94796 6708 94836 6722
rect 95420 6708 95920 6722
rect 94796 6702 94799 6708
rect 94261 6688 94264 6694
rect 91070 6674 91092 6688
rect 91280 6674 92950 6688
rect 92982 6674 93732 6688
rect 94241 6674 94264 6688
rect 91070 6668 91073 6674
rect 88189 6654 88192 6660
rect 87968 6638 88074 6652
rect 88169 6640 88192 6654
rect 88189 6634 88192 6640
rect 88218 6634 88221 6660
rect 90305 6634 90308 6660
rect 90334 6654 90337 6660
rect 92982 6658 92996 6674
rect 90996 6655 91025 6658
rect 90996 6654 91002 6655
rect 90334 6640 91002 6654
rect 90334 6634 90337 6640
rect 90996 6638 91002 6640
rect 91019 6654 91025 6655
rect 91456 6655 91485 6658
rect 91456 6654 91462 6655
rect 91019 6640 91462 6654
rect 91019 6638 91025 6640
rect 90996 6635 91025 6638
rect 91456 6638 91462 6640
rect 91479 6638 91485 6655
rect 91456 6635 91485 6638
rect 92974 6655 93003 6658
rect 92974 6638 92980 6655
rect 92997 6638 93003 6655
rect 92974 6635 93003 6638
rect 93664 6655 93693 6658
rect 93664 6638 93670 6655
rect 93687 6638 93693 6655
rect 93718 6654 93732 6674
rect 94261 6668 94264 6674
rect 94290 6668 94293 6694
rect 94822 6688 94836 6708
rect 95917 6702 95920 6708
rect 95946 6702 95949 6728
rect 98686 6722 98700 6742
rect 103553 6736 103556 6742
rect 103582 6736 103585 6762
rect 105163 6756 105166 6762
rect 103608 6742 103990 6756
rect 105143 6742 105166 6756
rect 97858 6708 98700 6722
rect 99920 6723 99949 6726
rect 94906 6689 94935 6692
rect 94906 6688 94912 6689
rect 94822 6674 94912 6688
rect 94906 6672 94912 6674
rect 94929 6672 94935 6689
rect 94906 6669 94935 6672
rect 94951 6668 94954 6694
rect 94980 6688 94983 6694
rect 97858 6688 97872 6708
rect 99920 6706 99926 6723
rect 99943 6722 99949 6723
rect 100977 6722 100980 6728
rect 99943 6708 100980 6722
rect 99943 6706 99949 6708
rect 99920 6703 99949 6706
rect 100977 6702 100980 6708
rect 101006 6702 101009 6728
rect 101713 6702 101716 6728
rect 101742 6722 101745 6728
rect 101944 6723 101973 6726
rect 101944 6722 101950 6723
rect 101742 6708 101950 6722
rect 101742 6702 101745 6708
rect 101944 6706 101950 6708
rect 101967 6706 101973 6723
rect 101944 6703 101973 6706
rect 103001 6702 103004 6728
rect 103030 6722 103033 6728
rect 103608 6722 103622 6742
rect 103030 6708 103622 6722
rect 103030 6702 103033 6708
rect 103875 6702 103878 6728
rect 103904 6722 103907 6728
rect 103904 6708 103944 6722
rect 103904 6702 103907 6708
rect 94980 6674 97872 6688
rect 94980 6668 94983 6674
rect 98815 6668 98818 6694
rect 98844 6688 98847 6694
rect 99368 6689 99397 6692
rect 99368 6688 99374 6689
rect 98844 6674 99374 6688
rect 98844 6668 98847 6674
rect 99368 6672 99374 6674
rect 99391 6672 99397 6689
rect 99368 6669 99397 6672
rect 100564 6689 100593 6692
rect 100564 6672 100570 6689
rect 100587 6688 100593 6689
rect 101023 6688 101026 6694
rect 100587 6674 101026 6688
rect 100587 6672 100593 6674
rect 100564 6669 100593 6672
rect 101023 6668 101026 6674
rect 101052 6668 101055 6694
rect 103930 6692 103944 6708
rect 102358 6689 102387 6692
rect 102358 6688 102364 6689
rect 101078 6674 102364 6688
rect 101078 6660 101092 6674
rect 102358 6672 102364 6674
rect 102381 6688 102387 6689
rect 103922 6689 103951 6692
rect 102381 6674 103898 6688
rect 102381 6672 102387 6674
rect 102358 6669 102387 6672
rect 94216 6655 94245 6658
rect 94216 6654 94222 6655
rect 93718 6640 94222 6654
rect 93664 6635 93693 6638
rect 94216 6638 94222 6640
rect 94239 6638 94245 6655
rect 94767 6654 94770 6660
rect 94747 6640 94770 6654
rect 94216 6635 94245 6638
rect 87867 6600 87870 6626
rect 87896 6620 87899 6626
rect 88328 6621 88357 6624
rect 88328 6620 88334 6621
rect 87896 6606 88334 6620
rect 87896 6600 87899 6606
rect 88328 6604 88334 6606
rect 88351 6604 88357 6621
rect 88328 6601 88357 6604
rect 88833 6600 88836 6626
rect 88862 6600 88865 6626
rect 89616 6621 89645 6624
rect 89616 6620 89622 6621
rect 88980 6606 89622 6620
rect 83690 6572 87292 6586
rect 87499 6566 87502 6592
rect 87528 6586 87531 6592
rect 88980 6586 88994 6606
rect 89616 6604 89622 6606
rect 89639 6604 89645 6621
rect 89616 6601 89645 6604
rect 89983 6600 89986 6626
rect 90012 6600 90015 6626
rect 90443 6600 90446 6626
rect 90472 6620 90475 6626
rect 90950 6621 90979 6624
rect 90950 6620 90956 6621
rect 90472 6606 90956 6620
rect 90472 6600 90475 6606
rect 90950 6604 90956 6606
rect 90973 6620 90979 6621
rect 92982 6620 92996 6635
rect 90973 6606 92996 6620
rect 90973 6604 90979 6606
rect 90950 6601 90979 6604
rect 90351 6586 90354 6592
rect 87528 6572 88994 6586
rect 90331 6572 90354 6586
rect 87528 6566 87531 6572
rect 90351 6566 90354 6572
rect 90380 6566 90383 6592
rect 93672 6586 93686 6635
rect 94767 6634 94770 6640
rect 94796 6634 94799 6660
rect 95918 6655 95947 6658
rect 95918 6638 95924 6655
rect 95941 6638 95947 6655
rect 95918 6635 95947 6638
rect 97206 6655 97235 6658
rect 97206 6638 97212 6655
rect 97229 6638 97235 6655
rect 97206 6635 97235 6638
rect 100012 6655 100041 6658
rect 100012 6638 100018 6655
rect 100035 6654 100041 6655
rect 100747 6654 100750 6660
rect 100035 6640 100750 6654
rect 100035 6638 100041 6640
rect 100012 6635 100041 6638
rect 93710 6621 93739 6624
rect 93710 6604 93716 6621
rect 93733 6620 93739 6621
rect 95926 6620 95940 6635
rect 93733 6606 95151 6620
rect 95604 6606 95940 6620
rect 93733 6604 93739 6606
rect 93710 6601 93739 6604
rect 93893 6586 93896 6592
rect 93672 6572 93896 6586
rect 93893 6566 93896 6572
rect 93922 6566 93925 6592
rect 93985 6586 93988 6592
rect 93965 6572 93988 6586
rect 93985 6566 93988 6572
rect 94014 6566 94017 6592
rect 94169 6586 94172 6592
rect 94149 6572 94172 6586
rect 94169 6566 94172 6572
rect 94198 6566 94201 6592
rect 94767 6566 94770 6592
rect 94796 6586 94799 6592
rect 95604 6586 95618 6606
rect 94796 6572 95618 6586
rect 95642 6587 95671 6590
rect 94796 6566 94799 6572
rect 95642 6570 95648 6587
rect 95665 6586 95671 6587
rect 95687 6586 95690 6592
rect 95665 6572 95690 6586
rect 95665 6570 95671 6572
rect 95642 6567 95671 6570
rect 95687 6566 95690 6572
rect 95716 6566 95719 6592
rect 95926 6586 95940 6606
rect 96056 6621 96085 6624
rect 96056 6604 96062 6621
rect 96079 6620 96085 6621
rect 96193 6620 96196 6626
rect 96079 6606 96196 6620
rect 96079 6604 96085 6606
rect 96056 6601 96085 6604
rect 96193 6600 96196 6606
rect 96222 6600 96225 6626
rect 96699 6620 96702 6626
rect 96669 6606 96702 6620
rect 96699 6600 96702 6606
rect 96728 6600 96731 6626
rect 96930 6621 96959 6624
rect 96930 6604 96936 6621
rect 96953 6620 96959 6621
rect 96975 6620 96978 6626
rect 96953 6606 96978 6620
rect 96953 6604 96959 6606
rect 96930 6601 96959 6604
rect 96975 6600 96978 6606
rect 97004 6600 97007 6626
rect 97214 6586 97228 6635
rect 100747 6634 100750 6640
rect 100776 6634 100779 6660
rect 101069 6654 101072 6660
rect 101049 6640 101072 6654
rect 101069 6634 101072 6640
rect 101098 6634 101101 6660
rect 103599 6654 103602 6660
rect 103148 6640 103602 6654
rect 97297 6600 97300 6626
rect 97326 6620 97329 6626
rect 97344 6621 97373 6624
rect 97344 6620 97350 6621
rect 97326 6606 97350 6620
rect 97326 6600 97329 6606
rect 97344 6604 97350 6606
rect 97367 6604 97373 6621
rect 97344 6601 97373 6604
rect 97389 6600 97392 6626
rect 97418 6620 97421 6626
rect 98217 6620 98220 6626
rect 97418 6606 97589 6620
rect 98173 6606 98220 6620
rect 97418 6600 97421 6606
rect 98217 6600 98220 6606
rect 98246 6620 98249 6626
rect 98677 6620 98680 6626
rect 98246 6606 98680 6620
rect 98246 6600 98249 6606
rect 98677 6600 98680 6606
rect 98706 6600 98709 6626
rect 98908 6621 98937 6624
rect 98908 6604 98914 6621
rect 98931 6620 98937 6621
rect 99322 6621 99351 6624
rect 98931 6606 99298 6620
rect 98931 6604 98937 6606
rect 98908 6601 98937 6604
rect 99284 6592 99298 6606
rect 99322 6604 99328 6621
rect 99345 6620 99351 6621
rect 101207 6620 101210 6626
rect 99345 6606 101092 6620
rect 101187 6606 101210 6620
rect 99345 6604 99351 6606
rect 99322 6601 99351 6604
rect 98861 6586 98864 6592
rect 95926 6572 98864 6586
rect 98861 6566 98864 6572
rect 98890 6566 98893 6592
rect 98953 6566 98956 6592
rect 98982 6586 98985 6592
rect 99092 6587 99121 6590
rect 99092 6586 99098 6587
rect 98982 6572 99098 6586
rect 98982 6566 98985 6572
rect 99092 6570 99098 6572
rect 99115 6570 99121 6587
rect 99275 6586 99278 6592
rect 99255 6572 99278 6586
rect 99092 6567 99121 6570
rect 99275 6566 99278 6572
rect 99304 6566 99307 6592
rect 100241 6586 100244 6592
rect 100221 6572 100244 6586
rect 100241 6566 100244 6572
rect 100270 6566 100273 6592
rect 100425 6586 100428 6592
rect 100405 6572 100428 6586
rect 100425 6566 100428 6572
rect 100454 6566 100457 6592
rect 100472 6587 100501 6590
rect 100472 6570 100478 6587
rect 100495 6586 100501 6587
rect 100655 6586 100658 6592
rect 100495 6572 100658 6586
rect 100495 6570 100501 6572
rect 100472 6567 100501 6570
rect 100655 6566 100658 6572
rect 100684 6566 100687 6592
rect 101078 6586 101092 6606
rect 101207 6600 101210 6606
rect 101236 6600 101239 6626
rect 101575 6600 101578 6626
rect 101604 6600 101607 6626
rect 101906 6606 102012 6620
rect 101906 6586 101920 6606
rect 101078 6572 101920 6586
rect 101998 6586 102012 6606
rect 102127 6600 102130 6626
rect 102156 6620 102159 6626
rect 102496 6621 102525 6624
rect 102496 6620 102502 6621
rect 102156 6606 102502 6620
rect 102156 6600 102159 6606
rect 102496 6604 102502 6606
rect 102519 6604 102525 6621
rect 102496 6601 102525 6604
rect 102725 6600 102728 6626
rect 102754 6600 102757 6626
rect 102817 6586 102820 6592
rect 101998 6572 102820 6586
rect 102817 6566 102820 6572
rect 102846 6566 102849 6592
rect 102863 6566 102866 6592
rect 102892 6586 102895 6592
rect 103148 6586 103162 6640
rect 103599 6634 103602 6640
rect 103628 6634 103631 6660
rect 103830 6655 103859 6658
rect 103830 6654 103836 6655
rect 103792 6640 103836 6654
rect 103792 6626 103806 6640
rect 103830 6638 103836 6640
rect 103853 6638 103859 6655
rect 103830 6635 103859 6638
rect 103185 6600 103188 6626
rect 103214 6620 103217 6626
rect 103214 6606 103438 6620
rect 103214 6600 103217 6606
rect 103232 6587 103261 6590
rect 103232 6586 103238 6587
rect 102892 6572 103238 6586
rect 102892 6566 102895 6572
rect 103232 6570 103238 6572
rect 103255 6570 103261 6587
rect 103424 6586 103438 6606
rect 103783 6600 103786 6626
rect 103812 6600 103815 6626
rect 103884 6620 103898 6674
rect 103922 6672 103928 6689
rect 103945 6672 103951 6689
rect 103976 6688 103990 6742
rect 105163 6736 105166 6742
rect 105192 6736 105195 6762
rect 106681 6756 106684 6762
rect 106661 6742 106684 6756
rect 106681 6736 106684 6742
rect 106710 6736 106713 6762
rect 134465 6756 134468 6762
rect 106736 6742 134468 6756
rect 104013 6702 104016 6728
rect 104042 6722 104045 6728
rect 106635 6722 106638 6728
rect 104042 6708 106638 6722
rect 104042 6702 104045 6708
rect 106635 6702 106638 6708
rect 106664 6702 106667 6728
rect 106736 6688 106750 6742
rect 134465 6736 134468 6742
rect 134494 6736 134497 6762
rect 134690 6757 134719 6760
rect 134690 6740 134696 6757
rect 134713 6756 134719 6757
rect 134787 6756 134790 6762
rect 134713 6742 134790 6756
rect 134713 6740 134719 6742
rect 134690 6737 134719 6740
rect 134787 6736 134790 6742
rect 134816 6736 134819 6762
rect 135891 6736 135894 6762
rect 135920 6756 135923 6762
rect 137134 6757 137163 6760
rect 137134 6756 137140 6757
rect 135920 6742 137140 6756
rect 135920 6736 135923 6742
rect 137134 6740 137140 6742
rect 137157 6740 137163 6757
rect 137455 6756 137458 6762
rect 137435 6742 137458 6756
rect 137134 6737 137163 6740
rect 137455 6736 137458 6742
rect 137484 6736 137487 6762
rect 138927 6756 138930 6762
rect 138907 6742 138930 6756
rect 138927 6736 138930 6742
rect 138956 6736 138959 6762
rect 140445 6756 140448 6762
rect 140425 6742 140448 6756
rect 140445 6736 140448 6742
rect 140474 6736 140477 6762
rect 142147 6736 142150 6762
rect 142176 6756 142179 6762
rect 142286 6757 142315 6760
rect 142286 6756 142292 6757
rect 142176 6742 142292 6756
rect 142176 6736 142179 6742
rect 142286 6740 142292 6742
rect 142309 6740 142315 6757
rect 142286 6737 142315 6740
rect 143527 6736 143530 6762
rect 143556 6756 143559 6762
rect 143574 6757 143603 6760
rect 143574 6756 143580 6757
rect 143556 6742 143580 6756
rect 143556 6736 143559 6742
rect 143574 6740 143580 6742
rect 143597 6740 143603 6757
rect 145045 6756 145048 6762
rect 145025 6742 145048 6756
rect 143574 6737 143603 6740
rect 145045 6736 145048 6742
rect 145074 6736 145077 6762
rect 146609 6756 146612 6762
rect 146589 6742 146612 6756
rect 146609 6736 146612 6742
rect 146638 6736 146641 6762
rect 148127 6756 148130 6762
rect 148107 6742 148130 6756
rect 148127 6736 148130 6742
rect 148156 6736 148159 6762
rect 149645 6756 149648 6762
rect 149625 6742 149648 6756
rect 149645 6736 149648 6742
rect 149674 6736 149677 6762
rect 150703 6756 150706 6762
rect 150683 6742 150706 6756
rect 150703 6736 150706 6742
rect 150732 6756 150735 6762
rect 150888 6757 150917 6760
rect 150888 6756 150894 6757
rect 150732 6742 150894 6756
rect 150732 6736 150735 6742
rect 150888 6740 150894 6742
rect 150911 6756 150917 6757
rect 151072 6757 151101 6760
rect 151072 6756 151078 6757
rect 150911 6742 151078 6756
rect 150911 6740 150917 6742
rect 150888 6737 150917 6740
rect 151072 6740 151078 6742
rect 151095 6756 151101 6757
rect 151486 6757 151515 6760
rect 151486 6756 151492 6757
rect 151095 6742 151492 6756
rect 151095 6740 151101 6742
rect 151072 6737 151101 6740
rect 151486 6740 151492 6742
rect 151509 6756 151515 6757
rect 151670 6757 151699 6760
rect 151670 6756 151676 6757
rect 151509 6742 151676 6756
rect 151509 6740 151515 6742
rect 151486 6737 151515 6740
rect 151670 6740 151676 6742
rect 151693 6740 151699 6757
rect 151670 6737 151699 6740
rect 108199 6722 108202 6728
rect 108179 6708 108202 6722
rect 108199 6702 108202 6708
rect 108228 6702 108231 6728
rect 109717 6702 109720 6728
rect 109746 6722 109749 6728
rect 110086 6723 110115 6726
rect 110086 6722 110092 6723
rect 109746 6708 110092 6722
rect 109746 6702 109749 6708
rect 110086 6706 110092 6708
rect 110109 6706 110115 6723
rect 112063 6722 112066 6728
rect 110086 6703 110115 6706
rect 110140 6708 112066 6722
rect 103976 6674 106750 6688
rect 103922 6669 103951 6672
rect 103967 6634 103970 6660
rect 103996 6654 103999 6660
rect 105256 6655 105285 6658
rect 105256 6654 105262 6655
rect 103996 6640 105262 6654
rect 103996 6634 103999 6640
rect 105256 6638 105262 6640
rect 105279 6638 105285 6655
rect 106773 6654 106776 6660
rect 106753 6640 106776 6654
rect 105256 6635 105285 6638
rect 106773 6634 106776 6640
rect 106802 6634 106805 6660
rect 108291 6654 108294 6660
rect 108247 6640 108294 6654
rect 108291 6634 108294 6640
rect 108320 6654 108323 6660
rect 110140 6654 110154 6708
rect 112063 6702 112066 6708
rect 112092 6702 112095 6728
rect 113213 6722 113216 6728
rect 112164 6708 113216 6722
rect 112017 6688 112020 6694
rect 110186 6674 112020 6688
rect 110186 6658 110200 6674
rect 112017 6668 112020 6674
rect 112046 6668 112049 6694
rect 112164 6692 112178 6708
rect 113213 6702 113216 6708
rect 113242 6702 113245 6728
rect 113305 6702 113308 6728
rect 113334 6722 113337 6728
rect 113334 6708 113356 6722
rect 113334 6702 113337 6708
rect 113443 6702 113446 6728
rect 113472 6722 113475 6728
rect 113949 6722 113952 6728
rect 113472 6708 113952 6722
rect 113472 6702 113475 6708
rect 113949 6702 113952 6708
rect 113978 6702 113981 6728
rect 114593 6702 114596 6728
rect 114622 6722 114625 6728
rect 114824 6723 114853 6726
rect 114824 6722 114830 6723
rect 114622 6708 114830 6722
rect 114622 6702 114625 6708
rect 114824 6706 114830 6708
rect 114847 6706 114853 6723
rect 114824 6703 114853 6706
rect 115890 6708 119170 6722
rect 112156 6689 112185 6692
rect 112156 6672 112162 6689
rect 112179 6672 112185 6689
rect 112156 6669 112185 6672
rect 112201 6668 112204 6694
rect 112230 6688 112233 6694
rect 113535 6688 113538 6694
rect 112230 6674 113538 6688
rect 112230 6668 112233 6674
rect 113535 6668 113538 6674
rect 113564 6668 113567 6694
rect 113581 6668 113584 6694
rect 113610 6688 113613 6694
rect 115238 6689 115267 6692
rect 115238 6688 115244 6689
rect 113610 6674 113632 6688
rect 113912 6674 115244 6688
rect 113610 6668 113613 6674
rect 108320 6640 110154 6654
rect 110178 6655 110207 6658
rect 108320 6634 108323 6640
rect 110178 6638 110184 6655
rect 110201 6638 110207 6655
rect 110178 6635 110207 6638
rect 111466 6655 111495 6658
rect 111466 6638 111472 6655
rect 111489 6654 111495 6655
rect 112938 6655 112967 6658
rect 112808 6654 112868 6655
rect 111489 6640 112178 6654
rect 111489 6638 111495 6640
rect 111466 6635 111495 6638
rect 112109 6620 112112 6626
rect 103884 6606 112112 6620
rect 112109 6600 112112 6606
rect 112138 6600 112141 6626
rect 103646 6587 103675 6590
rect 103646 6586 103652 6587
rect 103424 6572 103652 6586
rect 103232 6567 103261 6570
rect 103646 6570 103652 6572
rect 103669 6570 103675 6587
rect 103646 6567 103675 6570
rect 103691 6566 103694 6592
rect 103720 6586 103723 6592
rect 103876 6587 103905 6590
rect 103876 6586 103882 6587
rect 103720 6572 103882 6586
rect 103720 6566 103723 6572
rect 103876 6570 103882 6572
rect 103899 6586 103905 6587
rect 106773 6586 106776 6592
rect 103899 6572 106776 6586
rect 103899 6570 103905 6572
rect 103876 6567 103905 6570
rect 106773 6566 106776 6572
rect 106802 6566 106805 6592
rect 111373 6586 111376 6592
rect 111353 6572 111376 6586
rect 111373 6566 111376 6572
rect 111402 6566 111405 6592
rect 111833 6586 111836 6592
rect 111813 6572 111836 6586
rect 111833 6566 111836 6572
rect 111862 6566 111865 6592
rect 112017 6586 112020 6592
rect 111997 6572 112020 6586
rect 112017 6566 112020 6572
rect 112046 6566 112049 6592
rect 112063 6566 112066 6592
rect 112092 6586 112095 6592
rect 112164 6586 112178 6640
rect 112716 6641 112914 6654
rect 112716 6640 112822 6641
rect 112854 6640 112914 6641
rect 112201 6600 112204 6626
rect 112230 6620 112233 6626
rect 112716 6620 112730 6640
rect 112230 6606 112730 6620
rect 112900 6620 112914 6640
rect 112938 6638 112944 6655
rect 112961 6654 112967 6655
rect 113857 6654 113860 6660
rect 112961 6640 113860 6654
rect 112961 6638 112967 6640
rect 112938 6635 112967 6638
rect 113857 6634 113860 6640
rect 113886 6634 113889 6660
rect 113912 6620 113926 6674
rect 115238 6672 115244 6674
rect 115261 6688 115267 6689
rect 115890 6688 115904 6708
rect 115261 6674 115904 6688
rect 115261 6672 115267 6674
rect 115238 6669 115267 6672
rect 115973 6668 115976 6694
rect 116002 6688 116005 6694
rect 116112 6689 116141 6692
rect 116112 6688 116118 6689
rect 116002 6674 116118 6688
rect 116002 6668 116005 6674
rect 116112 6672 116118 6674
rect 116135 6672 116141 6689
rect 116571 6688 116574 6694
rect 116112 6669 116141 6672
rect 116350 6674 116574 6688
rect 113950 6655 113979 6658
rect 113950 6638 113956 6655
rect 113973 6638 113979 6655
rect 115191 6654 115194 6660
rect 114655 6640 115194 6654
rect 113950 6635 113979 6638
rect 112900 6606 113926 6620
rect 112230 6600 112233 6606
rect 113958 6592 113972 6635
rect 115191 6634 115194 6640
rect 115220 6634 115223 6660
rect 115927 6634 115930 6660
rect 115956 6634 115959 6660
rect 116019 6634 116022 6660
rect 116048 6654 116051 6660
rect 116350 6654 116364 6674
rect 116571 6668 116574 6674
rect 116600 6668 116603 6694
rect 116663 6668 116666 6694
rect 116692 6688 116695 6694
rect 118596 6689 118625 6692
rect 118596 6688 118602 6689
rect 116692 6674 118602 6688
rect 116692 6668 116695 6674
rect 116525 6654 116528 6660
rect 116048 6640 116364 6654
rect 116505 6640 116528 6654
rect 116048 6634 116051 6640
rect 116525 6634 116528 6640
rect 116554 6634 116557 6660
rect 116940 6655 116969 6658
rect 116580 6642 116870 6654
rect 116580 6640 116916 6642
rect 114041 6600 114044 6626
rect 114070 6620 114073 6626
rect 114088 6621 114117 6624
rect 114088 6620 114094 6621
rect 114070 6606 114094 6620
rect 114070 6600 114073 6606
rect 114088 6604 114094 6606
rect 114111 6604 114117 6621
rect 115375 6620 115378 6626
rect 115355 6606 115378 6620
rect 114088 6601 114117 6604
rect 115375 6600 115378 6606
rect 115404 6600 115407 6626
rect 116580 6620 116594 6640
rect 116856 6628 116916 6640
rect 116940 6638 116946 6655
rect 116963 6654 116969 6655
rect 116994 6654 117008 6674
rect 118596 6672 118602 6674
rect 118619 6672 118625 6689
rect 118596 6669 118625 6672
rect 118642 6689 118671 6692
rect 118642 6672 118648 6689
rect 118665 6688 118671 6689
rect 118963 6688 118966 6694
rect 118665 6674 118966 6688
rect 118665 6672 118671 6674
rect 118642 6669 118671 6672
rect 118963 6668 118966 6674
rect 118992 6668 118995 6694
rect 119055 6688 119058 6694
rect 119018 6674 119058 6688
rect 116963 6640 117008 6654
rect 117538 6655 117567 6658
rect 116963 6638 116969 6640
rect 116940 6635 116969 6638
rect 117538 6638 117544 6655
rect 117561 6654 117567 6655
rect 118550 6655 118579 6658
rect 118550 6654 118556 6655
rect 117561 6640 118556 6654
rect 117561 6638 117567 6640
rect 117538 6635 117567 6638
rect 118550 6638 118556 6640
rect 118573 6654 118579 6655
rect 119018 6654 119032 6674
rect 119055 6668 119058 6674
rect 119084 6668 119087 6694
rect 119156 6688 119170 6708
rect 119745 6702 119748 6728
rect 119774 6722 119777 6728
rect 119976 6723 120005 6726
rect 119976 6722 119982 6723
rect 119774 6708 119982 6722
rect 119774 6702 119777 6708
rect 119976 6706 119982 6708
rect 119999 6706 120005 6723
rect 119976 6703 120005 6706
rect 122321 6702 122324 6728
rect 122350 6722 122353 6728
rect 122689 6722 122692 6728
rect 122350 6708 122692 6722
rect 122350 6702 122353 6708
rect 122689 6702 122692 6708
rect 122718 6702 122721 6728
rect 123563 6722 123566 6728
rect 123543 6708 123566 6722
rect 123563 6702 123566 6708
rect 123592 6702 123595 6728
rect 124760 6723 124789 6726
rect 124760 6706 124766 6723
rect 124783 6722 124789 6723
rect 125541 6722 125544 6728
rect 124783 6708 125544 6722
rect 124783 6706 124789 6708
rect 124760 6703 124789 6706
rect 125541 6702 125544 6708
rect 125570 6702 125573 6728
rect 126231 6702 126234 6728
rect 126260 6722 126263 6728
rect 126416 6723 126445 6726
rect 126416 6722 126422 6723
rect 126260 6708 126422 6722
rect 126260 6702 126263 6708
rect 126416 6706 126422 6708
rect 126439 6706 126445 6723
rect 126416 6703 126445 6706
rect 127473 6702 127476 6728
rect 127502 6722 127505 6728
rect 127704 6723 127733 6726
rect 127704 6722 127710 6723
rect 127502 6708 127710 6722
rect 127502 6702 127505 6708
rect 127704 6706 127710 6708
rect 127727 6706 127733 6723
rect 129727 6722 129730 6728
rect 129707 6708 129730 6722
rect 127704 6703 127733 6706
rect 129727 6702 129730 6708
rect 129756 6702 129759 6728
rect 131338 6723 131367 6726
rect 131338 6706 131344 6723
rect 131361 6722 131367 6723
rect 131751 6722 131754 6728
rect 131361 6708 131754 6722
rect 131361 6706 131367 6708
rect 131338 6703 131367 6706
rect 131751 6702 131754 6708
rect 131780 6702 131783 6728
rect 132763 6702 132766 6728
rect 132792 6722 132795 6728
rect 132994 6723 133023 6726
rect 132994 6722 133000 6723
rect 132792 6708 133000 6722
rect 132792 6702 132795 6708
rect 132994 6706 133000 6708
rect 133017 6706 133023 6723
rect 132994 6703 133023 6706
rect 135201 6702 135204 6728
rect 135230 6722 135233 6728
rect 135230 6708 135914 6722
rect 135230 6702 135233 6708
rect 120390 6689 120419 6692
rect 120390 6688 120396 6689
rect 119156 6674 120396 6688
rect 120390 6672 120396 6674
rect 120413 6688 120419 6689
rect 121678 6689 121707 6692
rect 121678 6688 121684 6689
rect 120413 6674 121684 6688
rect 120413 6672 120419 6674
rect 120390 6669 120419 6672
rect 121678 6672 121684 6674
rect 121701 6672 121707 6689
rect 121678 6669 121707 6672
rect 122045 6668 122048 6694
rect 122074 6688 122077 6694
rect 122552 6689 122581 6692
rect 122552 6688 122558 6689
rect 122074 6674 122558 6688
rect 122074 6668 122077 6674
rect 122552 6672 122558 6674
rect 122575 6672 122581 6689
rect 122552 6669 122581 6672
rect 125082 6689 125111 6692
rect 125082 6672 125088 6689
rect 125105 6688 125111 6689
rect 125495 6688 125498 6694
rect 125105 6674 125498 6688
rect 125105 6672 125111 6674
rect 125082 6669 125111 6672
rect 119101 6654 119104 6660
rect 118573 6640 119032 6654
rect 119081 6640 119104 6654
rect 118573 6638 118579 6640
rect 118550 6635 118579 6638
rect 119101 6634 119104 6640
rect 119130 6634 119133 6660
rect 119883 6654 119886 6660
rect 119807 6640 119886 6654
rect 119883 6634 119886 6640
rect 119912 6634 119915 6660
rect 122560 6654 122574 6669
rect 125495 6668 125498 6674
rect 125524 6668 125527 6694
rect 131016 6689 131045 6692
rect 125550 6674 129888 6688
rect 125550 6660 125564 6674
rect 123656 6655 123685 6658
rect 123656 6654 123662 6655
rect 122560 6640 123662 6654
rect 123656 6638 123662 6640
rect 123679 6654 123685 6655
rect 124990 6655 125019 6658
rect 124990 6654 124996 6655
rect 123679 6640 124996 6654
rect 123679 6638 123685 6640
rect 123656 6635 123685 6638
rect 124990 6638 124996 6640
rect 125013 6638 125019 6655
rect 125541 6654 125544 6660
rect 125521 6640 125544 6654
rect 124990 6635 125019 6638
rect 125541 6634 125544 6640
rect 125570 6634 125573 6660
rect 126830 6655 126859 6658
rect 126830 6654 126836 6655
rect 126470 6640 126836 6654
rect 116028 6606 116594 6620
rect 116902 6620 116916 6628
rect 116902 6606 119216 6620
rect 112707 6586 112710 6592
rect 112092 6572 112114 6586
rect 112164 6572 112710 6586
rect 112092 6566 112095 6572
rect 112707 6566 112710 6572
rect 112736 6566 112739 6592
rect 112845 6586 112848 6592
rect 112825 6572 112848 6586
rect 112845 6566 112848 6572
rect 112874 6566 112877 6592
rect 113490 6587 113519 6590
rect 113490 6570 113496 6587
rect 113513 6586 113519 6587
rect 113535 6586 113538 6592
rect 113513 6572 113538 6586
rect 113513 6570 113519 6572
rect 113490 6567 113519 6570
rect 113535 6566 113538 6572
rect 113564 6586 113567 6592
rect 113811 6586 113814 6592
rect 113564 6572 113814 6586
rect 113564 6566 113567 6572
rect 113811 6566 113814 6572
rect 113840 6566 113843 6592
rect 113949 6586 113952 6592
rect 113905 6572 113952 6586
rect 113949 6566 113952 6572
rect 113978 6586 113981 6592
rect 116028 6586 116042 6606
rect 113978 6572 116042 6586
rect 113978 6566 113981 6572
rect 116065 6566 116068 6592
rect 116094 6586 116097 6592
rect 116572 6587 116601 6590
rect 116572 6586 116578 6587
rect 116094 6572 116578 6586
rect 116094 6566 116097 6572
rect 116572 6570 116578 6572
rect 116595 6570 116601 6587
rect 116572 6567 116601 6570
rect 116617 6566 116620 6592
rect 116646 6586 116649 6592
rect 116848 6587 116877 6590
rect 116848 6586 116854 6587
rect 116646 6572 116854 6586
rect 116646 6566 116649 6572
rect 116848 6570 116854 6572
rect 116871 6570 116877 6587
rect 117445 6586 117448 6592
rect 117425 6572 117448 6586
rect 116848 6567 116877 6570
rect 117445 6566 117448 6572
rect 117474 6566 117477 6592
rect 118366 6587 118395 6590
rect 118366 6570 118372 6587
rect 118389 6586 118395 6587
rect 118503 6586 118506 6592
rect 118389 6572 118506 6586
rect 118389 6570 118395 6572
rect 118366 6567 118395 6570
rect 118503 6566 118506 6572
rect 118532 6566 118535 6592
rect 119202 6586 119216 6606
rect 119239 6600 119242 6626
rect 119268 6620 119271 6626
rect 120527 6620 120530 6626
rect 119268 6606 119290 6620
rect 119892 6606 120044 6620
rect 120507 6606 120530 6620
rect 119268 6600 119271 6606
rect 119892 6586 119906 6606
rect 119202 6572 119906 6586
rect 120030 6586 120044 6606
rect 120527 6600 120530 6606
rect 120556 6600 120559 6626
rect 120895 6600 120898 6626
rect 120924 6600 120927 6626
rect 121815 6620 121818 6626
rect 121180 6606 121332 6620
rect 121795 6606 121818 6620
rect 121180 6586 121194 6606
rect 121263 6586 121266 6592
rect 120030 6572 121194 6586
rect 121243 6572 121266 6586
rect 121263 6566 121266 6572
rect 121292 6566 121295 6592
rect 121318 6586 121332 6606
rect 121815 6600 121818 6606
rect 121844 6600 121847 6626
rect 122459 6620 122462 6626
rect 122429 6606 122462 6620
rect 122459 6600 122462 6606
rect 122488 6600 122491 6626
rect 124860 6606 125656 6620
rect 124860 6586 124874 6606
rect 121318 6572 124874 6586
rect 124944 6587 124973 6590
rect 124944 6570 124950 6587
rect 124967 6586 124973 6587
rect 125587 6586 125590 6592
rect 124967 6572 125590 6586
rect 124967 6570 124973 6572
rect 124944 6567 124973 6570
rect 125587 6566 125590 6572
rect 125616 6566 125619 6592
rect 125642 6586 125656 6606
rect 125679 6600 125682 6626
rect 125708 6620 125711 6626
rect 125708 6606 125730 6620
rect 125708 6600 125711 6606
rect 126185 6600 126188 6626
rect 126214 6600 126217 6626
rect 126470 6586 126484 6640
rect 126830 6638 126836 6640
rect 126853 6638 126859 6655
rect 128117 6654 128120 6660
rect 126830 6635 126859 6638
rect 127620 6640 128120 6654
rect 126507 6600 126510 6626
rect 126536 6620 126539 6626
rect 126968 6621 126997 6624
rect 126968 6620 126974 6621
rect 126536 6606 126974 6620
rect 126536 6600 126539 6606
rect 126968 6604 126974 6606
rect 126991 6604 126997 6621
rect 126968 6601 126997 6604
rect 127473 6600 127476 6626
rect 127502 6600 127505 6626
rect 126737 6586 126740 6592
rect 125642 6572 126740 6586
rect 126737 6566 126740 6572
rect 126766 6586 126769 6592
rect 127620 6586 127634 6640
rect 128117 6634 128120 6640
rect 128146 6634 128149 6660
rect 129820 6655 129849 6658
rect 129820 6654 129826 6655
rect 128908 6640 129826 6654
rect 127657 6600 127660 6626
rect 127686 6620 127689 6626
rect 128256 6621 128285 6624
rect 128256 6620 128262 6621
rect 127686 6606 128262 6620
rect 127686 6600 127689 6606
rect 128256 6604 128262 6606
rect 128279 6604 128285 6621
rect 128256 6601 128285 6604
rect 128485 6600 128488 6626
rect 128514 6600 128517 6626
rect 126766 6572 127634 6586
rect 126766 6566 126769 6572
rect 128163 6566 128166 6592
rect 128192 6586 128195 6592
rect 128908 6586 128922 6640
rect 129820 6638 129826 6640
rect 129843 6638 129849 6655
rect 129874 6654 129888 6674
rect 131016 6672 131022 6689
rect 131039 6688 131045 6689
rect 131614 6689 131643 6692
rect 131614 6688 131620 6689
rect 131039 6674 131620 6688
rect 131039 6672 131045 6674
rect 131016 6669 131045 6672
rect 131614 6672 131620 6674
rect 131637 6688 131643 6689
rect 132073 6688 132076 6694
rect 131637 6674 132076 6688
rect 131637 6672 131643 6674
rect 131614 6669 131643 6672
rect 132073 6668 132076 6674
rect 132102 6668 132105 6694
rect 133270 6689 133299 6692
rect 133270 6688 133276 6689
rect 132128 6674 133276 6688
rect 132128 6658 132142 6674
rect 133270 6672 133276 6674
rect 133293 6688 133299 6689
rect 134558 6689 134587 6692
rect 134558 6688 134564 6689
rect 133293 6674 134564 6688
rect 133293 6672 133299 6674
rect 133270 6669 133299 6672
rect 134558 6672 134564 6674
rect 134581 6688 134587 6689
rect 135846 6689 135875 6692
rect 135846 6688 135852 6689
rect 134581 6674 135852 6688
rect 134581 6672 134587 6674
rect 134558 6669 134587 6672
rect 135846 6672 135852 6674
rect 135869 6672 135875 6689
rect 135900 6688 135914 6708
rect 136489 6702 136492 6728
rect 136518 6722 136521 6728
rect 136518 6708 139042 6722
rect 136518 6702 136521 6708
rect 135900 6674 136558 6688
rect 135846 6669 135875 6672
rect 132120 6655 132149 6658
rect 132120 6654 132126 6655
rect 129874 6640 132126 6654
rect 129820 6635 129849 6638
rect 132120 6638 132126 6640
rect 132143 6638 132149 6655
rect 132120 6635 132149 6638
rect 134282 6655 134311 6658
rect 134282 6638 134288 6655
rect 134305 6654 134311 6655
rect 134465 6654 134468 6660
rect 134305 6640 134468 6654
rect 134305 6638 134311 6640
rect 134282 6635 134311 6638
rect 134465 6634 134468 6640
rect 134494 6634 134497 6660
rect 136544 6647 136558 6674
rect 136581 6668 136584 6694
rect 136610 6688 136613 6694
rect 136610 6674 138996 6688
rect 136610 6668 136613 6674
rect 136627 6634 136630 6660
rect 136656 6654 136659 6660
rect 137226 6655 137255 6658
rect 137226 6654 137232 6655
rect 136656 6640 137232 6654
rect 136656 6634 136659 6640
rect 137226 6638 137232 6640
rect 137249 6638 137255 6655
rect 137547 6654 137550 6660
rect 137527 6640 137550 6654
rect 137226 6635 137255 6638
rect 137547 6634 137550 6640
rect 137576 6634 137579 6660
rect 130923 6620 130926 6626
rect 130903 6606 130926 6620
rect 130923 6600 130926 6606
rect 130952 6600 130955 6626
rect 131522 6621 131551 6624
rect 131522 6604 131528 6621
rect 131545 6620 131551 6621
rect 131705 6620 131708 6626
rect 131545 6606 131708 6620
rect 131545 6604 131551 6606
rect 131522 6601 131551 6604
rect 131705 6600 131708 6606
rect 131734 6600 131737 6626
rect 131751 6600 131754 6626
rect 131780 6620 131783 6626
rect 132211 6620 132214 6626
rect 131780 6606 132214 6620
rect 131780 6600 131783 6606
rect 132211 6600 132214 6606
rect 132240 6600 132243 6626
rect 132258 6621 132287 6624
rect 132258 6604 132264 6621
rect 132281 6620 132287 6621
rect 132303 6620 132306 6626
rect 132281 6606 132306 6620
rect 132281 6604 132287 6606
rect 132258 6601 132287 6604
rect 132303 6600 132306 6606
rect 132332 6600 132335 6626
rect 132487 6600 132490 6626
rect 132516 6600 132519 6626
rect 133408 6621 133437 6624
rect 132956 6606 133384 6620
rect 128192 6572 128922 6586
rect 128192 6566 128195 6572
rect 128991 6566 128994 6592
rect 129020 6586 129023 6592
rect 131475 6586 131478 6592
rect 129020 6572 131478 6586
rect 129020 6566 129023 6572
rect 131475 6566 131478 6572
rect 131504 6586 131507 6592
rect 131568 6587 131597 6590
rect 131568 6586 131574 6587
rect 131504 6572 131574 6586
rect 131504 6566 131507 6572
rect 131568 6570 131574 6572
rect 131591 6570 131597 6587
rect 131568 6567 131597 6570
rect 131659 6566 131662 6592
rect 131688 6586 131691 6592
rect 132956 6586 132970 6606
rect 131688 6572 132970 6586
rect 133370 6586 133384 6606
rect 133408 6604 133414 6621
rect 133431 6620 133437 6621
rect 133453 6620 133456 6626
rect 133431 6606 133456 6620
rect 133431 6604 133437 6606
rect 133408 6601 133437 6604
rect 133453 6600 133456 6606
rect 133482 6600 133485 6626
rect 134021 6606 134258 6620
rect 133821 6586 133824 6592
rect 133370 6572 133824 6586
rect 131688 6566 131691 6572
rect 133821 6566 133824 6572
rect 133850 6566 133853 6592
rect 134244 6586 134258 6606
rect 134373 6600 134376 6626
rect 134402 6620 134405 6626
rect 134402 6606 134941 6620
rect 134402 6600 134405 6606
rect 135339 6600 135342 6626
rect 135368 6620 135371 6626
rect 135368 6606 135454 6620
rect 135368 6600 135371 6606
rect 135385 6586 135388 6592
rect 134244 6572 135388 6586
rect 135385 6566 135388 6572
rect 135414 6566 135417 6592
rect 135440 6590 135454 6606
rect 135477 6600 135480 6626
rect 135506 6620 135509 6626
rect 135984 6621 136013 6624
rect 135984 6620 135990 6621
rect 135506 6606 135990 6620
rect 135506 6600 135509 6606
rect 135984 6604 135990 6606
rect 136007 6604 136013 6621
rect 138982 6620 138996 6674
rect 139028 6658 139042 6708
rect 151678 6688 151692 6737
rect 152222 6689 152251 6692
rect 152222 6688 152228 6689
rect 139074 6674 146724 6688
rect 151678 6674 152228 6688
rect 139020 6655 139049 6658
rect 139020 6638 139026 6655
rect 139043 6638 139049 6655
rect 139020 6635 139049 6638
rect 139074 6620 139088 6674
rect 140537 6654 140540 6660
rect 140517 6640 140540 6654
rect 140537 6634 140540 6640
rect 140566 6634 140569 6660
rect 142377 6654 142380 6660
rect 142357 6640 142380 6654
rect 142377 6634 142380 6640
rect 142406 6634 142409 6660
rect 143666 6655 143695 6658
rect 143666 6654 143672 6655
rect 143513 6640 143672 6654
rect 143513 6620 143527 6640
rect 143666 6638 143672 6640
rect 143689 6638 143695 6655
rect 145137 6654 145140 6660
rect 145117 6640 145140 6654
rect 143666 6635 143695 6638
rect 145137 6634 145140 6640
rect 145166 6634 145169 6660
rect 146710 6658 146724 6674
rect 152222 6672 152228 6674
rect 152245 6688 152251 6689
rect 152452 6689 152481 6692
rect 152452 6688 152458 6689
rect 152245 6674 152458 6688
rect 152245 6672 152251 6674
rect 152222 6669 152251 6672
rect 152452 6672 152458 6674
rect 152475 6688 152481 6689
rect 152497 6688 152500 6694
rect 152475 6674 152500 6688
rect 152475 6672 152481 6674
rect 152452 6669 152481 6672
rect 152497 6668 152500 6674
rect 152526 6688 152529 6694
rect 152682 6689 152711 6692
rect 152682 6688 152688 6689
rect 152526 6674 152688 6688
rect 152526 6668 152529 6674
rect 152682 6672 152688 6674
rect 152705 6672 152711 6689
rect 152682 6669 152711 6672
rect 146702 6655 146731 6658
rect 146702 6638 146708 6655
rect 146725 6638 146731 6655
rect 148220 6655 148249 6658
rect 148220 6654 148226 6655
rect 146702 6635 146731 6638
rect 147952 6640 148226 6654
rect 138982 6606 139088 6620
rect 141443 6606 143527 6620
rect 135984 6601 136013 6604
rect 135432 6587 135461 6590
rect 135432 6570 135438 6587
rect 135455 6586 135461 6587
rect 135891 6586 135894 6592
rect 135455 6572 135894 6586
rect 135455 6570 135461 6572
rect 135432 6567 135461 6570
rect 135891 6566 135894 6572
rect 135920 6566 135923 6592
rect 136443 6566 136446 6592
rect 136472 6586 136475 6592
rect 136720 6587 136749 6590
rect 136720 6586 136726 6587
rect 136472 6572 136726 6586
rect 136472 6566 136475 6572
rect 136720 6570 136726 6572
rect 136743 6586 136749 6587
rect 141443 6586 141457 6606
rect 147952 6592 147966 6640
rect 148220 6638 148226 6640
rect 148243 6638 148249 6655
rect 149737 6654 149740 6660
rect 149717 6640 149740 6654
rect 148220 6635 148249 6638
rect 149737 6634 149740 6640
rect 149766 6634 149769 6660
rect 151761 6634 151764 6660
rect 151790 6654 151793 6660
rect 151854 6655 151883 6658
rect 151854 6654 151860 6655
rect 151790 6640 151860 6654
rect 151790 6634 151793 6640
rect 151854 6638 151860 6640
rect 151877 6638 151883 6655
rect 151854 6635 151883 6638
rect 147943 6586 147946 6592
rect 136743 6572 141457 6586
rect 147923 6572 147946 6586
rect 136743 6570 136749 6572
rect 136720 6567 136749 6570
rect 147943 6566 147946 6572
rect 147972 6566 147975 6592
rect 552 6541 152904 6552
rect 552 6515 38574 6541
rect 38600 6515 38606 6541
rect 38632 6515 38638 6541
rect 38664 6515 38670 6541
rect 38696 6515 38702 6541
rect 38728 6515 76673 6541
rect 76699 6515 76705 6541
rect 76731 6515 76737 6541
rect 76763 6515 76769 6541
rect 76795 6515 76801 6541
rect 76827 6515 114772 6541
rect 114798 6515 114804 6541
rect 114830 6515 114836 6541
rect 114862 6515 114868 6541
rect 114894 6515 114900 6541
rect 114926 6515 152904 6541
rect 552 6504 152904 6515
rect 13025 6484 13028 6490
rect 13005 6470 13028 6484
rect 13025 6464 13028 6470
rect 13054 6464 13057 6490
rect 13716 6485 13745 6488
rect 13716 6468 13722 6485
rect 13739 6468 13745 6485
rect 16107 6484 16110 6490
rect 13716 6465 13745 6468
rect 13816 6470 16110 6484
rect 10081 6430 10084 6456
rect 10110 6450 10113 6456
rect 10110 6436 11047 6450
rect 10110 6430 10113 6436
rect 11033 6314 11047 6436
rect 13669 6430 13672 6456
rect 13698 6450 13701 6456
rect 13724 6450 13738 6465
rect 13698 6436 13738 6450
rect 13698 6430 13701 6436
rect 13118 6417 13147 6420
rect 13118 6400 13124 6417
rect 13141 6416 13147 6417
rect 13816 6416 13830 6470
rect 16107 6464 16110 6470
rect 16136 6484 16139 6490
rect 16936 6485 16965 6488
rect 16936 6484 16942 6485
rect 16136 6470 16942 6484
rect 16136 6464 16139 6470
rect 16936 6468 16942 6470
rect 16959 6468 16965 6485
rect 16936 6465 16965 6468
rect 17073 6464 17076 6490
rect 17102 6484 17105 6490
rect 17396 6485 17425 6488
rect 17396 6484 17402 6485
rect 17102 6470 17402 6484
rect 17102 6464 17105 6470
rect 17396 6468 17402 6470
rect 17419 6468 17425 6485
rect 17763 6484 17766 6490
rect 17743 6470 17766 6484
rect 17396 6465 17425 6468
rect 17763 6464 17766 6470
rect 17792 6464 17795 6490
rect 18316 6485 18345 6488
rect 18316 6484 18322 6485
rect 17818 6470 18322 6484
rect 14497 6450 14500 6456
rect 13141 6402 13830 6416
rect 13862 6436 14500 6450
rect 13141 6400 13147 6402
rect 13118 6397 13147 6400
rect 11599 6362 11602 6388
rect 11628 6382 11631 6388
rect 13862 6382 13876 6436
rect 14497 6430 14500 6436
rect 14526 6430 14529 6456
rect 15187 6450 15190 6456
rect 14552 6436 15190 6450
rect 13900 6417 13929 6420
rect 13900 6400 13906 6417
rect 13923 6416 13929 6417
rect 13991 6416 13994 6422
rect 13923 6402 13994 6416
rect 13923 6400 13929 6402
rect 13900 6397 13929 6400
rect 13991 6396 13994 6402
rect 14020 6396 14023 6422
rect 11628 6368 13876 6382
rect 13946 6383 13975 6386
rect 11628 6362 11631 6368
rect 13946 6366 13952 6383
rect 13969 6366 13975 6383
rect 14037 6382 14040 6388
rect 14017 6368 14040 6382
rect 13946 6363 13975 6366
rect 13577 6328 13580 6354
rect 13606 6348 13609 6354
rect 13954 6348 13968 6363
rect 14037 6362 14040 6368
rect 14066 6362 14069 6388
rect 14552 6386 14566 6436
rect 15187 6430 15190 6436
rect 15216 6430 15219 6456
rect 15785 6450 15788 6456
rect 15663 6436 15788 6450
rect 15785 6430 15788 6436
rect 15814 6430 15817 6456
rect 17211 6450 17214 6456
rect 16813 6436 17214 6450
rect 17211 6430 17214 6436
rect 17240 6430 17243 6456
rect 17818 6450 17832 6470
rect 18316 6468 18322 6470
rect 18339 6468 18345 6485
rect 21260 6485 21289 6488
rect 18316 6465 18345 6468
rect 18692 6470 20707 6484
rect 18692 6454 18706 6470
rect 17266 6436 17832 6450
rect 18270 6451 18299 6454
rect 16843 6396 16846 6422
rect 16872 6416 16875 6422
rect 17266 6416 17280 6436
rect 18270 6434 18276 6451
rect 18293 6450 18299 6451
rect 18684 6451 18713 6454
rect 18684 6450 18690 6451
rect 18293 6436 18690 6450
rect 18293 6434 18299 6436
rect 18270 6431 18299 6434
rect 18684 6434 18690 6436
rect 18707 6434 18713 6451
rect 18684 6431 18713 6434
rect 18729 6430 18732 6456
rect 18758 6450 18761 6456
rect 19236 6451 19265 6454
rect 19236 6450 19242 6451
rect 18758 6436 19242 6450
rect 18758 6430 18761 6436
rect 19236 6434 19242 6436
rect 19259 6434 19265 6451
rect 19236 6431 19265 6434
rect 19833 6430 19836 6456
rect 19862 6450 19865 6456
rect 19880 6451 19909 6454
rect 19880 6450 19886 6451
rect 19862 6436 19886 6450
rect 19862 6430 19865 6436
rect 19880 6434 19886 6436
rect 19903 6434 19909 6451
rect 20523 6450 20526 6456
rect 20493 6436 20526 6450
rect 19880 6431 19909 6434
rect 20523 6430 20526 6436
rect 20552 6430 20555 6456
rect 20693 6450 20707 6470
rect 21260 6468 21266 6485
rect 21283 6484 21289 6485
rect 21627 6484 21630 6490
rect 21283 6470 21630 6484
rect 21283 6468 21289 6470
rect 21260 6465 21289 6468
rect 21627 6464 21630 6470
rect 21656 6464 21659 6490
rect 21720 6485 21749 6488
rect 21720 6468 21726 6485
rect 21743 6484 21749 6485
rect 22133 6484 22136 6490
rect 21743 6470 22136 6484
rect 21743 6468 21749 6470
rect 21720 6465 21749 6468
rect 22133 6464 22136 6470
rect 22162 6464 22165 6490
rect 22271 6484 22274 6490
rect 22251 6470 22274 6484
rect 22271 6464 22274 6470
rect 22300 6464 22303 6490
rect 25998 6485 26027 6488
rect 25998 6468 26004 6485
rect 26021 6484 26027 6485
rect 26641 6484 26644 6490
rect 26021 6470 26644 6484
rect 26021 6468 26027 6470
rect 25998 6465 26027 6468
rect 26641 6464 26644 6470
rect 26670 6464 26673 6490
rect 26780 6485 26809 6488
rect 26780 6468 26786 6485
rect 26803 6468 26809 6485
rect 26780 6465 26809 6468
rect 26964 6485 26993 6488
rect 26964 6468 26970 6485
rect 26987 6484 26993 6485
rect 27331 6484 27334 6490
rect 26987 6470 27334 6484
rect 26987 6468 26993 6470
rect 26964 6465 26993 6468
rect 21489 6450 21492 6456
rect 20693 6436 21492 6450
rect 21489 6430 21492 6436
rect 21518 6430 21521 6456
rect 26788 6450 26802 6465
rect 27331 6464 27334 6470
rect 27360 6464 27363 6490
rect 27929 6464 27932 6490
rect 27958 6484 27961 6490
rect 28987 6484 28990 6490
rect 27958 6470 28990 6484
rect 27958 6464 27961 6470
rect 28987 6464 28990 6470
rect 29016 6464 29019 6490
rect 29264 6485 29293 6488
rect 29264 6468 29270 6485
rect 29287 6484 29293 6485
rect 29815 6484 29818 6490
rect 29287 6470 29818 6484
rect 29287 6468 29293 6470
rect 29264 6465 29293 6468
rect 29815 6464 29818 6470
rect 29844 6464 29847 6490
rect 36071 6484 36074 6490
rect 36051 6470 36074 6484
rect 36071 6464 36074 6470
rect 36100 6464 36103 6490
rect 36163 6464 36166 6490
rect 36192 6484 36195 6490
rect 37359 6484 37362 6490
rect 36192 6470 37362 6484
rect 36192 6464 36195 6470
rect 37359 6464 37362 6470
rect 37388 6464 37391 6490
rect 41959 6484 41962 6490
rect 37782 6470 41962 6484
rect 26098 6436 26802 6450
rect 16872 6402 17280 6416
rect 17350 6417 17379 6420
rect 16872 6396 16875 6402
rect 17350 6400 17356 6417
rect 17373 6400 17379 6417
rect 17350 6397 17379 6400
rect 17856 6417 17885 6420
rect 17856 6400 17862 6417
rect 17879 6416 17885 6417
rect 19190 6417 19219 6420
rect 19190 6416 19196 6417
rect 17879 6402 19196 6416
rect 17879 6400 17885 6402
rect 17856 6397 17885 6400
rect 19190 6400 19196 6402
rect 19213 6416 19219 6417
rect 19649 6416 19652 6422
rect 19213 6402 19652 6416
rect 19213 6400 19219 6402
rect 19190 6397 19219 6400
rect 14544 6383 14573 6386
rect 14544 6382 14550 6383
rect 14138 6368 14550 6382
rect 13606 6334 13968 6348
rect 13606 6328 13609 6334
rect 14138 6314 14152 6368
rect 14544 6366 14550 6368
rect 14567 6366 14573 6383
rect 14544 6363 14573 6366
rect 14636 6383 14665 6386
rect 14636 6366 14642 6383
rect 14659 6382 14665 6383
rect 14819 6382 14822 6388
rect 14659 6368 14822 6382
rect 14659 6366 14665 6368
rect 14636 6363 14665 6366
rect 14819 6362 14822 6368
rect 14848 6362 14851 6388
rect 14911 6382 14914 6388
rect 14867 6368 14914 6382
rect 14911 6362 14914 6368
rect 14940 6362 14943 6388
rect 15049 6382 15052 6388
rect 15029 6368 15052 6382
rect 15049 6362 15052 6368
rect 15078 6362 15081 6388
rect 16062 6383 16091 6386
rect 16062 6366 16068 6383
rect 16085 6366 16091 6383
rect 16062 6363 16091 6366
rect 16200 6383 16229 6386
rect 16200 6366 16206 6383
rect 16223 6382 16229 6383
rect 16521 6382 16524 6388
rect 16223 6368 16524 6382
rect 16223 6366 16229 6368
rect 16200 6363 16229 6366
rect 11033 6300 14152 6314
rect 14314 6315 14343 6318
rect 14314 6298 14320 6315
rect 14337 6314 14343 6315
rect 14451 6314 14454 6320
rect 14337 6300 14454 6314
rect 14337 6298 14343 6300
rect 14314 6295 14343 6298
rect 14451 6294 14454 6300
rect 14480 6294 14483 6320
rect 14920 6314 14934 6362
rect 16070 6348 16084 6363
rect 16521 6362 16524 6368
rect 16550 6362 16553 6388
rect 16705 6362 16708 6388
rect 16734 6382 16737 6388
rect 17165 6382 17168 6388
rect 16734 6368 17168 6382
rect 16734 6362 16737 6368
rect 17165 6362 17168 6368
rect 17194 6382 17197 6388
rect 17358 6382 17372 6397
rect 19649 6396 19652 6402
rect 19678 6396 19681 6422
rect 20753 6396 20756 6422
rect 20782 6416 20785 6422
rect 20846 6417 20875 6420
rect 20846 6416 20852 6417
rect 20782 6402 20852 6416
rect 20782 6396 20785 6402
rect 20846 6400 20852 6402
rect 20869 6416 20875 6417
rect 21214 6417 21243 6420
rect 21214 6416 21220 6417
rect 20869 6402 21220 6416
rect 20869 6400 20875 6402
rect 20846 6397 20875 6400
rect 21214 6400 21220 6402
rect 21237 6400 21243 6417
rect 22364 6417 22393 6420
rect 22364 6416 22370 6417
rect 21214 6397 21243 6400
rect 21774 6402 22370 6416
rect 17194 6368 17372 6382
rect 17194 6362 17197 6368
rect 17441 6362 17444 6388
rect 17470 6382 17473 6388
rect 17470 6368 17492 6382
rect 17470 6362 17473 6368
rect 17671 6362 17674 6388
rect 17700 6382 17703 6388
rect 18776 6383 18805 6386
rect 18776 6382 18782 6383
rect 17700 6368 18782 6382
rect 17700 6362 17703 6368
rect 18776 6366 18782 6368
rect 18799 6366 18805 6383
rect 18776 6363 18805 6366
rect 19282 6383 19311 6386
rect 19282 6366 19288 6383
rect 19305 6382 19311 6383
rect 19695 6382 19698 6388
rect 19305 6368 19698 6382
rect 19305 6366 19311 6368
rect 19282 6363 19311 6366
rect 19695 6362 19698 6368
rect 19724 6362 19727 6388
rect 19742 6383 19771 6386
rect 19742 6366 19748 6383
rect 19765 6366 19771 6383
rect 19742 6363 19771 6366
rect 19750 6348 19764 6363
rect 20477 6362 20480 6388
rect 20506 6382 20509 6388
rect 21535 6382 21538 6388
rect 20506 6368 21538 6382
rect 20506 6362 20509 6368
rect 21535 6362 21538 6368
rect 21564 6362 21567 6388
rect 21581 6362 21584 6388
rect 21610 6382 21613 6388
rect 21774 6386 21788 6402
rect 22364 6400 22370 6402
rect 22387 6416 22393 6417
rect 22685 6416 22688 6422
rect 22387 6402 22688 6416
rect 22387 6400 22393 6402
rect 22364 6397 22393 6400
rect 22685 6396 22688 6402
rect 22714 6396 22717 6422
rect 26098 6420 26112 6436
rect 27745 6430 27748 6456
rect 27774 6430 27777 6456
rect 28665 6430 28668 6456
rect 28694 6450 28697 6456
rect 29310 6451 29339 6454
rect 29310 6450 29316 6451
rect 28694 6436 29316 6450
rect 28694 6430 28697 6436
rect 29310 6434 29316 6436
rect 29333 6450 29339 6451
rect 30321 6450 30324 6456
rect 29333 6436 30324 6450
rect 29333 6434 29339 6436
rect 29310 6431 29339 6434
rect 30321 6430 30324 6436
rect 30350 6430 30353 6456
rect 32943 6430 32946 6456
rect 32972 6450 32975 6456
rect 37782 6450 37796 6470
rect 38924 6451 38953 6454
rect 38924 6450 38930 6451
rect 32972 6436 37796 6450
rect 38525 6436 38930 6450
rect 32972 6430 32975 6436
rect 26090 6417 26119 6420
rect 26090 6400 26096 6417
rect 26113 6400 26119 6417
rect 26090 6397 26119 6400
rect 26458 6417 26487 6420
rect 26458 6400 26464 6417
rect 26481 6416 26487 6417
rect 26871 6416 26874 6422
rect 26481 6402 26874 6416
rect 26481 6400 26487 6402
rect 26458 6397 26487 6400
rect 26871 6396 26874 6402
rect 26900 6396 26903 6422
rect 27009 6419 27012 6422
rect 26972 6416 27012 6419
rect 26926 6402 27012 6416
rect 21766 6383 21795 6386
rect 21766 6382 21772 6383
rect 21610 6368 21772 6382
rect 21610 6362 21613 6368
rect 21766 6366 21772 6368
rect 21789 6366 21795 6383
rect 21766 6363 21795 6366
rect 21858 6383 21887 6386
rect 21858 6366 21864 6383
rect 21881 6382 21887 6383
rect 21903 6382 21906 6388
rect 21881 6368 21906 6382
rect 21881 6366 21887 6368
rect 21858 6363 21887 6366
rect 21903 6362 21906 6368
rect 21932 6382 21935 6388
rect 22731 6382 22734 6388
rect 21932 6368 22734 6382
rect 21932 6362 21935 6368
rect 22731 6362 22734 6368
rect 22760 6362 22763 6388
rect 25675 6362 25678 6388
rect 25704 6382 25707 6388
rect 26926 6382 26940 6402
rect 27009 6396 27012 6402
rect 27038 6396 27041 6422
rect 27377 6418 27380 6422
rect 27340 6416 27380 6418
rect 27333 6402 27380 6416
rect 27055 6382 27058 6388
rect 25704 6368 26940 6382
rect 27035 6368 27058 6382
rect 25704 6362 25707 6368
rect 27055 6362 27058 6368
rect 27084 6362 27087 6388
rect 27340 6348 27354 6402
rect 27377 6396 27380 6402
rect 27406 6396 27409 6422
rect 28528 6417 28557 6420
rect 28528 6400 28534 6417
rect 28551 6416 28557 6417
rect 28711 6416 28714 6422
rect 28551 6402 28714 6416
rect 28551 6400 28557 6402
rect 28528 6397 28557 6400
rect 28711 6396 28714 6402
rect 28740 6396 28743 6422
rect 36164 6417 36193 6420
rect 36164 6400 36170 6417
rect 36187 6416 36193 6417
rect 37405 6416 37408 6422
rect 36187 6402 37408 6416
rect 36187 6400 36193 6402
rect 36164 6397 36193 6400
rect 37405 6396 37408 6402
rect 37434 6396 37437 6422
rect 37544 6417 37573 6420
rect 37544 6400 37550 6417
rect 37567 6416 37573 6417
rect 37727 6416 37730 6422
rect 37567 6402 37730 6416
rect 37567 6400 37573 6402
rect 37544 6397 37573 6400
rect 37727 6396 37730 6402
rect 37756 6396 37759 6422
rect 37782 6420 37796 6436
rect 38924 6434 38930 6436
rect 38947 6434 38953 6451
rect 38924 6431 38953 6434
rect 39199 6430 39202 6456
rect 39228 6450 39231 6456
rect 39292 6451 39321 6454
rect 39292 6450 39298 6451
rect 39228 6436 39298 6450
rect 39228 6430 39231 6436
rect 39292 6434 39298 6436
rect 39315 6434 39321 6451
rect 39292 6431 39321 6434
rect 37774 6417 37803 6420
rect 37774 6400 37780 6417
rect 37797 6400 37803 6417
rect 37774 6397 37803 6400
rect 38878 6417 38907 6420
rect 38878 6400 38884 6417
rect 38901 6416 38907 6417
rect 39246 6417 39275 6420
rect 39246 6416 39252 6417
rect 38901 6402 39252 6416
rect 38901 6400 38907 6402
rect 38878 6397 38907 6400
rect 39246 6400 39252 6402
rect 39269 6416 39275 6417
rect 39660 6417 39689 6420
rect 39269 6402 39314 6416
rect 39269 6400 39275 6402
rect 39246 6397 39275 6400
rect 39300 6388 39314 6402
rect 39660 6400 39666 6417
rect 39683 6416 39689 6417
rect 39843 6416 39846 6422
rect 39683 6402 39846 6416
rect 39683 6400 39689 6402
rect 39660 6397 39689 6400
rect 39843 6396 39846 6402
rect 39872 6396 39875 6422
rect 39898 6420 39912 6470
rect 41959 6464 41962 6470
rect 41988 6464 41991 6490
rect 43247 6484 43250 6490
rect 42336 6470 43250 6484
rect 40257 6430 40260 6456
rect 40286 6430 40289 6456
rect 41453 6430 41456 6456
rect 41482 6450 41485 6456
rect 42336 6450 42350 6470
rect 43247 6464 43250 6470
rect 43276 6464 43279 6490
rect 43569 6484 43572 6490
rect 43440 6470 43572 6484
rect 43440 6450 43454 6470
rect 43569 6464 43572 6470
rect 43598 6464 43601 6490
rect 44766 6485 44795 6488
rect 44766 6468 44772 6485
rect 44789 6484 44795 6485
rect 44789 6470 44857 6484
rect 44789 6468 44795 6470
rect 44766 6465 44795 6468
rect 44843 6450 44857 6470
rect 45225 6464 45228 6490
rect 45254 6484 45257 6490
rect 45548 6485 45577 6488
rect 45548 6484 45554 6485
rect 45254 6470 45554 6484
rect 45254 6464 45257 6470
rect 45548 6468 45554 6470
rect 45571 6468 45577 6485
rect 45548 6465 45577 6468
rect 45823 6464 45826 6490
rect 45852 6484 45855 6490
rect 48997 6484 49000 6490
rect 45852 6470 49000 6484
rect 45852 6464 45855 6470
rect 48997 6464 49000 6470
rect 49026 6464 49029 6490
rect 49673 6470 54172 6484
rect 45271 6450 45274 6456
rect 41482 6436 42350 6450
rect 42757 6436 43454 6450
rect 43861 6436 44788 6450
rect 44843 6436 45274 6450
rect 41482 6430 41485 6436
rect 39890 6417 39919 6420
rect 39890 6400 39896 6417
rect 39913 6400 39919 6417
rect 43110 6417 43139 6420
rect 43110 6416 43116 6417
rect 39890 6397 39919 6400
rect 42750 6402 43116 6416
rect 27515 6382 27518 6388
rect 27495 6368 27518 6382
rect 27515 6362 27518 6368
rect 27544 6362 27547 6388
rect 29356 6383 29385 6386
rect 29356 6366 29362 6383
rect 29379 6366 29385 6383
rect 37912 6383 37941 6386
rect 37912 6382 37918 6383
rect 29356 6363 29385 6366
rect 37460 6368 37918 6382
rect 29364 6348 29378 6363
rect 37460 6352 37474 6368
rect 37912 6366 37918 6368
rect 37935 6366 37941 6383
rect 37912 6363 37941 6366
rect 39291 6362 39294 6388
rect 39320 6362 39323 6388
rect 40028 6383 40057 6386
rect 40028 6382 40034 6383
rect 39576 6368 40034 6382
rect 15564 6334 16084 6348
rect 15564 6314 15578 6334
rect 14920 6300 15578 6314
rect 15693 6294 15696 6320
rect 15722 6314 15725 6320
rect 15786 6315 15815 6318
rect 15786 6314 15792 6315
rect 15722 6300 15792 6314
rect 15722 6294 15725 6300
rect 15786 6298 15792 6300
rect 15809 6298 15815 6315
rect 16070 6314 16084 6334
rect 16714 6334 19764 6348
rect 16199 6314 16202 6320
rect 16070 6300 16202 6314
rect 15786 6295 15815 6298
rect 16199 6294 16202 6300
rect 16228 6314 16231 6320
rect 16714 6314 16728 6334
rect 16228 6300 16728 6314
rect 16228 6294 16231 6300
rect 17073 6294 17076 6320
rect 17102 6314 17105 6320
rect 17166 6315 17195 6318
rect 17166 6314 17172 6315
rect 17102 6300 17172 6314
rect 17102 6294 17105 6300
rect 17166 6298 17172 6300
rect 17189 6298 17195 6315
rect 19005 6314 19008 6320
rect 18985 6300 19008 6314
rect 17166 6295 17195 6298
rect 19005 6294 19008 6300
rect 19034 6294 19037 6320
rect 19750 6314 19764 6334
rect 20394 6334 27354 6348
rect 28168 6334 29378 6348
rect 37452 6349 37481 6352
rect 20394 6314 20408 6334
rect 28168 6320 28182 6334
rect 20615 6314 20618 6320
rect 19750 6300 20408 6314
rect 20595 6300 20618 6314
rect 20615 6294 20618 6300
rect 20644 6294 20647 6320
rect 20891 6314 20894 6320
rect 20871 6300 20894 6314
rect 20891 6294 20894 6300
rect 20920 6294 20923 6320
rect 21397 6294 21400 6320
rect 21426 6314 21429 6320
rect 21536 6315 21565 6318
rect 21536 6314 21542 6315
rect 21426 6300 21542 6314
rect 21426 6294 21429 6300
rect 21536 6298 21542 6300
rect 21559 6298 21565 6315
rect 21536 6295 21565 6298
rect 21627 6294 21630 6320
rect 21656 6314 21659 6320
rect 21903 6314 21906 6320
rect 21656 6300 21906 6314
rect 21656 6294 21659 6300
rect 21903 6294 21906 6300
rect 21932 6294 21935 6320
rect 26504 6315 26533 6318
rect 26504 6298 26510 6315
rect 26527 6314 26533 6315
rect 26549 6314 26552 6320
rect 26527 6300 26552 6314
rect 26527 6298 26533 6300
rect 26504 6295 26533 6298
rect 26549 6294 26552 6300
rect 26578 6294 26581 6320
rect 27055 6294 27058 6320
rect 27084 6314 27087 6320
rect 27791 6314 27794 6320
rect 27084 6300 27794 6314
rect 27084 6294 27087 6300
rect 27791 6294 27794 6300
rect 27820 6314 27823 6320
rect 28159 6314 28162 6320
rect 27820 6300 28162 6314
rect 27820 6294 27823 6300
rect 28159 6294 28162 6300
rect 28188 6294 28191 6320
rect 28251 6314 28254 6320
rect 28231 6300 28254 6314
rect 28251 6294 28254 6300
rect 28280 6294 28283 6320
rect 28582 6318 28596 6334
rect 37452 6332 37458 6349
rect 37475 6332 37481 6349
rect 38923 6348 38926 6354
rect 37452 6329 37481 6332
rect 38426 6334 38926 6348
rect 28574 6315 28603 6318
rect 28574 6298 28580 6315
rect 28597 6298 28603 6315
rect 28574 6295 28603 6298
rect 28619 6294 28622 6320
rect 28648 6314 28651 6320
rect 29080 6315 29109 6318
rect 29080 6314 29086 6315
rect 28648 6300 29086 6314
rect 28648 6294 28651 6300
rect 29080 6298 29086 6300
rect 29103 6298 29109 6315
rect 29080 6295 29109 6298
rect 36347 6294 36350 6320
rect 36376 6314 36379 6320
rect 37497 6314 37500 6320
rect 36376 6300 37500 6314
rect 36376 6294 36379 6300
rect 37497 6294 37500 6300
rect 37526 6294 37529 6320
rect 37589 6294 37592 6320
rect 37618 6314 37621 6320
rect 38426 6314 38440 6334
rect 38923 6328 38926 6334
rect 38952 6328 38955 6354
rect 39061 6328 39064 6354
rect 39090 6348 39093 6354
rect 39576 6352 39590 6368
rect 40028 6366 40034 6368
rect 40051 6366 40057 6383
rect 40028 6363 40057 6366
rect 40395 6362 40398 6388
rect 40424 6382 40427 6388
rect 42006 6383 42035 6386
rect 42006 6382 42012 6383
rect 40424 6368 42012 6382
rect 40424 6362 40427 6368
rect 42006 6366 42012 6368
rect 42029 6366 42035 6383
rect 42006 6363 42035 6366
rect 42144 6383 42173 6386
rect 42144 6366 42150 6383
rect 42167 6382 42173 6383
rect 42419 6382 42422 6388
rect 42167 6368 42422 6382
rect 42167 6366 42173 6368
rect 42144 6363 42173 6366
rect 39568 6349 39597 6352
rect 39090 6334 39360 6348
rect 39090 6328 39093 6334
rect 37618 6300 38440 6314
rect 37618 6294 37621 6300
rect 38601 6294 38604 6320
rect 38630 6314 38633 6320
rect 38648 6315 38677 6318
rect 38648 6314 38654 6315
rect 38630 6300 38654 6314
rect 38630 6294 38633 6300
rect 38648 6298 38654 6300
rect 38671 6298 38677 6315
rect 39346 6314 39360 6334
rect 39568 6332 39574 6349
rect 39591 6332 39597 6349
rect 39568 6329 39597 6332
rect 40717 6328 40720 6354
rect 40746 6348 40749 6354
rect 40764 6349 40793 6352
rect 40764 6348 40770 6349
rect 40746 6334 40770 6348
rect 40746 6328 40749 6334
rect 40764 6332 40770 6334
rect 40787 6332 40793 6349
rect 40764 6329 40793 6332
rect 40809 6314 40812 6320
rect 39346 6300 40812 6314
rect 38648 6295 38677 6298
rect 40809 6294 40812 6300
rect 40838 6294 40841 6320
rect 42014 6314 42028 6363
rect 42419 6362 42422 6368
rect 42448 6362 42451 6388
rect 42750 6382 42764 6402
rect 42658 6368 42764 6382
rect 42658 6314 42672 6368
rect 42879 6314 42882 6320
rect 42014 6300 42672 6314
rect 42859 6300 42882 6314
rect 42879 6294 42882 6300
rect 42908 6294 42911 6320
rect 43072 6314 43086 6402
rect 43110 6400 43116 6402
rect 43133 6400 43139 6417
rect 44774 6416 44788 6436
rect 45271 6430 45274 6436
rect 45300 6430 45303 6456
rect 45363 6430 45366 6456
rect 45392 6450 45395 6456
rect 49673 6450 49687 6470
rect 49733 6450 49736 6456
rect 45392 6436 49687 6450
rect 49713 6436 49736 6450
rect 45392 6430 45395 6436
rect 49733 6430 49736 6436
rect 49762 6430 49765 6456
rect 49963 6430 49966 6456
rect 49992 6430 49995 6456
rect 52309 6450 52312 6456
rect 52289 6436 52312 6450
rect 52309 6430 52312 6436
rect 52338 6430 52341 6456
rect 52355 6430 52358 6456
rect 52384 6450 52387 6456
rect 52384 6436 53068 6450
rect 52384 6430 52387 6436
rect 45087 6416 45090 6422
rect 44774 6402 45090 6416
rect 43110 6397 43139 6400
rect 45087 6396 45090 6402
rect 45116 6396 45119 6422
rect 45225 6416 45228 6422
rect 45181 6402 45228 6416
rect 45225 6396 45228 6402
rect 45254 6416 45257 6422
rect 45317 6416 45320 6422
rect 45254 6402 45320 6416
rect 45254 6396 45257 6402
rect 45317 6396 45320 6402
rect 45346 6396 45349 6422
rect 45640 6417 45669 6420
rect 45640 6400 45646 6417
rect 45663 6400 45669 6417
rect 45640 6397 45669 6400
rect 49274 6417 49303 6420
rect 49274 6400 49280 6417
rect 49297 6400 49303 6417
rect 52585 6416 52588 6422
rect 51405 6402 52588 6416
rect 49274 6397 49303 6400
rect 43247 6382 43250 6388
rect 43227 6368 43250 6382
rect 43247 6362 43250 6368
rect 43276 6362 43279 6388
rect 44121 6362 44124 6388
rect 44150 6382 44153 6388
rect 44812 6383 44841 6386
rect 44812 6382 44818 6383
rect 44150 6368 44818 6382
rect 44150 6362 44153 6368
rect 44812 6366 44818 6368
rect 44835 6382 44841 6383
rect 44857 6382 44860 6388
rect 44835 6368 44860 6382
rect 44835 6366 44841 6368
rect 44812 6363 44841 6366
rect 44857 6362 44860 6368
rect 44886 6362 44889 6388
rect 44904 6383 44933 6386
rect 44904 6366 44910 6383
rect 44927 6382 44933 6383
rect 44927 6368 44972 6382
rect 44927 6366 44933 6368
rect 44904 6363 44933 6366
rect 44958 6320 44972 6368
rect 45041 6362 45044 6388
rect 45070 6382 45073 6388
rect 45648 6382 45662 6397
rect 45070 6368 45662 6382
rect 45070 6362 45073 6368
rect 49282 6348 49296 6397
rect 52585 6396 52588 6402
rect 52614 6396 52617 6422
rect 53054 6420 53068 6436
rect 53046 6417 53075 6420
rect 53046 6400 53052 6417
rect 53069 6400 53075 6417
rect 53046 6397 53075 6400
rect 49595 6382 49598 6388
rect 49551 6368 49598 6382
rect 49595 6362 49598 6368
rect 49624 6382 49627 6388
rect 50699 6382 50702 6388
rect 49624 6368 50702 6382
rect 49624 6362 49627 6368
rect 50699 6362 50702 6368
rect 50728 6362 50731 6388
rect 50837 6382 50840 6388
rect 50817 6368 50840 6382
rect 50837 6362 50840 6368
rect 50866 6362 50869 6388
rect 52402 6383 52431 6386
rect 52402 6366 52408 6383
rect 52425 6366 52431 6383
rect 52402 6363 52431 6366
rect 50470 6349 50499 6352
rect 49282 6334 49664 6348
rect 43891 6314 43894 6320
rect 43072 6300 43894 6314
rect 43891 6294 43894 6300
rect 43920 6294 43923 6320
rect 43983 6314 43986 6320
rect 43963 6300 43986 6314
rect 43983 6294 43986 6300
rect 44012 6294 44015 6320
rect 44213 6294 44216 6320
rect 44242 6314 44245 6320
rect 44582 6315 44611 6318
rect 44582 6314 44588 6315
rect 44242 6300 44588 6314
rect 44242 6294 44245 6300
rect 44582 6298 44588 6300
rect 44605 6298 44611 6315
rect 44949 6314 44952 6320
rect 44905 6300 44952 6314
rect 44582 6295 44611 6298
rect 44949 6294 44952 6300
rect 44978 6314 44981 6320
rect 45272 6315 45301 6318
rect 45272 6314 45278 6315
rect 44978 6300 45278 6314
rect 44978 6294 44981 6300
rect 45272 6298 45278 6300
rect 45295 6298 45301 6315
rect 45272 6295 45301 6298
rect 49182 6315 49211 6318
rect 49182 6298 49188 6315
rect 49205 6314 49211 6315
rect 49595 6314 49598 6320
rect 49205 6300 49598 6314
rect 49205 6298 49211 6300
rect 49182 6295 49211 6298
rect 49595 6294 49598 6300
rect 49624 6294 49627 6320
rect 49650 6314 49664 6334
rect 50470 6332 50476 6349
rect 50493 6348 50499 6349
rect 50515 6348 50518 6354
rect 50493 6334 50518 6348
rect 50493 6332 50499 6334
rect 50470 6329 50499 6332
rect 50515 6328 50518 6334
rect 50544 6328 50547 6354
rect 51619 6328 51622 6354
rect 51648 6348 51651 6354
rect 52410 6348 52424 6363
rect 52953 6348 52956 6354
rect 51648 6334 52424 6348
rect 52933 6334 52956 6348
rect 51648 6328 51651 6334
rect 52953 6328 52956 6334
rect 52982 6328 52985 6354
rect 54158 6348 54172 6470
rect 55713 6464 55716 6490
rect 55742 6484 55745 6490
rect 56128 6485 56157 6488
rect 56128 6484 56134 6485
rect 55742 6470 56134 6484
rect 55742 6464 55745 6470
rect 56128 6468 56134 6470
rect 56151 6484 56157 6485
rect 57277 6484 57280 6490
rect 56151 6470 57280 6484
rect 56151 6468 56157 6470
rect 56128 6465 56157 6468
rect 57277 6464 57280 6470
rect 57306 6464 57309 6490
rect 57369 6464 57372 6490
rect 57398 6484 57401 6490
rect 58703 6484 58706 6490
rect 57398 6470 58706 6484
rect 57398 6464 57401 6470
rect 58703 6464 58706 6470
rect 58732 6464 58735 6490
rect 59117 6484 59120 6490
rect 59097 6470 59120 6484
rect 59117 6464 59120 6470
rect 59146 6464 59149 6490
rect 59347 6484 59350 6490
rect 59327 6470 59350 6484
rect 59347 6464 59350 6470
rect 59376 6464 59379 6490
rect 63350 6485 63379 6488
rect 63350 6468 63356 6485
rect 63373 6484 63379 6485
rect 63441 6484 63444 6490
rect 63373 6470 63444 6484
rect 63373 6468 63379 6470
rect 63350 6465 63379 6468
rect 63441 6464 63444 6470
rect 63470 6464 63473 6490
rect 64039 6484 64042 6490
rect 64019 6470 64042 6484
rect 64039 6464 64042 6470
rect 64068 6464 64071 6490
rect 64315 6464 64318 6490
rect 64344 6484 64347 6490
rect 64362 6485 64391 6488
rect 64362 6484 64368 6485
rect 64344 6470 64368 6484
rect 64344 6464 64347 6470
rect 64362 6468 64368 6470
rect 64385 6468 64391 6485
rect 64591 6484 64594 6490
rect 64571 6470 64594 6484
rect 64362 6465 64391 6468
rect 64591 6464 64594 6470
rect 64620 6464 64623 6490
rect 65144 6485 65173 6488
rect 65144 6468 65150 6485
rect 65167 6484 65173 6485
rect 66661 6484 66664 6490
rect 65167 6470 66664 6484
rect 65167 6468 65173 6470
rect 65144 6465 65173 6468
rect 66661 6464 66664 6470
rect 66690 6464 66693 6490
rect 66754 6485 66783 6488
rect 66754 6468 66760 6485
rect 66777 6484 66783 6485
rect 66777 6470 66914 6484
rect 66777 6468 66783 6470
rect 66754 6465 66783 6468
rect 54793 6430 54796 6456
rect 54822 6450 54825 6456
rect 56174 6451 56203 6454
rect 56174 6450 56180 6451
rect 54822 6436 56180 6450
rect 54822 6430 54825 6436
rect 56174 6434 56180 6436
rect 56197 6434 56203 6451
rect 57002 6451 57031 6454
rect 57002 6450 57008 6451
rect 56174 6431 56203 6434
rect 56274 6436 57008 6450
rect 56274 6386 56288 6436
rect 57002 6434 57008 6436
rect 57025 6450 57031 6451
rect 57830 6451 57859 6454
rect 57025 6436 57806 6450
rect 57025 6434 57031 6436
rect 57002 6431 57031 6434
rect 56541 6416 56544 6422
rect 56521 6402 56544 6416
rect 56541 6396 56544 6402
rect 56570 6396 56573 6422
rect 56909 6416 56912 6422
rect 56889 6402 56912 6416
rect 56909 6396 56912 6402
rect 56938 6396 56941 6422
rect 57323 6396 57326 6422
rect 57352 6416 57355 6422
rect 57792 6416 57806 6436
rect 57830 6434 57836 6451
rect 57853 6450 57859 6451
rect 57875 6450 57878 6456
rect 57853 6436 57878 6450
rect 57853 6434 57859 6436
rect 57830 6431 57859 6434
rect 57875 6430 57878 6436
rect 57904 6430 57907 6456
rect 58657 6430 58660 6456
rect 58686 6430 58689 6456
rect 63257 6430 63260 6456
rect 63286 6450 63289 6456
rect 64600 6450 64614 6464
rect 66201 6450 66204 6456
rect 63286 6436 64614 6450
rect 66171 6436 66204 6450
rect 63286 6430 63289 6436
rect 57352 6402 57374 6416
rect 57792 6402 57944 6416
rect 57352 6396 57355 6402
rect 57930 6388 57944 6402
rect 59025 6396 59028 6422
rect 59054 6416 59057 6422
rect 63450 6420 63464 6436
rect 66201 6430 66204 6436
rect 66230 6430 66233 6456
rect 66799 6450 66802 6456
rect 66779 6436 66802 6450
rect 66799 6430 66802 6436
rect 66828 6430 66831 6456
rect 66900 6450 66914 6470
rect 66937 6464 66940 6490
rect 66966 6484 66969 6490
rect 67168 6485 67197 6488
rect 67168 6484 67174 6485
rect 66966 6470 67174 6484
rect 66966 6464 66969 6470
rect 67168 6468 67174 6470
rect 67191 6468 67197 6485
rect 67168 6465 67197 6468
rect 72734 6485 72763 6488
rect 72734 6468 72740 6485
rect 72757 6484 72763 6485
rect 73837 6484 73840 6490
rect 72757 6470 73840 6484
rect 72757 6468 72763 6470
rect 72734 6465 72763 6468
rect 73837 6464 73840 6470
rect 73866 6464 73869 6490
rect 75724 6485 75753 6488
rect 74076 6470 74918 6484
rect 67075 6450 67078 6456
rect 66900 6436 67078 6450
rect 67075 6430 67078 6436
rect 67104 6430 67107 6456
rect 71537 6430 71540 6456
rect 71566 6450 71569 6456
rect 72963 6450 72966 6456
rect 71566 6436 72894 6450
rect 72943 6436 72966 6450
rect 71566 6430 71569 6436
rect 59440 6417 59469 6420
rect 59440 6416 59446 6417
rect 59054 6402 59446 6416
rect 59054 6396 59057 6402
rect 59440 6400 59446 6402
rect 59463 6400 59469 6417
rect 59440 6397 59469 6400
rect 63442 6417 63471 6420
rect 63442 6400 63448 6417
rect 63465 6400 63471 6417
rect 63717 6416 63720 6422
rect 63697 6402 63720 6416
rect 63442 6397 63471 6400
rect 63717 6396 63720 6402
rect 63746 6416 63749 6422
rect 64132 6417 64161 6420
rect 63746 6402 64108 6416
rect 63746 6396 63749 6402
rect 56266 6383 56295 6386
rect 56266 6366 56272 6383
rect 56289 6366 56295 6383
rect 56266 6363 56295 6366
rect 56588 6383 56617 6386
rect 56588 6366 56594 6383
rect 56611 6382 56617 6383
rect 56955 6382 56958 6388
rect 56611 6368 56958 6382
rect 56611 6366 56617 6368
rect 56588 6363 56617 6366
rect 56955 6362 56958 6368
rect 56984 6362 56987 6388
rect 57369 6362 57372 6388
rect 57398 6362 57401 6388
rect 57829 6362 57832 6388
rect 57858 6382 57861 6388
rect 57876 6383 57905 6386
rect 57876 6382 57882 6383
rect 57858 6368 57882 6382
rect 57858 6362 57861 6368
rect 57876 6366 57882 6368
rect 57899 6366 57905 6383
rect 57876 6363 57905 6366
rect 57921 6362 57924 6388
rect 57950 6382 57953 6388
rect 58244 6383 58273 6386
rect 57950 6368 57972 6382
rect 57950 6362 57953 6368
rect 58244 6366 58250 6383
rect 58267 6366 58273 6383
rect 58381 6382 58384 6388
rect 58361 6368 58384 6382
rect 58244 6363 58273 6366
rect 57378 6348 57392 6362
rect 54158 6334 57392 6348
rect 57415 6328 57418 6354
rect 57444 6348 57447 6354
rect 58252 6348 58266 6363
rect 58381 6362 58384 6368
rect 58410 6362 58413 6388
rect 63763 6382 63766 6388
rect 58896 6368 63766 6382
rect 57444 6334 58266 6348
rect 57444 6328 57447 6334
rect 50377 6314 50380 6320
rect 49650 6300 50380 6314
rect 50377 6294 50380 6300
rect 50406 6294 50409 6320
rect 51527 6294 51530 6320
rect 51556 6314 51559 6320
rect 51574 6315 51603 6318
rect 51574 6314 51580 6315
rect 51556 6300 51580 6314
rect 51556 6294 51559 6300
rect 51574 6298 51580 6300
rect 51597 6298 51603 6315
rect 51574 6295 51603 6298
rect 51803 6294 51806 6320
rect 51832 6314 51835 6320
rect 52126 6315 52155 6318
rect 52126 6314 52132 6315
rect 51832 6300 52132 6314
rect 51832 6294 51835 6300
rect 52126 6298 52132 6300
rect 52149 6298 52155 6315
rect 55943 6314 55946 6320
rect 55923 6300 55946 6314
rect 52126 6295 52155 6298
rect 55943 6294 55946 6300
rect 55972 6294 55975 6320
rect 56541 6294 56544 6320
rect 56570 6314 56573 6320
rect 57369 6314 57372 6320
rect 56570 6300 57372 6314
rect 56570 6294 56573 6300
rect 57369 6294 57372 6300
rect 57398 6294 57401 6320
rect 57646 6315 57675 6318
rect 57646 6298 57652 6315
rect 57669 6314 57675 6315
rect 57921 6314 57924 6320
rect 57669 6300 57924 6314
rect 57669 6298 57675 6300
rect 57646 6295 57675 6298
rect 57921 6294 57924 6300
rect 57950 6294 57953 6320
rect 58252 6314 58266 6334
rect 58896 6314 58910 6368
rect 63763 6362 63766 6368
rect 63792 6362 63795 6388
rect 58252 6300 58910 6314
rect 63764 6315 63793 6318
rect 63764 6298 63770 6315
rect 63787 6314 63793 6315
rect 64039 6314 64042 6320
rect 63787 6300 64042 6314
rect 63787 6298 63793 6300
rect 63764 6295 63793 6298
rect 64039 6294 64042 6300
rect 64068 6294 64071 6320
rect 64094 6314 64108 6402
rect 64132 6400 64138 6417
rect 64155 6400 64161 6417
rect 64545 6416 64548 6422
rect 64525 6402 64548 6416
rect 64132 6397 64161 6400
rect 64140 6348 64154 6397
rect 64545 6396 64548 6402
rect 64574 6396 64577 6422
rect 65098 6417 65127 6420
rect 65098 6416 65104 6417
rect 64600 6402 65104 6416
rect 64177 6362 64180 6388
rect 64206 6382 64209 6388
rect 64600 6382 64614 6402
rect 65098 6400 65104 6402
rect 65121 6400 65127 6417
rect 65098 6397 65127 6400
rect 65143 6396 65146 6422
rect 65172 6416 65175 6422
rect 65420 6417 65449 6420
rect 65420 6416 65426 6417
rect 65172 6402 65426 6416
rect 65172 6396 65175 6402
rect 65420 6400 65426 6402
rect 65443 6400 65449 6417
rect 65420 6397 65449 6400
rect 64206 6368 64614 6382
rect 64684 6383 64713 6386
rect 64206 6362 64209 6368
rect 64684 6366 64690 6383
rect 64707 6382 64713 6383
rect 64867 6382 64870 6388
rect 64707 6368 64870 6382
rect 64707 6366 64713 6368
rect 64684 6363 64713 6366
rect 64867 6362 64870 6368
rect 64896 6362 64899 6388
rect 65557 6382 65560 6388
rect 65537 6368 65560 6382
rect 65557 6362 65560 6368
rect 65586 6362 65589 6388
rect 66293 6362 66296 6388
rect 66322 6382 66325 6388
rect 66808 6382 66822 6430
rect 66845 6396 66848 6422
rect 66874 6418 66877 6422
rect 66874 6416 66914 6418
rect 67260 6417 67289 6420
rect 67260 6416 67266 6417
rect 66874 6404 67266 6416
rect 66874 6396 66877 6404
rect 66900 6402 67266 6404
rect 67260 6400 67266 6402
rect 67283 6400 67289 6417
rect 67260 6397 67289 6400
rect 67674 6417 67703 6420
rect 67674 6400 67680 6417
rect 67697 6416 67703 6417
rect 71492 6417 71521 6420
rect 71492 6416 71498 6417
rect 67697 6402 71498 6416
rect 67697 6400 67703 6402
rect 67674 6397 67703 6400
rect 71492 6400 71498 6402
rect 71515 6416 71521 6417
rect 72880 6416 72894 6436
rect 72963 6430 72966 6436
rect 72992 6430 72995 6456
rect 74076 6450 74090 6470
rect 73018 6436 74090 6450
rect 74904 6450 74918 6470
rect 75724 6468 75730 6485
rect 75747 6484 75753 6485
rect 76321 6484 76324 6490
rect 75747 6470 76324 6484
rect 75747 6468 75753 6470
rect 75724 6465 75753 6468
rect 76321 6464 76324 6470
rect 76350 6464 76353 6490
rect 76368 6485 76397 6488
rect 76368 6468 76374 6485
rect 76391 6484 76397 6485
rect 76413 6484 76416 6490
rect 76391 6470 76416 6484
rect 76391 6468 76397 6470
rect 76368 6465 76397 6468
rect 76413 6464 76416 6470
rect 76442 6484 76445 6490
rect 76552 6485 76581 6488
rect 76552 6484 76558 6485
rect 76442 6470 76558 6484
rect 76442 6464 76445 6470
rect 76552 6468 76558 6470
rect 76575 6484 76581 6485
rect 76736 6485 76765 6488
rect 76736 6484 76742 6485
rect 76575 6470 76742 6484
rect 76575 6468 76581 6470
rect 76552 6465 76581 6468
rect 76736 6468 76742 6470
rect 76759 6484 76765 6485
rect 76920 6485 76949 6488
rect 76920 6484 76926 6485
rect 76759 6470 76926 6484
rect 76759 6468 76765 6470
rect 76736 6465 76765 6468
rect 76920 6468 76926 6470
rect 76943 6484 76949 6485
rect 77104 6485 77133 6488
rect 77104 6484 77110 6485
rect 76943 6470 77110 6484
rect 76943 6468 76949 6470
rect 76920 6465 76949 6468
rect 77104 6468 77110 6470
rect 77127 6484 77133 6485
rect 77472 6485 77501 6488
rect 77472 6484 77478 6485
rect 77127 6470 77478 6484
rect 77127 6468 77133 6470
rect 77104 6465 77133 6468
rect 77472 6468 77478 6470
rect 77495 6484 77501 6485
rect 78024 6485 78053 6488
rect 78024 6484 78030 6485
rect 77495 6470 78030 6484
rect 77495 6468 77501 6470
rect 77472 6465 77501 6468
rect 78024 6468 78030 6470
rect 78047 6484 78053 6485
rect 78208 6485 78237 6488
rect 78208 6484 78214 6485
rect 78047 6470 78214 6484
rect 78047 6468 78053 6470
rect 78024 6465 78053 6468
rect 78208 6468 78214 6470
rect 78231 6484 78237 6485
rect 78392 6485 78421 6488
rect 78392 6484 78398 6485
rect 78231 6470 78398 6484
rect 78231 6468 78237 6470
rect 78208 6465 78237 6468
rect 78392 6468 78398 6470
rect 78415 6484 78421 6485
rect 78575 6484 78578 6490
rect 78415 6470 78578 6484
rect 78415 6468 78421 6470
rect 78392 6465 78421 6468
rect 78575 6464 78578 6470
rect 78604 6464 78607 6490
rect 79311 6464 79314 6490
rect 79340 6484 79343 6490
rect 81749 6484 81752 6490
rect 79340 6470 81752 6484
rect 79340 6464 79343 6470
rect 78299 6450 78302 6456
rect 74904 6436 78302 6450
rect 72917 6416 72920 6422
rect 71515 6402 72848 6416
rect 72873 6402 72920 6416
rect 71515 6400 71521 6402
rect 71492 6397 71521 6400
rect 66322 6368 66822 6382
rect 66892 6383 66921 6386
rect 66322 6362 66325 6368
rect 66892 6366 66898 6383
rect 66915 6366 66921 6383
rect 71629 6382 71632 6388
rect 71609 6368 71632 6382
rect 66892 6363 66921 6366
rect 65143 6348 65146 6354
rect 64140 6334 65146 6348
rect 65143 6328 65146 6334
rect 65172 6328 65175 6354
rect 66845 6348 66848 6354
rect 66233 6334 66848 6348
rect 66233 6314 66247 6334
rect 66845 6328 66848 6334
rect 66874 6328 66877 6354
rect 66569 6314 66572 6320
rect 64094 6300 66247 6314
rect 66549 6300 66572 6314
rect 66569 6294 66572 6300
rect 66598 6294 66601 6320
rect 66615 6294 66618 6320
rect 66644 6314 66647 6320
rect 66900 6314 66914 6363
rect 71629 6362 71632 6368
rect 71658 6362 71661 6388
rect 72834 6382 72848 6402
rect 72917 6396 72920 6402
rect 72946 6396 72949 6422
rect 73018 6416 73032 6436
rect 78299 6430 78302 6436
rect 78328 6430 78331 6456
rect 79634 6451 79663 6454
rect 79634 6450 79640 6451
rect 78653 6436 79640 6450
rect 72972 6402 73032 6416
rect 73516 6417 73545 6420
rect 72972 6382 72986 6402
rect 73516 6400 73522 6417
rect 73539 6416 73545 6417
rect 73653 6416 73656 6422
rect 73539 6402 73656 6416
rect 73539 6400 73545 6402
rect 73516 6397 73545 6400
rect 73653 6396 73656 6402
rect 73682 6396 73685 6422
rect 74451 6402 74504 6416
rect 74490 6388 74504 6402
rect 74665 6396 74668 6422
rect 74694 6416 74697 6422
rect 74942 6417 74971 6420
rect 74942 6416 74948 6417
rect 74694 6402 74948 6416
rect 74694 6396 74697 6402
rect 74942 6400 74948 6402
rect 74965 6416 74971 6417
rect 74965 6402 75194 6416
rect 74965 6400 74971 6402
rect 74942 6397 74971 6400
rect 72834 6368 72986 6382
rect 73056 6383 73085 6386
rect 73056 6366 73062 6383
rect 73079 6382 73085 6383
rect 73699 6382 73702 6388
rect 73079 6368 73702 6382
rect 73079 6366 73085 6368
rect 73056 6363 73085 6366
rect 73699 6362 73702 6368
rect 73728 6362 73731 6388
rect 73746 6383 73775 6386
rect 73746 6366 73752 6383
rect 73769 6366 73775 6383
rect 73883 6382 73886 6388
rect 73863 6368 73886 6382
rect 73746 6363 73775 6366
rect 66937 6328 66940 6354
rect 66966 6348 66969 6354
rect 67766 6349 67795 6352
rect 67766 6348 67772 6349
rect 66966 6334 67772 6348
rect 66966 6328 66969 6334
rect 67766 6332 67772 6334
rect 67789 6332 67795 6349
rect 67766 6329 67795 6332
rect 72871 6328 72874 6354
rect 72900 6348 72903 6354
rect 73754 6348 73768 6363
rect 73883 6362 73886 6368
rect 73912 6362 73915 6388
rect 74481 6362 74484 6388
rect 74510 6362 74513 6388
rect 74619 6382 74622 6388
rect 74599 6368 74622 6382
rect 74619 6362 74622 6368
rect 74648 6362 74651 6388
rect 75180 6354 75194 6402
rect 75217 6396 75220 6422
rect 75246 6416 75249 6422
rect 77426 6417 77455 6420
rect 77426 6416 77432 6417
rect 75246 6402 77432 6416
rect 75246 6396 75249 6402
rect 77426 6400 77432 6402
rect 77449 6400 77455 6417
rect 77426 6397 77455 6400
rect 77931 6396 77934 6422
rect 77960 6416 77963 6422
rect 78653 6416 78667 6436
rect 79634 6434 79640 6436
rect 79657 6434 79663 6451
rect 80185 6450 80188 6456
rect 79634 6431 79663 6434
rect 79964 6436 80188 6450
rect 77960 6402 78667 6416
rect 77960 6396 77963 6402
rect 78897 6396 78900 6422
rect 78926 6416 78929 6422
rect 79588 6417 79617 6420
rect 79588 6416 79594 6417
rect 78926 6402 79594 6416
rect 78926 6396 78929 6402
rect 79588 6400 79594 6402
rect 79611 6416 79617 6417
rect 79964 6416 79978 6436
rect 80185 6430 80188 6436
rect 80214 6430 80217 6456
rect 80562 6436 80898 6450
rect 79611 6402 79978 6416
rect 80002 6417 80031 6420
rect 79611 6400 79617 6402
rect 79588 6397 79617 6400
rect 80002 6400 80008 6417
rect 80025 6416 80031 6417
rect 80562 6416 80576 6436
rect 80025 6402 80576 6416
rect 80600 6417 80629 6420
rect 80025 6400 80031 6402
rect 80002 6397 80031 6400
rect 80600 6400 80606 6417
rect 80623 6416 80629 6417
rect 80829 6416 80832 6422
rect 80623 6402 80832 6416
rect 80623 6400 80629 6402
rect 80600 6397 80629 6400
rect 80829 6396 80832 6402
rect 80858 6396 80861 6422
rect 75769 6382 75772 6388
rect 75749 6368 75772 6382
rect 75769 6362 75772 6368
rect 75798 6362 75801 6388
rect 75862 6383 75891 6386
rect 75862 6366 75868 6383
rect 75885 6366 75891 6383
rect 75862 6363 75891 6366
rect 72900 6334 73768 6348
rect 72900 6328 72903 6334
rect 75171 6328 75174 6354
rect 75200 6348 75203 6354
rect 75815 6348 75818 6354
rect 75200 6334 75818 6348
rect 75200 6328 75203 6334
rect 75815 6328 75818 6334
rect 75844 6328 75847 6354
rect 66644 6300 66914 6314
rect 73424 6315 73453 6318
rect 66644 6294 66647 6300
rect 73424 6298 73430 6315
rect 73447 6314 73453 6315
rect 74251 6314 74254 6320
rect 73447 6300 74254 6314
rect 73447 6298 73453 6300
rect 73424 6295 73453 6298
rect 74251 6294 74254 6300
rect 74280 6294 74283 6320
rect 74987 6314 74990 6320
rect 74967 6300 74990 6314
rect 74987 6294 74990 6300
rect 75016 6294 75019 6320
rect 75540 6315 75569 6318
rect 75540 6298 75546 6315
rect 75563 6314 75569 6315
rect 75631 6314 75634 6320
rect 75563 6300 75634 6314
rect 75563 6298 75569 6300
rect 75540 6295 75569 6298
rect 75631 6294 75634 6300
rect 75660 6294 75663 6320
rect 75677 6294 75680 6320
rect 75706 6314 75709 6320
rect 75870 6314 75884 6363
rect 76367 6362 76370 6388
rect 76396 6382 76399 6388
rect 76396 6368 77494 6382
rect 76396 6362 76399 6368
rect 76184 6349 76213 6352
rect 76184 6332 76190 6349
rect 76207 6348 76213 6349
rect 76413 6348 76416 6354
rect 76207 6334 76416 6348
rect 76207 6332 76213 6334
rect 76184 6329 76213 6332
rect 76413 6328 76416 6334
rect 76442 6328 76445 6354
rect 76551 6328 76554 6354
rect 76580 6348 76583 6354
rect 77242 6349 77271 6352
rect 77242 6348 77248 6349
rect 76580 6334 77248 6348
rect 76580 6328 76583 6334
rect 77242 6332 77248 6334
rect 77265 6332 77271 6349
rect 77480 6348 77494 6368
rect 77517 6362 77520 6388
rect 77546 6382 77549 6388
rect 79725 6382 79728 6388
rect 77546 6368 77568 6382
rect 77618 6368 79656 6382
rect 79705 6368 79728 6382
rect 77546 6362 77549 6368
rect 77618 6348 77632 6368
rect 79403 6348 79406 6354
rect 77480 6334 77632 6348
rect 79383 6334 79406 6348
rect 77242 6329 77271 6332
rect 79403 6328 79406 6334
rect 79432 6328 79435 6354
rect 79642 6348 79656 6368
rect 79725 6362 79728 6368
rect 79754 6362 79757 6388
rect 79771 6362 79774 6388
rect 79800 6382 79803 6388
rect 80783 6382 80786 6388
rect 79800 6368 80786 6382
rect 79800 6362 79803 6368
rect 80783 6362 80786 6368
rect 80812 6362 80815 6388
rect 80094 6349 80123 6352
rect 80094 6348 80100 6349
rect 79642 6334 80100 6348
rect 80094 6332 80100 6334
rect 80117 6332 80123 6349
rect 80094 6329 80123 6332
rect 77057 6314 77060 6320
rect 75706 6300 77060 6314
rect 75706 6294 75709 6300
rect 77057 6294 77060 6300
rect 77086 6314 77089 6320
rect 78943 6314 78946 6320
rect 77086 6300 78946 6314
rect 77086 6294 77089 6300
rect 78943 6294 78946 6300
rect 78972 6294 78975 6320
rect 80139 6294 80142 6320
rect 80168 6314 80171 6320
rect 80646 6315 80675 6318
rect 80646 6314 80652 6315
rect 80168 6300 80652 6314
rect 80168 6294 80171 6300
rect 80646 6298 80652 6300
rect 80669 6298 80675 6315
rect 80884 6314 80898 6436
rect 80930 6420 80944 6470
rect 81749 6464 81752 6470
rect 81778 6464 81781 6490
rect 81796 6485 81825 6488
rect 81796 6468 81802 6485
rect 81819 6468 81825 6485
rect 81796 6465 81825 6468
rect 82210 6485 82239 6488
rect 82210 6468 82216 6485
rect 82233 6484 82239 6485
rect 82623 6484 82626 6490
rect 82233 6470 82626 6484
rect 82233 6468 82239 6470
rect 82210 6465 82239 6468
rect 81703 6450 81706 6456
rect 81673 6436 81706 6450
rect 81703 6430 81706 6436
rect 81732 6430 81735 6456
rect 81804 6450 81818 6465
rect 82623 6464 82626 6470
rect 82652 6484 82655 6490
rect 82652 6470 83497 6484
rect 82652 6464 82655 6470
rect 82256 6451 82285 6454
rect 82256 6450 82262 6451
rect 81804 6436 82262 6450
rect 80922 6417 80951 6420
rect 80922 6400 80928 6417
rect 80945 6400 80951 6417
rect 80922 6397 80951 6400
rect 81059 6382 81062 6388
rect 81039 6368 81062 6382
rect 81059 6362 81062 6368
rect 81088 6362 81091 6388
rect 81427 6362 81430 6388
rect 81456 6382 81459 6388
rect 81804 6382 81818 6436
rect 82256 6434 82262 6436
rect 82279 6450 82285 6451
rect 83483 6450 83497 6470
rect 83589 6464 83592 6490
rect 83618 6484 83621 6490
rect 83912 6485 83941 6488
rect 83912 6484 83918 6485
rect 83618 6470 83918 6484
rect 83618 6464 83621 6470
rect 83912 6468 83918 6470
rect 83935 6468 83941 6485
rect 87499 6484 87502 6490
rect 87479 6470 87502 6484
rect 83912 6465 83941 6468
rect 87499 6464 87502 6470
rect 87528 6464 87531 6490
rect 87822 6485 87851 6488
rect 87822 6468 87828 6485
rect 87845 6484 87851 6485
rect 87867 6484 87870 6490
rect 87845 6470 87870 6484
rect 87845 6468 87851 6470
rect 87822 6465 87851 6468
rect 87867 6464 87870 6470
rect 87896 6464 87899 6490
rect 88189 6464 88192 6490
rect 88218 6484 88221 6490
rect 90075 6484 90078 6490
rect 88218 6470 90078 6484
rect 88218 6464 88221 6470
rect 82279 6436 83336 6450
rect 83483 6436 84026 6450
rect 82279 6434 82285 6436
rect 82256 6431 82285 6434
rect 82670 6417 82699 6420
rect 82670 6400 82676 6417
rect 82693 6416 82699 6417
rect 82715 6416 82718 6422
rect 82693 6402 82718 6416
rect 82693 6400 82699 6402
rect 82670 6397 82699 6400
rect 82715 6396 82718 6402
rect 82744 6396 82747 6422
rect 83083 6396 83086 6422
rect 83112 6416 83115 6422
rect 83267 6416 83270 6422
rect 83112 6402 83270 6416
rect 83112 6396 83115 6402
rect 83267 6396 83270 6402
rect 83296 6396 83299 6422
rect 83322 6416 83336 6436
rect 84012 6420 84026 6436
rect 86901 6430 86904 6456
rect 86930 6450 86933 6456
rect 86930 6436 87936 6450
rect 86930 6430 86933 6436
rect 87922 6420 87936 6436
rect 87959 6430 87962 6456
rect 87988 6450 87991 6456
rect 88465 6450 88468 6456
rect 87988 6436 88468 6450
rect 87988 6430 87991 6436
rect 88465 6430 88468 6436
rect 88494 6430 88497 6456
rect 88971 6450 88974 6456
rect 88941 6436 88974 6450
rect 88971 6430 88974 6436
rect 89000 6430 89003 6456
rect 83682 6417 83711 6420
rect 83682 6416 83688 6417
rect 83322 6402 83688 6416
rect 83682 6400 83688 6402
rect 83705 6400 83711 6417
rect 83682 6397 83711 6400
rect 84004 6417 84033 6420
rect 84004 6400 84010 6417
rect 84027 6400 84033 6417
rect 84004 6397 84033 6400
rect 87592 6417 87621 6420
rect 87592 6400 87598 6417
rect 87615 6400 87621 6417
rect 87592 6397 87621 6400
rect 87914 6417 87943 6420
rect 87914 6400 87920 6417
rect 87937 6400 87943 6417
rect 88189 6416 88192 6422
rect 88169 6402 88192 6416
rect 87914 6397 87943 6400
rect 82301 6382 82304 6388
rect 81456 6368 81818 6382
rect 82281 6368 82304 6382
rect 81456 6362 81459 6368
rect 82301 6362 82304 6368
rect 82330 6362 82333 6388
rect 81804 6334 82094 6348
rect 81804 6314 81818 6334
rect 80884 6300 81818 6314
rect 80646 6295 80675 6298
rect 81841 6294 81844 6320
rect 81870 6314 81873 6320
rect 82026 6315 82055 6318
rect 82026 6314 82032 6315
rect 81870 6300 82032 6314
rect 81870 6294 81873 6300
rect 82026 6298 82032 6300
rect 82049 6298 82055 6315
rect 82080 6314 82094 6334
rect 82117 6328 82120 6354
rect 82146 6348 82149 6354
rect 83590 6349 83619 6352
rect 83590 6348 83596 6349
rect 82146 6334 83596 6348
rect 82146 6328 82149 6334
rect 83590 6332 83596 6334
rect 83613 6332 83619 6349
rect 87600 6348 87614 6397
rect 88189 6396 88192 6402
rect 88218 6396 88221 6422
rect 89302 6420 89316 6470
rect 90075 6464 90078 6470
rect 90104 6464 90107 6490
rect 90121 6464 90124 6490
rect 90150 6484 90153 6490
rect 90398 6485 90427 6488
rect 90398 6484 90404 6485
rect 90150 6470 90404 6484
rect 90150 6464 90153 6470
rect 90398 6468 90404 6470
rect 90421 6468 90427 6485
rect 94169 6484 94172 6490
rect 90398 6465 90427 6468
rect 94040 6470 94172 6484
rect 90812 6451 90841 6454
rect 90812 6450 90818 6451
rect 90130 6436 90818 6450
rect 89294 6417 89323 6420
rect 89294 6400 89300 6417
rect 89317 6400 89323 6417
rect 90130 6416 90144 6436
rect 90812 6434 90818 6436
rect 90835 6434 90841 6451
rect 90812 6431 90841 6434
rect 89999 6402 90144 6416
rect 89294 6397 89323 6400
rect 90167 6396 90170 6422
rect 90196 6416 90199 6422
rect 90490 6417 90519 6420
rect 90490 6416 90496 6417
rect 90196 6402 90496 6416
rect 90196 6396 90199 6402
rect 90490 6400 90496 6402
rect 90513 6400 90519 6417
rect 90765 6416 90768 6422
rect 90721 6402 90768 6416
rect 90490 6397 90519 6400
rect 90765 6396 90768 6402
rect 90794 6416 90797 6422
rect 94040 6420 94054 6470
rect 94169 6464 94172 6470
rect 94198 6484 94201 6490
rect 95687 6484 95690 6490
rect 94198 6470 95690 6484
rect 94198 6464 94201 6470
rect 95687 6464 95690 6470
rect 95716 6484 95719 6490
rect 96148 6485 96177 6488
rect 96148 6484 96154 6485
rect 95716 6470 96154 6484
rect 95716 6464 95719 6470
rect 96148 6468 96154 6470
rect 96171 6468 96177 6485
rect 96148 6465 96177 6468
rect 96239 6464 96242 6490
rect 96268 6484 96271 6490
rect 96268 6470 96722 6484
rect 96268 6464 96271 6470
rect 94261 6430 94264 6456
rect 94290 6450 94293 6456
rect 94768 6451 94797 6454
rect 94768 6450 94774 6451
rect 94290 6436 94774 6450
rect 94290 6430 94293 6436
rect 94768 6434 94774 6436
rect 94791 6450 94797 6451
rect 95457 6450 95460 6456
rect 94791 6436 95227 6450
rect 95437 6436 95460 6450
rect 94791 6434 94797 6436
rect 94768 6431 94797 6434
rect 91088 6417 91117 6420
rect 91088 6416 91094 6417
rect 90794 6402 91094 6416
rect 90794 6396 90797 6402
rect 91088 6400 91094 6402
rect 91111 6400 91117 6417
rect 91088 6397 91117 6400
rect 94032 6417 94061 6420
rect 94032 6400 94038 6417
rect 94055 6400 94061 6417
rect 94032 6397 94061 6400
rect 94169 6396 94172 6422
rect 94198 6416 94201 6422
rect 94308 6417 94337 6420
rect 94308 6416 94314 6417
rect 94198 6402 94314 6416
rect 94198 6396 94201 6402
rect 94308 6400 94314 6402
rect 94331 6416 94337 6417
rect 94399 6416 94402 6422
rect 94331 6402 94402 6416
rect 94331 6400 94337 6402
rect 94308 6397 94337 6400
rect 94399 6396 94402 6402
rect 94428 6396 94431 6422
rect 94675 6416 94678 6422
rect 94655 6402 94678 6416
rect 94675 6396 94678 6402
rect 94704 6396 94707 6422
rect 88328 6383 88357 6386
rect 88328 6366 88334 6383
rect 88351 6382 88357 6383
rect 88373 6382 88376 6388
rect 88351 6368 88376 6382
rect 88351 6366 88357 6368
rect 88328 6363 88357 6366
rect 88373 6362 88376 6368
rect 88402 6362 88405 6388
rect 89432 6383 89461 6386
rect 89432 6366 89438 6383
rect 89455 6382 89461 6383
rect 89455 6368 90052 6382
rect 89455 6366 89461 6368
rect 89432 6363 89461 6366
rect 90038 6348 90052 6368
rect 90075 6362 90078 6388
rect 90104 6382 90107 6388
rect 94767 6382 94770 6388
rect 90104 6368 94770 6382
rect 90104 6362 90107 6368
rect 94767 6362 94770 6368
rect 94796 6362 94799 6388
rect 95213 6382 95227 6436
rect 95457 6430 95460 6436
rect 95486 6430 95489 6456
rect 95871 6430 95874 6456
rect 95900 6450 95903 6456
rect 96654 6451 96683 6454
rect 96654 6450 96660 6451
rect 95900 6436 96660 6450
rect 95900 6430 95903 6436
rect 96654 6434 96660 6436
rect 96677 6434 96683 6451
rect 96708 6450 96722 6470
rect 96975 6464 96978 6490
rect 97004 6484 97007 6490
rect 97435 6484 97438 6490
rect 97004 6470 97438 6484
rect 97004 6464 97007 6470
rect 97435 6464 97438 6470
rect 97464 6484 97467 6490
rect 97987 6484 97990 6490
rect 97464 6470 97990 6484
rect 97464 6464 97467 6470
rect 97987 6464 97990 6470
rect 98016 6464 98019 6490
rect 98861 6464 98864 6490
rect 98890 6484 98893 6490
rect 98890 6470 103254 6484
rect 98890 6464 98893 6470
rect 97942 6451 97971 6454
rect 97942 6450 97948 6451
rect 96708 6436 96899 6450
rect 97536 6436 97948 6450
rect 96654 6431 96683 6434
rect 97536 6422 97550 6436
rect 97942 6434 97948 6436
rect 97965 6434 97971 6451
rect 101483 6450 101486 6456
rect 97942 6431 97971 6434
rect 101262 6436 101486 6450
rect 95504 6417 95533 6420
rect 95504 6400 95510 6417
rect 95527 6416 95533 6417
rect 96102 6417 96131 6420
rect 96102 6416 96108 6417
rect 95527 6402 96108 6416
rect 95527 6400 95533 6402
rect 95504 6397 95533 6400
rect 96102 6400 96108 6402
rect 96125 6416 96131 6417
rect 96285 6416 96288 6422
rect 96125 6402 96288 6416
rect 96125 6400 96131 6402
rect 96102 6397 96131 6400
rect 96285 6396 96288 6402
rect 96314 6396 96317 6422
rect 97527 6416 97530 6422
rect 97507 6402 97530 6416
rect 97527 6396 97530 6402
rect 97556 6396 97559 6422
rect 98677 6416 98680 6422
rect 98657 6402 98680 6416
rect 98677 6396 98680 6402
rect 98706 6396 98709 6422
rect 98723 6396 98726 6422
rect 98752 6416 98755 6422
rect 99183 6416 99186 6422
rect 98752 6402 99068 6416
rect 99163 6402 99186 6416
rect 98752 6396 98755 6402
rect 95596 6383 95625 6386
rect 95596 6382 95602 6383
rect 95213 6368 95602 6382
rect 95596 6366 95602 6368
rect 95619 6382 95625 6383
rect 96194 6383 96223 6386
rect 96194 6382 96200 6383
rect 95619 6368 96200 6382
rect 95619 6366 95625 6368
rect 95596 6363 95625 6366
rect 96194 6366 96200 6368
rect 96217 6382 96223 6383
rect 96331 6382 96334 6388
rect 96217 6368 96334 6382
rect 96217 6366 96223 6368
rect 96194 6363 96223 6366
rect 96331 6362 96334 6368
rect 96360 6362 96363 6388
rect 96515 6382 96518 6388
rect 96495 6368 96518 6382
rect 96515 6362 96518 6368
rect 96544 6362 96547 6388
rect 97389 6382 97392 6388
rect 96570 6368 97392 6382
rect 90121 6348 90124 6354
rect 87600 6334 88074 6348
rect 90038 6334 90124 6348
rect 83590 6329 83619 6332
rect 82716 6315 82745 6318
rect 82716 6314 82722 6315
rect 82080 6300 82722 6314
rect 82026 6295 82055 6298
rect 82716 6298 82722 6300
rect 82739 6314 82745 6315
rect 83083 6314 83086 6320
rect 82739 6300 83086 6314
rect 82739 6298 82745 6300
rect 82716 6295 82745 6298
rect 83083 6294 83086 6300
rect 83112 6294 83115 6320
rect 83313 6314 83316 6320
rect 83293 6300 83316 6314
rect 83313 6294 83316 6300
rect 83342 6294 83345 6320
rect 88060 6314 88074 6334
rect 90121 6328 90124 6334
rect 90150 6328 90153 6354
rect 90259 6328 90262 6354
rect 90288 6348 90291 6354
rect 91041 6348 91044 6354
rect 90288 6334 91044 6348
rect 90288 6328 90291 6334
rect 91041 6328 91044 6334
rect 91070 6328 91073 6354
rect 93940 6349 93969 6352
rect 93940 6332 93946 6349
rect 93963 6348 93969 6349
rect 94307 6348 94310 6354
rect 93963 6334 94310 6348
rect 93963 6332 93969 6334
rect 93940 6329 93969 6332
rect 94307 6328 94310 6334
rect 94336 6328 94339 6354
rect 94583 6328 94586 6354
rect 94612 6348 94615 6354
rect 95871 6348 95874 6354
rect 94612 6334 95874 6348
rect 94612 6328 94615 6334
rect 95871 6328 95874 6334
rect 95900 6328 95903 6354
rect 95963 6328 95966 6354
rect 95992 6348 95995 6354
rect 96239 6348 96242 6354
rect 95992 6334 96242 6348
rect 95992 6328 95995 6334
rect 96239 6328 96242 6334
rect 96268 6328 96271 6354
rect 96570 6348 96584 6368
rect 97389 6362 97392 6368
rect 97418 6362 97421 6388
rect 97895 6362 97898 6388
rect 97924 6382 97927 6388
rect 98080 6383 98109 6386
rect 98080 6382 98086 6383
rect 97924 6368 98086 6382
rect 97924 6362 97927 6368
rect 98080 6366 98086 6368
rect 98103 6382 98109 6383
rect 98815 6382 98818 6388
rect 98103 6368 98818 6382
rect 98103 6366 98109 6368
rect 98080 6363 98109 6366
rect 98815 6362 98818 6368
rect 98844 6362 98847 6388
rect 99054 6386 99068 6402
rect 99183 6396 99186 6402
rect 99212 6396 99215 6422
rect 100242 6417 100271 6420
rect 100242 6400 100248 6417
rect 100265 6416 100271 6417
rect 100333 6416 100336 6422
rect 100265 6402 100336 6416
rect 100265 6400 100271 6402
rect 100242 6397 100271 6400
rect 100333 6396 100336 6402
rect 100362 6396 100365 6422
rect 100655 6416 100658 6422
rect 100635 6402 100658 6416
rect 100655 6396 100658 6402
rect 100684 6396 100687 6422
rect 99046 6383 99075 6386
rect 99046 6366 99052 6383
rect 99069 6382 99075 6383
rect 99275 6382 99278 6388
rect 99069 6368 99278 6382
rect 99069 6366 99075 6368
rect 99046 6363 99075 6366
rect 99275 6362 99278 6368
rect 99304 6382 99307 6388
rect 100195 6382 100198 6388
rect 99304 6368 100198 6382
rect 99304 6362 99307 6368
rect 100195 6362 100198 6368
rect 100224 6362 100227 6388
rect 100288 6383 100317 6386
rect 100288 6366 100294 6383
rect 100311 6382 100317 6383
rect 101262 6382 101276 6436
rect 101483 6430 101486 6436
rect 101512 6430 101515 6456
rect 101667 6430 101670 6456
rect 101696 6430 101699 6456
rect 102412 6420 102426 6470
rect 102817 6430 102820 6456
rect 102846 6430 102849 6456
rect 102404 6417 102433 6420
rect 102404 6400 102410 6417
rect 102427 6400 102433 6417
rect 103240 6416 103254 6470
rect 103277 6464 103280 6490
rect 103306 6484 103309 6490
rect 103691 6484 103694 6490
rect 103306 6470 103694 6484
rect 103306 6464 103309 6470
rect 103691 6464 103694 6470
rect 103720 6464 103723 6490
rect 103921 6464 103924 6490
rect 103950 6484 103953 6490
rect 103950 6470 109878 6484
rect 103950 6464 103953 6470
rect 103332 6436 103806 6450
rect 103332 6416 103346 6436
rect 103240 6402 103346 6416
rect 103738 6417 103767 6420
rect 102404 6397 102433 6400
rect 103738 6400 103744 6417
rect 103761 6400 103767 6417
rect 103738 6397 103767 6400
rect 100311 6368 101276 6382
rect 101300 6383 101329 6386
rect 100311 6366 100317 6368
rect 100288 6363 100317 6366
rect 101300 6366 101306 6383
rect 101323 6366 101329 6383
rect 101437 6382 101440 6388
rect 101417 6368 101440 6382
rect 101300 6363 101329 6366
rect 101069 6348 101072 6354
rect 96294 6334 96584 6348
rect 97168 6334 101072 6348
rect 88695 6314 88698 6320
rect 88060 6300 88698 6314
rect 88695 6294 88698 6300
rect 88724 6294 88727 6320
rect 88925 6294 88928 6320
rect 88954 6314 88957 6320
rect 89064 6315 89093 6318
rect 89064 6314 89070 6315
rect 88954 6300 89070 6314
rect 88954 6294 88957 6300
rect 89064 6298 89070 6300
rect 89087 6298 89093 6315
rect 89064 6295 89093 6298
rect 89937 6294 89940 6320
rect 89966 6314 89969 6320
rect 90168 6315 90197 6318
rect 90168 6314 90174 6315
rect 89966 6300 90174 6314
rect 89966 6294 89969 6300
rect 90168 6298 90174 6300
rect 90191 6314 90197 6315
rect 90305 6314 90308 6320
rect 90191 6300 90308 6314
rect 90191 6298 90197 6300
rect 90168 6295 90197 6298
rect 90305 6294 90308 6300
rect 90334 6294 90337 6320
rect 90719 6294 90722 6320
rect 90748 6314 90751 6320
rect 91134 6315 91163 6318
rect 91134 6314 91140 6315
rect 90748 6300 91140 6314
rect 90748 6294 90751 6300
rect 91134 6298 91140 6300
rect 91157 6298 91163 6315
rect 91134 6295 91163 6298
rect 93893 6294 93896 6320
rect 93922 6314 93925 6320
rect 94354 6315 94383 6318
rect 94354 6314 94360 6315
rect 93922 6300 94360 6314
rect 93922 6294 93925 6300
rect 94354 6298 94360 6300
rect 94377 6314 94383 6315
rect 94491 6314 94494 6320
rect 94377 6300 94494 6314
rect 94377 6298 94383 6300
rect 94354 6295 94383 6298
rect 94491 6294 94494 6300
rect 94520 6294 94523 6320
rect 95273 6314 95276 6320
rect 95253 6300 95276 6314
rect 95273 6294 95276 6300
rect 95302 6294 95305 6320
rect 95918 6315 95947 6318
rect 95918 6298 95924 6315
rect 95941 6314 95947 6315
rect 96009 6314 96012 6320
rect 95941 6300 96012 6314
rect 95941 6298 95947 6300
rect 95918 6295 95947 6298
rect 96009 6294 96012 6300
rect 96038 6294 96041 6320
rect 96055 6294 96058 6320
rect 96084 6314 96087 6320
rect 96294 6314 96308 6334
rect 96084 6300 96308 6314
rect 96084 6294 96087 6300
rect 96515 6294 96518 6320
rect 96544 6314 96547 6320
rect 97168 6314 97182 6334
rect 101069 6328 101072 6334
rect 101098 6348 101101 6354
rect 101308 6348 101322 6363
rect 101437 6362 101440 6368
rect 101466 6362 101469 6388
rect 101483 6362 101486 6388
rect 101512 6382 101515 6388
rect 102081 6382 102084 6388
rect 101512 6368 102084 6382
rect 101512 6362 101515 6368
rect 102081 6362 102084 6368
rect 102110 6362 102113 6388
rect 102541 6382 102544 6388
rect 102521 6368 102544 6382
rect 102541 6362 102544 6368
rect 102570 6362 102573 6388
rect 102587 6362 102590 6388
rect 102616 6382 102619 6388
rect 103746 6382 103760 6397
rect 102616 6368 103760 6382
rect 103792 6382 103806 6436
rect 105301 6430 105304 6456
rect 105330 6450 105333 6456
rect 109864 6450 109878 6470
rect 109901 6464 109904 6490
rect 109930 6484 109933 6490
rect 119101 6484 119104 6490
rect 109930 6470 119104 6484
rect 109930 6464 109933 6470
rect 114133 6450 114136 6456
rect 105330 6436 108682 6450
rect 109864 6436 114136 6450
rect 105330 6430 105333 6436
rect 103829 6396 103832 6422
rect 103858 6416 103861 6422
rect 105172 6416 105232 6418
rect 108291 6416 108294 6422
rect 103858 6404 108294 6416
rect 103858 6402 105186 6404
rect 105218 6402 108294 6404
rect 103858 6396 103861 6402
rect 108291 6396 108294 6402
rect 108320 6396 108323 6422
rect 108668 6416 108682 6436
rect 114133 6430 114136 6436
rect 114162 6430 114165 6456
rect 115191 6450 115194 6456
rect 114701 6436 115194 6450
rect 115191 6430 115194 6436
rect 115220 6430 115223 6456
rect 109901 6416 109904 6422
rect 108668 6402 109904 6416
rect 109901 6396 109904 6402
rect 109930 6396 109933 6422
rect 111833 6396 111836 6422
rect 111862 6416 111865 6422
rect 113352 6417 113381 6420
rect 113352 6416 113358 6417
rect 111862 6402 113358 6416
rect 111862 6396 111865 6402
rect 113352 6400 113358 6402
rect 113375 6400 113381 6417
rect 113352 6397 113381 6400
rect 113397 6396 113400 6422
rect 113426 6416 113429 6422
rect 113674 6417 113703 6420
rect 113674 6416 113680 6417
rect 113426 6402 113680 6416
rect 113426 6396 113429 6402
rect 113674 6400 113680 6402
rect 113697 6400 113703 6417
rect 113949 6416 113952 6422
rect 113929 6402 113952 6416
rect 113674 6397 113703 6400
rect 113949 6396 113952 6402
rect 113978 6396 113981 6422
rect 115145 6416 115148 6422
rect 115125 6402 115148 6416
rect 115145 6396 115148 6402
rect 115174 6396 115177 6422
rect 115384 6420 115398 6470
rect 119101 6464 119104 6470
rect 119130 6484 119133 6490
rect 125541 6484 125544 6490
rect 119130 6470 125544 6484
rect 119130 6464 119133 6470
rect 115513 6450 115516 6456
rect 115493 6436 115516 6450
rect 115513 6430 115516 6436
rect 115542 6430 115545 6456
rect 116157 6430 116160 6456
rect 116186 6450 116189 6456
rect 119147 6450 119150 6456
rect 116186 6436 119150 6450
rect 116186 6430 116189 6436
rect 119147 6430 119150 6436
rect 119176 6430 119179 6456
rect 119294 6450 119308 6470
rect 119248 6436 119308 6450
rect 119378 6451 119407 6454
rect 115376 6417 115405 6420
rect 115376 6400 115382 6417
rect 115399 6400 115405 6417
rect 116525 6416 116528 6422
rect 116081 6402 116364 6416
rect 116505 6402 116528 6416
rect 115376 6397 115405 6400
rect 113958 6382 113972 6396
rect 114088 6383 114117 6386
rect 114088 6382 114094 6383
rect 103792 6368 107647 6382
rect 102616 6362 102619 6368
rect 103645 6348 103648 6354
rect 101098 6334 101322 6348
rect 103240 6334 103392 6348
rect 103625 6334 103648 6348
rect 101098 6328 101101 6334
rect 96544 6300 97182 6314
rect 96544 6294 96547 6300
rect 97205 6294 97208 6320
rect 97234 6314 97237 6320
rect 97758 6315 97787 6318
rect 97758 6314 97764 6315
rect 97234 6300 97764 6314
rect 97234 6294 97237 6300
rect 97758 6298 97764 6300
rect 97781 6298 97787 6315
rect 97758 6295 97787 6298
rect 97987 6294 97990 6320
rect 98016 6314 98019 6320
rect 98494 6315 98523 6318
rect 98494 6314 98500 6315
rect 98016 6300 98500 6314
rect 98016 6294 98019 6300
rect 98494 6298 98500 6300
rect 98517 6298 98523 6315
rect 99091 6314 99094 6320
rect 99071 6300 99094 6314
rect 98494 6295 98523 6298
rect 99091 6294 99094 6300
rect 99120 6294 99123 6320
rect 100563 6314 100566 6320
rect 100543 6300 100566 6314
rect 100563 6294 100566 6300
rect 100592 6294 100595 6320
rect 100977 6294 100980 6320
rect 101006 6314 101009 6320
rect 102127 6314 102130 6320
rect 101006 6300 102130 6314
rect 101006 6294 101009 6300
rect 102127 6294 102130 6300
rect 102156 6294 102159 6320
rect 102174 6315 102203 6318
rect 102174 6298 102180 6315
rect 102197 6314 102203 6315
rect 102265 6314 102268 6320
rect 102197 6300 102268 6314
rect 102197 6298 102203 6300
rect 102174 6295 102203 6298
rect 102265 6294 102268 6300
rect 102294 6314 102297 6320
rect 102587 6314 102590 6320
rect 102294 6300 102590 6314
rect 102294 6294 102297 6300
rect 102587 6294 102590 6300
rect 102616 6294 102619 6320
rect 102633 6294 102636 6320
rect 102662 6314 102665 6320
rect 103240 6314 103254 6334
rect 102662 6300 103254 6314
rect 103378 6314 103392 6334
rect 103645 6328 103648 6334
rect 103674 6328 103677 6354
rect 105301 6314 105304 6320
rect 103378 6300 105304 6314
rect 102662 6294 102665 6300
rect 105301 6294 105304 6300
rect 105330 6294 105333 6320
rect 107633 6314 107647 6368
rect 109864 6368 113972 6382
rect 114004 6368 114094 6382
rect 109864 6314 109878 6368
rect 109901 6328 109904 6354
rect 109930 6348 109933 6354
rect 113582 6349 113611 6352
rect 109930 6334 113558 6348
rect 109930 6328 109933 6334
rect 107633 6300 109878 6314
rect 113260 6315 113289 6318
rect 113260 6298 113266 6315
rect 113283 6314 113289 6315
rect 113443 6314 113446 6320
rect 113283 6300 113446 6314
rect 113283 6298 113289 6300
rect 113260 6295 113289 6298
rect 113443 6294 113446 6300
rect 113472 6294 113475 6320
rect 113544 6314 113558 6334
rect 113582 6332 113588 6349
rect 113605 6348 113611 6349
rect 114004 6348 114018 6368
rect 114088 6366 114094 6368
rect 114111 6366 114117 6383
rect 114088 6363 114117 6366
rect 114133 6362 114136 6388
rect 114162 6382 114165 6388
rect 115099 6382 115102 6388
rect 114162 6368 115102 6382
rect 114162 6362 114165 6368
rect 115099 6362 115102 6368
rect 115128 6362 115131 6388
rect 116350 6382 116364 6402
rect 116525 6396 116528 6402
rect 116554 6396 116557 6422
rect 118503 6416 118506 6422
rect 118483 6402 118506 6416
rect 118503 6396 118506 6402
rect 118532 6396 118535 6422
rect 118826 6417 118855 6420
rect 118826 6400 118832 6417
rect 118849 6416 118855 6417
rect 119193 6416 119196 6422
rect 118849 6402 119196 6416
rect 118849 6400 118855 6402
rect 118826 6397 118855 6400
rect 119193 6396 119196 6402
rect 119222 6396 119225 6422
rect 119248 6420 119262 6436
rect 119378 6434 119384 6451
rect 119401 6450 119407 6451
rect 119515 6450 119518 6456
rect 119401 6436 119518 6450
rect 119401 6434 119407 6436
rect 119378 6431 119407 6434
rect 119515 6430 119518 6436
rect 119544 6430 119547 6456
rect 120021 6450 120024 6456
rect 119991 6436 120024 6450
rect 120021 6430 120024 6436
rect 120050 6430 120053 6456
rect 120352 6420 120366 6470
rect 125541 6464 125544 6470
rect 125570 6464 125573 6490
rect 126186 6485 126215 6488
rect 126186 6468 126192 6485
rect 126209 6484 126215 6485
rect 127335 6484 127338 6490
rect 126209 6470 127338 6484
rect 126209 6468 126215 6470
rect 126186 6465 126215 6468
rect 127335 6464 127338 6470
rect 127364 6464 127367 6490
rect 128117 6464 128120 6490
rect 128146 6484 128149 6490
rect 132303 6484 132306 6490
rect 128146 6470 131797 6484
rect 132283 6470 132306 6484
rect 128146 6464 128149 6470
rect 120481 6450 120484 6456
rect 120461 6436 120484 6450
rect 120481 6430 120484 6436
rect 120510 6430 120513 6456
rect 122321 6450 122324 6456
rect 122123 6436 122324 6450
rect 119240 6417 119269 6420
rect 119240 6400 119246 6417
rect 119263 6400 119269 6417
rect 119240 6397 119269 6400
rect 120344 6417 120373 6420
rect 120344 6400 120350 6417
rect 120367 6400 120373 6417
rect 120344 6397 120373 6400
rect 121033 6396 121036 6422
rect 121062 6396 121065 6422
rect 121125 6396 121128 6422
rect 121154 6416 121157 6422
rect 121908 6417 121937 6420
rect 121908 6416 121914 6417
rect 121154 6402 121914 6416
rect 121154 6396 121157 6402
rect 121908 6400 121914 6402
rect 121931 6416 121937 6417
rect 122123 6416 122137 6436
rect 122321 6430 122324 6436
rect 122350 6430 122353 6456
rect 122459 6430 122462 6456
rect 122488 6450 122491 6456
rect 122644 6451 122673 6454
rect 122644 6450 122650 6451
rect 122488 6436 122650 6450
rect 122488 6430 122491 6436
rect 122644 6434 122650 6436
rect 122667 6434 122673 6451
rect 122644 6431 122673 6434
rect 122689 6430 122692 6456
rect 122718 6450 122721 6456
rect 125680 6451 125709 6454
rect 125680 6450 125686 6451
rect 122718 6436 125686 6450
rect 122718 6430 122721 6436
rect 125680 6434 125686 6436
rect 125703 6450 125709 6451
rect 125817 6450 125820 6456
rect 125703 6436 125820 6450
rect 125703 6434 125709 6436
rect 125680 6431 125709 6434
rect 125817 6430 125820 6436
rect 125846 6430 125849 6456
rect 126231 6430 126234 6456
rect 126260 6450 126263 6456
rect 128623 6450 128626 6456
rect 126260 6436 126282 6450
rect 127581 6436 128370 6450
rect 126260 6430 126263 6436
rect 122275 6416 122278 6422
rect 121931 6402 122137 6416
rect 122255 6402 122278 6416
rect 121931 6400 121937 6402
rect 121908 6397 121937 6400
rect 122275 6396 122278 6402
rect 122304 6396 122307 6422
rect 122368 6417 122397 6420
rect 122368 6400 122374 6417
rect 122391 6416 122397 6417
rect 122413 6416 122416 6422
rect 122391 6402 122416 6416
rect 122391 6400 122397 6402
rect 122368 6397 122397 6400
rect 122413 6396 122416 6402
rect 122442 6416 122445 6422
rect 122598 6417 122627 6420
rect 122598 6416 122604 6417
rect 122442 6402 122604 6416
rect 122442 6396 122445 6402
rect 122598 6400 122604 6402
rect 122621 6400 122627 6417
rect 122598 6397 122627 6400
rect 125174 6417 125203 6420
rect 125174 6400 125180 6417
rect 125197 6416 125203 6417
rect 125587 6416 125590 6422
rect 125197 6402 125590 6416
rect 125197 6400 125203 6402
rect 125174 6397 125203 6400
rect 125573 6396 125590 6402
rect 125616 6396 125619 6422
rect 125771 6416 125774 6422
rect 125751 6402 125774 6416
rect 125771 6396 125774 6402
rect 125800 6396 125803 6422
rect 125826 6415 126208 6416
rect 126240 6415 126254 6430
rect 125826 6402 126254 6415
rect 116572 6383 116601 6386
rect 116572 6382 116578 6383
rect 115154 6368 116042 6382
rect 116350 6368 116578 6382
rect 115154 6348 115168 6368
rect 113605 6334 114018 6348
rect 114602 6334 115168 6348
rect 116028 6348 116042 6368
rect 116572 6366 116578 6368
rect 116595 6366 116601 6383
rect 125573 6382 125587 6396
rect 125826 6382 125840 6402
rect 126194 6401 126254 6402
rect 128118 6417 128147 6420
rect 128118 6400 128124 6417
rect 128141 6416 128147 6417
rect 128301 6416 128304 6422
rect 128141 6402 128304 6416
rect 128141 6400 128147 6402
rect 128118 6397 128147 6400
rect 128301 6396 128304 6402
rect 128330 6396 128333 6422
rect 116572 6363 116601 6366
rect 117293 6368 120274 6382
rect 117293 6348 117307 6368
rect 116028 6334 117307 6348
rect 118734 6349 118763 6352
rect 113605 6332 113611 6334
rect 113582 6329 113611 6332
rect 114602 6314 114616 6334
rect 118734 6332 118740 6349
rect 118757 6348 118763 6349
rect 118917 6348 118920 6354
rect 118757 6334 118920 6348
rect 118757 6332 118763 6334
rect 118734 6329 118763 6332
rect 118917 6328 118920 6334
rect 118946 6328 118949 6354
rect 118963 6328 118966 6354
rect 118992 6348 118995 6354
rect 118992 6334 119308 6348
rect 118992 6328 118995 6334
rect 113544 6300 114616 6314
rect 114777 6294 114780 6320
rect 114806 6314 114809 6320
rect 114824 6315 114853 6318
rect 114824 6314 114830 6315
rect 114806 6300 114830 6314
rect 114806 6294 114809 6300
rect 114824 6298 114830 6300
rect 114847 6298 114853 6315
rect 115053 6314 115056 6320
rect 115033 6300 115056 6314
rect 114824 6295 114853 6298
rect 115053 6294 115056 6300
rect 115082 6294 115085 6320
rect 115099 6294 115102 6320
rect 115128 6314 115131 6320
rect 116157 6314 116160 6320
rect 115128 6300 116160 6314
rect 115128 6294 115131 6300
rect 116157 6294 116160 6300
rect 116186 6294 116189 6320
rect 116249 6314 116252 6320
rect 116229 6300 116252 6314
rect 116249 6294 116252 6300
rect 116278 6314 116281 6320
rect 116571 6314 116574 6320
rect 116278 6300 116574 6314
rect 116278 6294 116281 6300
rect 116571 6294 116574 6300
rect 116600 6294 116603 6320
rect 118412 6315 118441 6318
rect 118412 6298 118418 6315
rect 118435 6314 118441 6315
rect 119239 6314 119242 6320
rect 118435 6300 119242 6314
rect 118435 6298 118441 6300
rect 118412 6295 118441 6298
rect 119239 6294 119242 6300
rect 119268 6294 119271 6320
rect 119294 6314 119308 6334
rect 119423 6314 119426 6320
rect 119294 6300 119426 6314
rect 119423 6294 119426 6300
rect 119452 6294 119455 6320
rect 119561 6294 119564 6320
rect 119590 6314 119593 6320
rect 120114 6315 120143 6318
rect 120114 6314 120120 6315
rect 119590 6300 120120 6314
rect 119590 6294 119593 6300
rect 120114 6298 120120 6300
rect 120137 6314 120143 6315
rect 120159 6314 120162 6320
rect 120137 6300 120162 6314
rect 120137 6298 120143 6300
rect 120114 6295 120143 6298
rect 120159 6294 120162 6300
rect 120188 6294 120191 6320
rect 120260 6314 120274 6368
rect 121042 6368 125150 6382
rect 125573 6368 125840 6382
rect 121042 6314 121056 6368
rect 121079 6328 121082 6354
rect 121108 6348 121111 6354
rect 121108 6334 122137 6348
rect 121108 6328 121111 6334
rect 121217 6314 121220 6320
rect 120260 6300 121056 6314
rect 121197 6300 121220 6314
rect 121217 6294 121220 6300
rect 121246 6294 121249 6320
rect 121447 6294 121450 6320
rect 121476 6314 121479 6320
rect 121954 6315 121983 6318
rect 121954 6314 121960 6315
rect 121476 6300 121960 6314
rect 121476 6294 121479 6300
rect 121954 6298 121960 6300
rect 121977 6298 121983 6315
rect 122123 6314 122137 6334
rect 122321 6328 122324 6354
rect 122350 6348 122353 6354
rect 124161 6348 124164 6354
rect 122350 6334 124164 6348
rect 122350 6328 122353 6334
rect 124161 6328 124164 6334
rect 124190 6328 124193 6354
rect 125081 6348 125084 6354
rect 125061 6334 125084 6348
rect 125081 6328 125084 6334
rect 125110 6328 125113 6354
rect 125136 6348 125150 6368
rect 126047 6362 126050 6388
rect 126076 6382 126079 6388
rect 126278 6383 126307 6386
rect 126278 6382 126284 6383
rect 126076 6368 126284 6382
rect 126076 6362 126079 6368
rect 126278 6366 126284 6368
rect 126301 6366 126307 6383
rect 126278 6363 126307 6366
rect 126829 6362 126832 6388
rect 126858 6382 126861 6388
rect 126858 6368 126880 6382
rect 126858 6362 126861 6368
rect 126967 6362 126970 6388
rect 126996 6382 126999 6388
rect 126996 6368 127018 6382
rect 126996 6362 126999 6368
rect 127565 6362 127568 6388
rect 127594 6382 127597 6388
rect 127704 6383 127733 6386
rect 127704 6382 127710 6383
rect 127594 6368 127710 6382
rect 127594 6362 127597 6368
rect 127704 6366 127710 6368
rect 127727 6382 127733 6383
rect 128163 6382 128166 6388
rect 127727 6368 128166 6382
rect 127727 6366 127733 6368
rect 127704 6363 127733 6366
rect 128163 6362 128166 6368
rect 128192 6362 128195 6388
rect 128209 6362 128212 6388
rect 128238 6382 128241 6388
rect 128238 6368 128260 6382
rect 128238 6362 128241 6368
rect 125909 6348 125912 6354
rect 125136 6334 125912 6348
rect 125909 6328 125912 6334
rect 125938 6328 125941 6354
rect 127519 6328 127522 6354
rect 127548 6348 127551 6354
rect 127934 6349 127963 6352
rect 127934 6348 127940 6349
rect 127548 6334 127940 6348
rect 127548 6328 127551 6334
rect 127934 6332 127940 6334
rect 127957 6332 127963 6349
rect 127934 6329 127963 6332
rect 125955 6314 125958 6320
rect 122123 6300 125958 6314
rect 121954 6295 121983 6298
rect 125955 6294 125958 6300
rect 125984 6294 125987 6320
rect 126001 6294 126004 6320
rect 126030 6314 126033 6320
rect 128356 6314 128370 6436
rect 128540 6436 128626 6450
rect 128540 6420 128554 6436
rect 128623 6430 128626 6436
rect 128652 6430 128655 6456
rect 130877 6450 130880 6456
rect 130833 6436 130880 6450
rect 130877 6430 130880 6436
rect 130906 6450 130909 6456
rect 131614 6451 131643 6454
rect 131614 6450 131620 6451
rect 130906 6436 131620 6450
rect 130906 6430 130909 6436
rect 131614 6434 131620 6436
rect 131637 6434 131643 6451
rect 131614 6431 131643 6434
rect 131659 6430 131662 6456
rect 131688 6450 131691 6456
rect 131706 6451 131735 6454
rect 131706 6450 131712 6451
rect 131688 6436 131712 6450
rect 131688 6430 131691 6436
rect 131706 6434 131712 6436
rect 131729 6434 131735 6451
rect 131783 6450 131797 6470
rect 132303 6464 132306 6470
rect 132332 6464 132335 6490
rect 134189 6484 134192 6490
rect 132634 6470 134192 6484
rect 132634 6450 132648 6470
rect 134189 6464 134192 6470
rect 134218 6464 134221 6490
rect 151301 6484 151304 6490
rect 134244 6470 148357 6484
rect 151281 6470 151304 6484
rect 132763 6450 132766 6456
rect 131783 6436 132648 6450
rect 132743 6436 132766 6450
rect 131706 6431 131735 6434
rect 128532 6417 128561 6420
rect 128532 6400 128538 6417
rect 128555 6400 128561 6417
rect 128532 6397 128561 6400
rect 130923 6396 130926 6422
rect 130952 6416 130955 6422
rect 131246 6417 131275 6420
rect 131246 6416 131252 6417
rect 130952 6402 131252 6416
rect 130952 6396 130955 6402
rect 131246 6400 131252 6402
rect 131269 6400 131275 6417
rect 131246 6397 131275 6400
rect 132074 6417 132103 6420
rect 132074 6400 132080 6417
rect 132097 6416 132103 6417
rect 132165 6416 132168 6422
rect 132097 6402 132168 6416
rect 132097 6400 132103 6402
rect 132074 6397 132103 6400
rect 132165 6396 132168 6402
rect 132194 6396 132197 6422
rect 132211 6396 132214 6422
rect 132240 6416 132243 6422
rect 132634 6420 132648 6436
rect 132763 6430 132766 6436
rect 132792 6430 132795 6456
rect 133269 6430 133272 6456
rect 133298 6430 133301 6456
rect 134244 6450 134258 6470
rect 135523 6450 135526 6456
rect 133416 6436 134258 6450
rect 135309 6436 135526 6450
rect 132396 6417 132425 6420
rect 132396 6416 132402 6417
rect 132240 6402 132402 6416
rect 132240 6396 132243 6402
rect 132396 6400 132402 6402
rect 132419 6400 132425 6417
rect 132396 6397 132425 6400
rect 132626 6417 132655 6420
rect 132626 6400 132632 6417
rect 132649 6400 132655 6417
rect 132626 6397 132655 6400
rect 128577 6362 128580 6388
rect 128606 6382 128609 6388
rect 131153 6382 131156 6388
rect 128606 6368 131156 6382
rect 128606 6362 128609 6368
rect 131153 6362 131156 6368
rect 131182 6362 131185 6388
rect 133416 6382 133430 6436
rect 135523 6430 135526 6436
rect 135552 6430 135555 6456
rect 135891 6450 135894 6456
rect 135847 6436 135894 6450
rect 135891 6430 135894 6436
rect 135920 6450 135923 6456
rect 136397 6450 136400 6456
rect 135920 6436 136400 6450
rect 135920 6430 135923 6436
rect 136397 6430 136400 6436
rect 136426 6430 136429 6456
rect 136444 6451 136473 6454
rect 136444 6434 136450 6451
rect 136467 6450 136473 6451
rect 136581 6450 136584 6456
rect 136467 6436 136584 6450
rect 136467 6434 136473 6436
rect 136444 6431 136473 6434
rect 136581 6430 136584 6436
rect 136610 6430 136613 6456
rect 147943 6450 147946 6456
rect 141443 6436 147946 6450
rect 133914 6417 133943 6420
rect 133914 6400 133920 6417
rect 133937 6416 133943 6417
rect 134143 6416 134146 6422
rect 133937 6402 134146 6416
rect 133937 6400 133943 6402
rect 133914 6397 133943 6400
rect 134143 6396 134146 6402
rect 134172 6416 134175 6422
rect 134511 6416 134514 6422
rect 134172 6402 134514 6416
rect 134172 6396 134175 6402
rect 134511 6396 134514 6402
rect 134540 6396 134543 6422
rect 134558 6417 134587 6420
rect 134558 6400 134564 6417
rect 134581 6400 134587 6417
rect 134558 6397 134587 6400
rect 131714 6368 133430 6382
rect 128531 6328 128534 6354
rect 128560 6348 128563 6354
rect 131337 6348 131340 6354
rect 128560 6334 131268 6348
rect 131317 6334 131340 6348
rect 128560 6328 128563 6334
rect 128578 6315 128607 6318
rect 128578 6314 128584 6315
rect 126030 6300 126052 6314
rect 128356 6300 128584 6314
rect 126030 6294 126033 6300
rect 128578 6298 128584 6300
rect 128601 6298 128607 6315
rect 128578 6295 128607 6298
rect 130924 6315 130953 6318
rect 130924 6298 130930 6315
rect 130947 6314 130953 6315
rect 131107 6314 131110 6320
rect 130947 6300 131110 6314
rect 130947 6298 130953 6300
rect 130924 6295 130953 6298
rect 131107 6294 131110 6300
rect 131136 6294 131139 6320
rect 131254 6314 131268 6334
rect 131337 6328 131340 6334
rect 131366 6328 131369 6354
rect 131714 6314 131728 6368
rect 133499 6362 133502 6388
rect 133528 6382 133531 6388
rect 133775 6382 133778 6388
rect 133528 6368 133778 6382
rect 133528 6362 133531 6368
rect 133775 6362 133778 6368
rect 133804 6382 133807 6388
rect 133960 6383 133989 6386
rect 133960 6382 133966 6383
rect 133804 6368 133966 6382
rect 133804 6362 133807 6368
rect 133960 6366 133966 6368
rect 133983 6366 133989 6383
rect 133960 6363 133989 6366
rect 134005 6362 134008 6388
rect 134034 6382 134037 6388
rect 134034 6368 134056 6382
rect 134034 6362 134037 6368
rect 134189 6362 134192 6388
rect 134218 6382 134221 6388
rect 134566 6382 134580 6397
rect 135431 6396 135434 6422
rect 135460 6416 135463 6422
rect 135846 6417 135875 6420
rect 135846 6416 135852 6417
rect 135460 6402 135852 6416
rect 135460 6396 135463 6402
rect 135846 6400 135852 6402
rect 135869 6416 135875 6417
rect 136305 6416 136308 6422
rect 135869 6402 136308 6416
rect 135869 6400 135875 6402
rect 135846 6397 135875 6400
rect 136305 6396 136308 6402
rect 136334 6396 136337 6422
rect 141443 6416 141457 6436
rect 147943 6430 147946 6436
rect 147972 6430 147975 6456
rect 148343 6450 148357 6470
rect 151301 6464 151304 6470
rect 151330 6464 151333 6490
rect 152222 6485 152251 6488
rect 152222 6468 152228 6485
rect 152245 6484 152251 6485
rect 152681 6484 152684 6490
rect 152245 6470 152684 6484
rect 152245 6468 152251 6470
rect 152222 6465 152251 6468
rect 152681 6464 152684 6470
rect 152710 6464 152713 6490
rect 152497 6450 152500 6456
rect 148343 6436 152336 6450
rect 152477 6436 152500 6450
rect 145137 6416 145140 6422
rect 136360 6402 141457 6416
rect 143513 6402 145140 6416
rect 134695 6382 134698 6388
rect 134218 6368 134580 6382
rect 134675 6368 134698 6382
rect 134218 6362 134221 6368
rect 134695 6362 134698 6368
rect 134724 6362 134727 6388
rect 135984 6383 136013 6386
rect 135440 6368 135730 6382
rect 131751 6328 131754 6354
rect 131780 6348 131783 6354
rect 135440 6348 135454 6368
rect 131780 6334 132050 6348
rect 131780 6328 131783 6334
rect 131981 6314 131984 6320
rect 131254 6300 131728 6314
rect 131961 6300 131984 6314
rect 131981 6294 131984 6300
rect 132010 6294 132013 6320
rect 132036 6314 132050 6334
rect 133278 6334 134626 6348
rect 133278 6314 133292 6334
rect 133499 6314 133502 6320
rect 132036 6300 133292 6314
rect 133479 6300 133502 6314
rect 133499 6294 133502 6300
rect 133528 6294 133531 6320
rect 133545 6294 133548 6320
rect 133574 6314 133577 6320
rect 133730 6315 133759 6318
rect 133730 6314 133736 6315
rect 133574 6300 133736 6314
rect 133574 6294 133577 6300
rect 133730 6298 133736 6300
rect 133753 6298 133759 6315
rect 133730 6295 133759 6298
rect 133775 6294 133778 6320
rect 133804 6314 133807 6320
rect 134557 6314 134560 6320
rect 133804 6300 134560 6314
rect 133804 6294 133807 6300
rect 134557 6294 134560 6300
rect 134586 6294 134589 6320
rect 134612 6314 134626 6334
rect 135210 6334 135454 6348
rect 135716 6348 135730 6368
rect 135984 6366 135990 6383
rect 136007 6382 136013 6383
rect 136121 6382 136124 6388
rect 136007 6368 136124 6382
rect 136007 6366 136013 6368
rect 135984 6363 136013 6366
rect 136121 6362 136124 6368
rect 136150 6362 136153 6388
rect 136360 6348 136374 6402
rect 136443 6362 136446 6388
rect 136472 6382 136475 6388
rect 136490 6383 136519 6386
rect 136490 6382 136496 6383
rect 136472 6368 136496 6382
rect 136472 6362 136475 6368
rect 136490 6366 136496 6368
rect 136513 6366 136519 6383
rect 136490 6363 136519 6366
rect 136536 6383 136565 6386
rect 136536 6366 136542 6383
rect 136559 6366 136565 6383
rect 136536 6363 136565 6366
rect 135716 6334 136374 6348
rect 135210 6314 135224 6334
rect 136397 6328 136400 6354
rect 136426 6348 136429 6354
rect 136544 6348 136558 6363
rect 136581 6362 136584 6388
rect 136610 6382 136613 6388
rect 143513 6382 143527 6402
rect 145137 6396 145140 6402
rect 145166 6396 145169 6422
rect 151393 6416 151396 6422
rect 151373 6402 151396 6416
rect 151393 6396 151396 6402
rect 151422 6396 151425 6422
rect 152322 6420 152336 6436
rect 152497 6430 152500 6436
rect 152526 6450 152529 6456
rect 152727 6450 152730 6456
rect 152526 6436 152730 6450
rect 152526 6430 152529 6436
rect 152727 6430 152730 6436
rect 152756 6430 152759 6456
rect 152314 6417 152343 6420
rect 152314 6400 152320 6417
rect 152337 6400 152343 6417
rect 152314 6397 152343 6400
rect 136610 6368 143527 6382
rect 136610 6362 136613 6368
rect 136426 6334 136558 6348
rect 136426 6328 136429 6334
rect 135431 6314 135434 6320
rect 134612 6300 135224 6314
rect 135411 6300 135434 6314
rect 135431 6294 135434 6300
rect 135460 6294 135463 6320
rect 135569 6294 135572 6320
rect 135598 6314 135601 6320
rect 135662 6315 135691 6318
rect 135662 6314 135668 6315
rect 135598 6300 135668 6314
rect 135598 6294 135601 6300
rect 135662 6298 135668 6300
rect 135685 6298 135691 6315
rect 136259 6314 136262 6320
rect 136239 6300 136262 6314
rect 135662 6295 135691 6298
rect 136259 6294 136262 6300
rect 136288 6294 136291 6320
rect 136305 6294 136308 6320
rect 136334 6314 136337 6320
rect 140537 6314 140540 6320
rect 136334 6300 140540 6314
rect 136334 6294 136337 6300
rect 140537 6294 140540 6300
rect 140566 6294 140569 6320
rect 552 6269 152904 6280
rect 552 6243 19524 6269
rect 19550 6243 19556 6269
rect 19582 6243 19588 6269
rect 19614 6243 19620 6269
rect 19646 6243 19652 6269
rect 19678 6243 57623 6269
rect 57649 6243 57655 6269
rect 57681 6243 57687 6269
rect 57713 6243 57719 6269
rect 57745 6243 57751 6269
rect 57777 6243 95722 6269
rect 95748 6243 95754 6269
rect 95780 6243 95786 6269
rect 95812 6243 95818 6269
rect 95844 6243 95850 6269
rect 95876 6243 133821 6269
rect 133847 6243 133853 6269
rect 133879 6243 133885 6269
rect 133911 6243 133917 6269
rect 133943 6243 133949 6269
rect 133975 6243 152904 6269
rect 552 6232 152904 6243
rect 13485 6192 13488 6218
rect 13514 6212 13517 6218
rect 14037 6212 14040 6218
rect 13514 6198 14040 6212
rect 13514 6192 13517 6198
rect 14037 6192 14040 6198
rect 14066 6212 14069 6218
rect 14066 6198 14244 6212
rect 14066 6192 14069 6198
rect 7137 6158 7140 6184
rect 7166 6178 7169 6184
rect 14230 6178 14244 6198
rect 14405 6192 14408 6218
rect 14434 6212 14437 6218
rect 15648 6213 15677 6216
rect 15648 6212 15654 6213
rect 14434 6198 15654 6212
rect 14434 6192 14437 6198
rect 15648 6196 15654 6198
rect 15671 6196 15677 6213
rect 15648 6193 15677 6196
rect 16291 6192 16294 6218
rect 16320 6212 16323 6218
rect 16982 6213 17011 6216
rect 16320 6198 16544 6212
rect 16320 6192 16323 6198
rect 16530 6178 16544 6198
rect 16982 6196 16988 6213
rect 17005 6212 17011 6213
rect 17257 6212 17260 6218
rect 17005 6198 17260 6212
rect 17005 6196 17011 6198
rect 16982 6193 17011 6196
rect 17257 6192 17260 6198
rect 17286 6192 17289 6218
rect 17396 6213 17425 6216
rect 17396 6196 17402 6213
rect 17419 6212 17425 6213
rect 17993 6212 17996 6218
rect 17419 6198 17996 6212
rect 17419 6196 17425 6198
rect 17396 6193 17425 6196
rect 17993 6192 17996 6198
rect 18022 6192 18025 6218
rect 18592 6213 18621 6216
rect 18592 6196 18598 6213
rect 18615 6196 18621 6213
rect 18592 6193 18621 6196
rect 17441 6178 17444 6184
rect 7166 6164 14198 6178
rect 14230 6164 14474 6178
rect 16530 6164 17444 6178
rect 7166 6158 7169 6164
rect 13439 6144 13442 6150
rect 8480 6130 13442 6144
rect 2399 6022 2402 6048
rect 2428 6042 2431 6048
rect 8480 6042 8494 6130
rect 13439 6124 13442 6130
rect 13468 6124 13471 6150
rect 13854 6145 13883 6148
rect 13854 6128 13860 6145
rect 13877 6144 13883 6145
rect 14037 6144 14040 6150
rect 13877 6130 14040 6144
rect 13877 6128 13883 6130
rect 13854 6125 13883 6128
rect 14037 6124 14040 6130
rect 14066 6124 14069 6150
rect 14184 6144 14198 6164
rect 14359 6144 14362 6150
rect 14184 6130 14362 6144
rect 14359 6124 14362 6130
rect 14388 6124 14391 6150
rect 14460 6148 14474 6164
rect 17441 6158 17444 6164
rect 17470 6178 17473 6184
rect 18600 6178 18614 6193
rect 18913 6192 18916 6218
rect 18942 6212 18945 6218
rect 19236 6213 19265 6216
rect 19236 6212 19242 6213
rect 18942 6198 19242 6212
rect 18942 6192 18945 6198
rect 19236 6196 19242 6198
rect 19259 6196 19265 6213
rect 19236 6193 19265 6196
rect 19465 6192 19468 6218
rect 19494 6212 19497 6218
rect 19604 6213 19633 6216
rect 19604 6212 19610 6213
rect 19494 6198 19610 6212
rect 19494 6192 19497 6198
rect 19604 6196 19610 6198
rect 19627 6196 19633 6213
rect 19604 6193 19633 6196
rect 19695 6192 19698 6218
rect 19724 6212 19727 6218
rect 20477 6212 20480 6218
rect 19724 6198 20480 6212
rect 19724 6192 19727 6198
rect 20477 6192 20480 6198
rect 20506 6192 20509 6218
rect 21581 6212 21584 6218
rect 20762 6198 21512 6212
rect 21561 6198 21584 6212
rect 20762 6178 20776 6198
rect 17470 6164 18614 6178
rect 18646 6164 20776 6178
rect 21498 6178 21512 6198
rect 21581 6192 21584 6198
rect 21610 6192 21613 6218
rect 21903 6212 21906 6218
rect 21883 6198 21906 6212
rect 21903 6192 21906 6198
rect 21932 6192 21935 6218
rect 27009 6192 27012 6218
rect 27038 6212 27041 6218
rect 27056 6213 27085 6216
rect 27056 6212 27062 6213
rect 27038 6198 27062 6212
rect 27038 6192 27041 6198
rect 27056 6196 27062 6198
rect 27079 6196 27085 6213
rect 27056 6193 27085 6196
rect 27332 6213 27361 6216
rect 27332 6196 27338 6213
rect 27355 6212 27361 6213
rect 27745 6212 27748 6218
rect 27355 6198 27748 6212
rect 27355 6196 27361 6198
rect 27332 6193 27361 6196
rect 27745 6192 27748 6198
rect 27774 6192 27777 6218
rect 28343 6192 28346 6218
rect 28372 6212 28375 6218
rect 28666 6213 28695 6216
rect 28666 6212 28672 6213
rect 28372 6198 28672 6212
rect 28372 6192 28375 6198
rect 28666 6196 28672 6198
rect 28689 6196 28695 6213
rect 28987 6212 28990 6218
rect 28967 6198 28990 6212
rect 28666 6193 28695 6196
rect 28987 6192 28990 6198
rect 29016 6192 29019 6218
rect 37543 6192 37546 6218
rect 37572 6212 37575 6218
rect 37590 6213 37619 6216
rect 37590 6212 37596 6213
rect 37572 6198 37596 6212
rect 37572 6192 37575 6198
rect 37590 6196 37596 6198
rect 37613 6196 37619 6213
rect 39659 6212 39662 6218
rect 37590 6193 37619 6196
rect 37644 6198 39268 6212
rect 39639 6198 39662 6212
rect 21857 6178 21860 6184
rect 21498 6164 21860 6178
rect 17470 6158 17473 6164
rect 14452 6145 14481 6148
rect 14452 6128 14458 6145
rect 14475 6144 14481 6145
rect 14497 6144 14500 6150
rect 14475 6130 14500 6144
rect 14475 6128 14481 6130
rect 14452 6125 14481 6128
rect 14497 6124 14500 6130
rect 14526 6124 14529 6150
rect 14773 6144 14776 6150
rect 14729 6130 14776 6144
rect 14773 6124 14776 6130
rect 14802 6144 14805 6150
rect 15878 6145 15907 6148
rect 15878 6144 15884 6145
rect 14802 6130 15884 6144
rect 14802 6124 14805 6130
rect 15878 6128 15884 6130
rect 15901 6144 15907 6145
rect 15901 6130 17786 6144
rect 15901 6128 15907 6130
rect 15878 6125 15907 6128
rect 8517 6090 8520 6116
rect 8546 6110 8549 6116
rect 8546 6096 11047 6110
rect 8546 6090 8549 6096
rect 11033 6076 11047 6096
rect 13540 6096 13692 6110
rect 13540 6076 13554 6096
rect 11033 6062 13554 6076
rect 13678 6076 13692 6096
rect 13715 6090 13718 6116
rect 13744 6110 13747 6116
rect 14314 6111 14343 6114
rect 14314 6110 14320 6111
rect 13744 6096 13766 6110
rect 14000 6096 14320 6110
rect 13744 6090 13747 6096
rect 14000 6076 14014 6096
rect 14314 6094 14320 6096
rect 14337 6110 14343 6111
rect 14681 6110 14684 6116
rect 14337 6096 14684 6110
rect 14337 6094 14343 6096
rect 14314 6091 14343 6094
rect 14681 6090 14684 6096
rect 14710 6090 14713 6116
rect 17073 6110 17076 6116
rect 17053 6096 17076 6110
rect 17073 6090 17076 6096
rect 17102 6090 17105 6116
rect 17349 6110 17352 6116
rect 17305 6096 17352 6110
rect 17349 6090 17352 6096
rect 17378 6110 17381 6116
rect 17671 6110 17674 6116
rect 17378 6096 17674 6110
rect 17378 6090 17381 6096
rect 17671 6090 17674 6096
rect 17700 6090 17703 6116
rect 14727 6076 14730 6082
rect 13678 6062 14014 6076
rect 14138 6062 14730 6076
rect 13531 6042 13534 6048
rect 2428 6028 8494 6042
rect 13511 6028 13534 6042
rect 2428 6022 2431 6028
rect 13531 6022 13534 6028
rect 13560 6022 13563 6048
rect 13577 6022 13580 6048
rect 13606 6042 13609 6048
rect 13762 6043 13791 6046
rect 13762 6042 13768 6043
rect 13606 6028 13768 6042
rect 13606 6022 13609 6028
rect 13762 6026 13768 6028
rect 13785 6042 13791 6043
rect 13991 6042 13994 6048
rect 13785 6028 13994 6042
rect 13785 6026 13791 6028
rect 13762 6023 13791 6026
rect 13991 6022 13994 6028
rect 14020 6022 14023 6048
rect 14138 6046 14152 6062
rect 14727 6056 14730 6062
rect 14756 6056 14759 6082
rect 14911 6076 14914 6082
rect 14891 6062 14914 6076
rect 14911 6056 14914 6062
rect 14940 6056 14943 6082
rect 15601 6076 15604 6082
rect 15525 6062 15604 6076
rect 15601 6056 15604 6062
rect 15630 6056 15633 6082
rect 16015 6076 16018 6082
rect 15995 6062 16018 6076
rect 16015 6056 16018 6062
rect 16044 6056 16047 6082
rect 17718 6077 17747 6080
rect 17718 6076 17724 6077
rect 16629 6062 17724 6076
rect 17718 6060 17724 6062
rect 17741 6060 17747 6077
rect 17772 6076 17786 6130
rect 18178 6111 18207 6114
rect 18178 6094 18184 6111
rect 18201 6110 18207 6111
rect 18546 6111 18575 6114
rect 18546 6110 18552 6111
rect 18201 6096 18552 6110
rect 18201 6094 18207 6096
rect 18178 6091 18207 6094
rect 18546 6094 18552 6096
rect 18569 6110 18575 6111
rect 18646 6110 18660 6164
rect 21857 6158 21860 6164
rect 21886 6158 21889 6184
rect 37644 6178 37658 6198
rect 26834 6164 37658 6178
rect 20432 6145 20461 6148
rect 20432 6128 20438 6145
rect 20455 6144 20461 6145
rect 20477 6144 20480 6150
rect 20455 6130 20480 6144
rect 20455 6128 20461 6130
rect 20432 6125 20461 6128
rect 20477 6124 20480 6130
rect 20506 6124 20509 6150
rect 26182 6145 26211 6148
rect 26182 6144 26188 6145
rect 20716 6130 26188 6144
rect 18569 6096 18660 6110
rect 18569 6094 18575 6096
rect 18546 6091 18575 6094
rect 19005 6090 19008 6116
rect 19034 6110 19037 6116
rect 19328 6111 19357 6114
rect 19328 6110 19334 6111
rect 19034 6096 19334 6110
rect 19034 6090 19037 6096
rect 19328 6094 19334 6096
rect 19351 6094 19357 6111
rect 19328 6091 19357 6094
rect 19558 6111 19587 6114
rect 19558 6094 19564 6111
rect 19581 6110 19587 6111
rect 20155 6110 20158 6116
rect 19581 6096 20158 6110
rect 19581 6094 19587 6096
rect 19558 6091 19587 6094
rect 20155 6090 20158 6096
rect 20184 6090 20187 6116
rect 20293 6110 20296 6116
rect 20273 6096 20296 6110
rect 20293 6090 20296 6096
rect 20322 6090 20325 6116
rect 20716 6114 20730 6130
rect 26182 6128 26188 6130
rect 26205 6144 26211 6145
rect 26834 6144 26848 6164
rect 38003 6158 38006 6184
rect 38032 6178 38035 6184
rect 38601 6178 38604 6184
rect 38032 6164 38604 6178
rect 38032 6158 38035 6164
rect 26205 6130 26848 6144
rect 26205 6128 26211 6130
rect 26182 6125 26211 6128
rect 26917 6124 26920 6150
rect 26946 6124 26949 6150
rect 27838 6145 27867 6148
rect 27838 6144 27844 6145
rect 27593 6130 27844 6144
rect 20708 6111 20737 6114
rect 20708 6094 20714 6111
rect 20731 6094 20737 6111
rect 21857 6110 21860 6116
rect 21837 6096 21860 6110
rect 20708 6091 20737 6094
rect 20716 6076 20730 6091
rect 21857 6090 21860 6096
rect 21886 6110 21889 6116
rect 26926 6110 26940 6124
rect 27286 6111 27315 6114
rect 27286 6110 27292 6111
rect 21886 6096 24157 6110
rect 26926 6096 27292 6110
rect 21886 6090 21889 6096
rect 17772 6062 20730 6076
rect 17718 6057 17747 6060
rect 20799 6056 20802 6082
rect 20828 6076 20831 6082
rect 20846 6077 20875 6080
rect 20846 6076 20852 6077
rect 20828 6062 20852 6076
rect 20828 6056 20831 6062
rect 20846 6060 20852 6062
rect 20869 6060 20875 6077
rect 20846 6057 20875 6060
rect 20891 6056 20894 6082
rect 20920 6076 20923 6082
rect 20920 6062 21091 6076
rect 20920 6056 20923 6062
rect 14130 6043 14159 6046
rect 14130 6026 14136 6043
rect 14153 6026 14159 6043
rect 14130 6023 14159 6026
rect 14451 6022 14454 6048
rect 14480 6042 14483 6048
rect 15555 6042 15558 6048
rect 14480 6028 15558 6042
rect 14480 6022 14483 6028
rect 15555 6022 15558 6028
rect 15584 6022 15587 6048
rect 16153 6022 16156 6048
rect 16182 6042 16185 6048
rect 16475 6042 16478 6048
rect 16182 6028 16478 6042
rect 16182 6022 16185 6028
rect 16475 6022 16478 6028
rect 16504 6042 16507 6048
rect 16752 6043 16781 6046
rect 16752 6042 16758 6043
rect 16504 6028 16758 6042
rect 16504 6022 16507 6028
rect 16752 6026 16758 6028
rect 16775 6026 16781 6043
rect 18223 6042 18226 6048
rect 18203 6028 18226 6042
rect 16752 6023 16781 6026
rect 18223 6022 18226 6028
rect 18252 6022 18255 6048
rect 20110 6043 20139 6046
rect 20110 6026 20116 6043
rect 20133 6042 20139 6043
rect 20247 6042 20250 6048
rect 20133 6028 20250 6042
rect 20133 6026 20139 6028
rect 20110 6023 20139 6026
rect 20247 6022 20250 6028
rect 20276 6022 20279 6048
rect 20339 6042 20342 6048
rect 20319 6028 20342 6042
rect 20339 6022 20342 6028
rect 20368 6022 20371 6048
rect 24143 6042 24157 6096
rect 27286 6094 27292 6096
rect 27309 6110 27315 6111
rect 27593 6110 27607 6130
rect 27838 6128 27844 6130
rect 27861 6128 27867 6145
rect 27838 6125 27867 6128
rect 28205 6124 28208 6150
rect 28234 6144 28237 6150
rect 28344 6145 28373 6148
rect 28344 6144 28350 6145
rect 28234 6130 28350 6144
rect 28234 6124 28237 6130
rect 28344 6128 28350 6130
rect 28367 6128 28373 6145
rect 28344 6125 28373 6128
rect 37405 6124 37408 6150
rect 37434 6144 37437 6150
rect 38380 6148 38394 6164
rect 38601 6158 38604 6164
rect 38630 6158 38633 6184
rect 38740 6179 38769 6182
rect 38740 6162 38746 6179
rect 38763 6178 38769 6179
rect 39199 6178 39202 6184
rect 38763 6164 39202 6178
rect 38763 6162 38769 6164
rect 38740 6159 38769 6162
rect 39199 6158 39202 6164
rect 39228 6158 39231 6184
rect 38372 6145 38401 6148
rect 37434 6130 38348 6144
rect 37434 6124 37437 6130
rect 27309 6096 27607 6110
rect 27309 6094 27315 6096
rect 27286 6091 27315 6094
rect 27653 6090 27656 6116
rect 27682 6110 27685 6116
rect 28251 6110 28254 6116
rect 27682 6096 28254 6110
rect 27682 6090 27685 6096
rect 28251 6090 28254 6096
rect 28280 6110 28283 6116
rect 38334 6114 38348 6130
rect 38372 6128 38378 6145
rect 38395 6128 38401 6145
rect 38372 6125 38401 6128
rect 38463 6124 38466 6150
rect 38492 6144 38495 6150
rect 39061 6144 39064 6150
rect 38492 6130 39064 6144
rect 38492 6124 38495 6130
rect 39061 6124 39064 6130
rect 39090 6124 39093 6150
rect 28298 6111 28327 6114
rect 28298 6110 28304 6111
rect 28280 6096 28304 6110
rect 28280 6090 28283 6096
rect 28298 6094 28304 6096
rect 28321 6110 28327 6111
rect 28758 6111 28787 6114
rect 28758 6110 28764 6111
rect 28321 6096 28764 6110
rect 28321 6094 28327 6096
rect 28298 6091 28327 6094
rect 28758 6094 28764 6096
rect 28781 6094 28787 6111
rect 28758 6091 28787 6094
rect 29080 6111 29109 6114
rect 29080 6094 29086 6111
rect 29103 6094 29109 6111
rect 29080 6091 29109 6094
rect 37682 6111 37711 6114
rect 37682 6094 37688 6111
rect 37705 6110 37711 6111
rect 38326 6111 38355 6114
rect 37705 6096 38302 6110
rect 37705 6094 37711 6096
rect 37682 6091 37711 6094
rect 26319 6076 26322 6082
rect 26299 6062 26322 6076
rect 26319 6056 26322 6062
rect 26348 6056 26351 6082
rect 26549 6056 26552 6082
rect 26578 6056 26581 6082
rect 27746 6077 27775 6080
rect 26972 6062 27607 6076
rect 26972 6042 26986 6062
rect 24143 6028 26986 6042
rect 27593 6042 27607 6062
rect 27746 6060 27752 6077
rect 27769 6076 27775 6077
rect 29088 6076 29102 6091
rect 27769 6062 28044 6076
rect 27769 6060 27775 6062
rect 27746 6057 27775 6060
rect 28030 6048 28044 6062
rect 28076 6062 29102 6076
rect 38288 6076 38302 6096
rect 38326 6094 38332 6111
rect 38349 6110 38355 6111
rect 38969 6110 38972 6116
rect 38349 6096 38972 6110
rect 38349 6094 38355 6096
rect 38326 6091 38355 6094
rect 38969 6090 38972 6096
rect 38998 6090 39001 6116
rect 39254 6076 39268 6198
rect 39659 6192 39662 6198
rect 39688 6192 39691 6218
rect 40120 6213 40149 6216
rect 40120 6196 40126 6213
rect 40143 6212 40149 6213
rect 40257 6212 40260 6218
rect 40143 6198 40260 6212
rect 40143 6196 40149 6198
rect 40120 6193 40149 6196
rect 40257 6192 40260 6198
rect 40286 6192 40289 6218
rect 42741 6192 42744 6218
rect 42770 6212 42773 6218
rect 42788 6213 42817 6216
rect 42788 6212 42794 6213
rect 42770 6198 42794 6212
rect 42770 6192 42773 6198
rect 42788 6196 42794 6198
rect 42811 6196 42817 6213
rect 43201 6212 43204 6218
rect 43181 6198 43204 6212
rect 42788 6193 42817 6196
rect 43201 6192 43204 6198
rect 43230 6192 43233 6218
rect 43937 6192 43940 6218
rect 43966 6212 43969 6218
rect 44444 6213 44473 6216
rect 44444 6212 44450 6213
rect 43966 6198 44450 6212
rect 43966 6192 43969 6198
rect 44444 6196 44450 6198
rect 44467 6196 44473 6213
rect 45087 6212 45090 6218
rect 45067 6198 45090 6212
rect 44444 6193 44473 6196
rect 45087 6192 45090 6198
rect 45116 6192 45119 6218
rect 49550 6213 49579 6216
rect 49550 6196 49556 6213
rect 49573 6212 49579 6213
rect 49733 6212 49736 6218
rect 49573 6198 49736 6212
rect 49573 6196 49579 6198
rect 49550 6193 49579 6196
rect 49733 6192 49736 6198
rect 49762 6192 49765 6218
rect 49918 6213 49947 6216
rect 49918 6196 49924 6213
rect 49941 6212 49947 6213
rect 49963 6212 49966 6218
rect 49941 6198 49966 6212
rect 49941 6196 49947 6198
rect 49918 6193 49947 6196
rect 49963 6192 49966 6198
rect 49992 6192 49995 6218
rect 51942 6213 51971 6216
rect 51942 6196 51948 6213
rect 51965 6212 51971 6213
rect 52493 6212 52496 6218
rect 51965 6198 52496 6212
rect 51965 6196 51971 6198
rect 51942 6193 51971 6196
rect 52493 6192 52496 6198
rect 52522 6192 52525 6218
rect 52585 6212 52588 6218
rect 52565 6198 52588 6212
rect 52585 6192 52588 6198
rect 52614 6192 52617 6218
rect 56265 6192 56268 6218
rect 56294 6212 56297 6218
rect 56542 6213 56571 6216
rect 56542 6212 56548 6213
rect 56294 6198 56548 6212
rect 56294 6192 56297 6198
rect 56542 6196 56548 6198
rect 56565 6196 56571 6213
rect 56542 6193 56571 6196
rect 56864 6213 56893 6216
rect 56864 6196 56870 6213
rect 56887 6212 56893 6213
rect 57507 6212 57510 6218
rect 56887 6198 57510 6212
rect 56887 6196 56893 6198
rect 56864 6193 56893 6196
rect 57507 6192 57510 6198
rect 57536 6192 57539 6218
rect 58473 6192 58476 6218
rect 58502 6212 58505 6218
rect 59210 6213 59239 6216
rect 59210 6212 59216 6213
rect 58502 6198 59216 6212
rect 58502 6192 58505 6198
rect 59210 6196 59216 6198
rect 59233 6196 59239 6213
rect 59210 6193 59239 6196
rect 63856 6213 63885 6216
rect 63856 6196 63862 6213
rect 63879 6212 63885 6213
rect 63901 6212 63904 6218
rect 63879 6198 63904 6212
rect 63879 6196 63885 6198
rect 63856 6193 63885 6196
rect 63901 6192 63904 6198
rect 63930 6192 63933 6218
rect 64545 6192 64548 6218
rect 64574 6212 64577 6218
rect 65420 6213 65449 6216
rect 65420 6212 65426 6213
rect 64574 6198 65426 6212
rect 64574 6192 64577 6198
rect 65420 6196 65426 6198
rect 65443 6212 65449 6213
rect 65465 6212 65468 6218
rect 65443 6198 65468 6212
rect 65443 6196 65449 6198
rect 65420 6193 65449 6196
rect 65465 6192 65468 6198
rect 65494 6192 65497 6218
rect 66201 6192 66204 6218
rect 66230 6212 66233 6218
rect 66340 6213 66369 6216
rect 66340 6212 66346 6213
rect 66230 6198 66346 6212
rect 66230 6192 66233 6198
rect 66340 6196 66346 6198
rect 66363 6196 66369 6213
rect 66340 6193 66369 6196
rect 73654 6213 73683 6216
rect 73654 6196 73660 6213
rect 73677 6212 73683 6213
rect 73883 6212 73886 6218
rect 73677 6198 73886 6212
rect 73677 6196 73683 6198
rect 73654 6193 73683 6196
rect 73883 6192 73886 6198
rect 73912 6192 73915 6218
rect 76229 6192 76232 6218
rect 76258 6212 76261 6218
rect 76276 6213 76305 6216
rect 76276 6212 76282 6213
rect 76258 6198 76282 6212
rect 76258 6192 76261 6198
rect 76276 6196 76282 6198
rect 76299 6196 76305 6213
rect 76276 6193 76305 6196
rect 76422 6198 76712 6212
rect 43063 6178 43066 6184
rect 40082 6164 43066 6178
rect 39291 6090 39294 6116
rect 39320 6110 39323 6116
rect 40082 6114 40096 6164
rect 43063 6158 43066 6164
rect 43092 6158 43095 6184
rect 43707 6158 43710 6184
rect 43736 6178 43739 6184
rect 44720 6179 44749 6182
rect 44720 6178 44726 6179
rect 43736 6164 44726 6178
rect 43736 6158 43739 6164
rect 44720 6162 44726 6164
rect 44743 6162 44749 6179
rect 44720 6159 44749 6162
rect 47258 6164 56587 6178
rect 40717 6124 40720 6150
rect 40746 6144 40749 6150
rect 42236 6145 42265 6148
rect 42236 6144 42242 6145
rect 40746 6130 42242 6144
rect 40746 6124 40749 6130
rect 42236 6128 42242 6130
rect 42259 6128 42265 6145
rect 42327 6144 42330 6150
rect 42307 6130 42330 6144
rect 42236 6125 42265 6128
rect 42327 6124 42330 6130
rect 42356 6124 42359 6150
rect 42879 6144 42882 6150
rect 42520 6130 42882 6144
rect 39614 6111 39643 6114
rect 39614 6110 39620 6111
rect 39320 6096 39620 6110
rect 39320 6090 39323 6096
rect 39614 6094 39620 6096
rect 39637 6110 39643 6111
rect 40074 6111 40103 6114
rect 40074 6110 40080 6111
rect 39637 6096 40080 6110
rect 39637 6094 39643 6096
rect 39614 6091 39643 6094
rect 40074 6094 40080 6096
rect 40097 6094 40103 6111
rect 40074 6091 40103 6094
rect 41913 6090 41916 6116
rect 41942 6110 41945 6116
rect 42190 6111 42219 6114
rect 42190 6110 42196 6111
rect 41942 6096 42196 6110
rect 41942 6090 41945 6096
rect 42190 6094 42196 6096
rect 42213 6110 42219 6111
rect 42520 6110 42534 6130
rect 42879 6124 42882 6130
rect 42908 6124 42911 6150
rect 43155 6124 43158 6150
rect 43184 6144 43187 6150
rect 43524 6145 43553 6148
rect 43524 6144 43530 6145
rect 43184 6130 43530 6144
rect 43184 6124 43187 6130
rect 43524 6128 43530 6130
rect 43547 6144 43553 6145
rect 44075 6144 44078 6150
rect 43547 6130 44078 6144
rect 43547 6128 43553 6130
rect 43524 6125 43553 6128
rect 44075 6124 44078 6130
rect 44104 6124 44107 6150
rect 44581 6144 44584 6150
rect 44452 6130 44584 6144
rect 42741 6110 42744 6116
rect 42213 6096 42534 6110
rect 42721 6096 42744 6110
rect 42213 6094 42219 6096
rect 42190 6091 42219 6094
rect 42741 6090 42744 6096
rect 42770 6090 42773 6116
rect 43017 6090 43020 6116
rect 43046 6110 43049 6116
rect 43432 6111 43461 6114
rect 43432 6110 43438 6111
rect 43046 6096 43438 6110
rect 43046 6090 43049 6096
rect 43432 6094 43438 6096
rect 43455 6094 43461 6111
rect 43432 6091 43461 6094
rect 43984 6111 44013 6114
rect 43984 6094 43990 6111
rect 44007 6110 44013 6111
rect 44121 6110 44124 6116
rect 44007 6096 44124 6110
rect 44007 6094 44013 6096
rect 43984 6091 44013 6094
rect 44121 6090 44124 6096
rect 44150 6090 44153 6116
rect 44398 6111 44427 6114
rect 44398 6094 44404 6111
rect 44421 6111 44427 6111
rect 44452 6111 44466 6130
rect 44581 6124 44584 6130
rect 44610 6144 44613 6150
rect 44610 6130 45064 6144
rect 44610 6124 44613 6130
rect 44421 6097 44466 6111
rect 44421 6094 44427 6097
rect 44398 6091 44427 6094
rect 44489 6090 44492 6116
rect 44518 6110 44521 6116
rect 45050 6114 45064 6130
rect 44812 6111 44841 6114
rect 44812 6110 44818 6111
rect 44518 6096 44818 6110
rect 44518 6090 44521 6096
rect 44812 6094 44818 6096
rect 44835 6094 44841 6111
rect 44812 6091 44841 6094
rect 45042 6111 45071 6114
rect 45042 6094 45048 6111
rect 45065 6110 45071 6111
rect 46007 6110 46010 6116
rect 45065 6096 46010 6110
rect 45065 6094 45071 6096
rect 45042 6091 45071 6094
rect 46007 6090 46010 6096
rect 46036 6090 46039 6116
rect 47258 6076 47272 6164
rect 49549 6124 49552 6150
rect 49578 6144 49581 6150
rect 50470 6145 50499 6148
rect 50470 6144 50476 6145
rect 49578 6130 50476 6144
rect 49578 6124 49581 6130
rect 50470 6128 50476 6130
rect 50493 6144 50499 6145
rect 51021 6144 51024 6150
rect 50493 6130 51024 6144
rect 50493 6128 50499 6130
rect 50470 6125 50499 6128
rect 51021 6124 51024 6130
rect 51050 6144 51053 6150
rect 51574 6145 51603 6148
rect 51574 6144 51580 6145
rect 51050 6130 51580 6144
rect 51050 6124 51053 6130
rect 51574 6128 51580 6130
rect 51597 6144 51603 6145
rect 51619 6144 51622 6150
rect 51597 6130 51622 6144
rect 51597 6128 51603 6130
rect 51574 6125 51603 6128
rect 51619 6124 51622 6130
rect 51648 6124 51651 6150
rect 51665 6124 51668 6150
rect 51694 6144 51697 6150
rect 52264 6145 52293 6148
rect 52264 6144 52270 6145
rect 51694 6130 52270 6144
rect 51694 6124 51697 6130
rect 52264 6128 52270 6130
rect 52287 6128 52293 6145
rect 56573 6144 56587 6164
rect 57875 6158 57878 6184
rect 57904 6178 57907 6184
rect 70985 6178 70988 6184
rect 57904 6164 58910 6178
rect 57904 6158 57907 6164
rect 58896 6148 58910 6164
rect 65198 6164 70988 6178
rect 57186 6145 57215 6148
rect 57186 6144 57192 6145
rect 56573 6130 57192 6144
rect 52264 6125 52293 6128
rect 57186 6128 57192 6130
rect 57209 6144 57215 6145
rect 58888 6145 58917 6148
rect 57209 6130 58404 6144
rect 57209 6128 57215 6130
rect 57186 6125 57215 6128
rect 48767 6090 48770 6116
rect 48796 6110 48799 6116
rect 49642 6111 49671 6114
rect 49642 6110 49648 6111
rect 48796 6096 49648 6110
rect 48796 6090 48799 6096
rect 49642 6094 49648 6096
rect 49665 6094 49671 6111
rect 49642 6091 49671 6094
rect 49872 6111 49901 6114
rect 49872 6094 49878 6111
rect 49895 6110 49901 6111
rect 51482 6111 51511 6114
rect 49895 6096 51090 6110
rect 49895 6094 49901 6096
rect 49872 6091 49901 6094
rect 51076 6082 51090 6096
rect 51482 6094 51488 6111
rect 51505 6110 51511 6111
rect 51849 6110 51852 6116
rect 51505 6096 51852 6110
rect 51505 6094 51511 6096
rect 51482 6091 51511 6094
rect 51849 6090 51852 6096
rect 51878 6090 51881 6116
rect 51896 6111 51925 6114
rect 51896 6094 51902 6111
rect 51919 6110 51925 6111
rect 52218 6111 52247 6114
rect 52218 6110 52224 6111
rect 51919 6096 52224 6110
rect 51919 6094 51925 6096
rect 51896 6091 51925 6094
rect 52218 6094 52224 6096
rect 52241 6110 52247 6111
rect 52540 6111 52569 6114
rect 52540 6110 52546 6111
rect 52241 6096 52546 6110
rect 52241 6094 52247 6096
rect 52218 6091 52247 6094
rect 52540 6094 52546 6096
rect 52563 6094 52569 6111
rect 52540 6091 52569 6094
rect 50377 6076 50380 6082
rect 38288 6062 38946 6076
rect 39254 6062 44420 6076
rect 27929 6042 27932 6048
rect 27593 6028 27932 6042
rect 27929 6022 27932 6028
rect 27958 6022 27961 6048
rect 28021 6042 28024 6048
rect 28001 6028 28024 6042
rect 28021 6022 28024 6028
rect 28050 6022 28053 6048
rect 28076 6046 28090 6062
rect 28068 6043 28097 6046
rect 28068 6026 28074 6043
rect 28091 6026 28097 6043
rect 28068 6023 28097 6026
rect 28252 6043 28281 6046
rect 28252 6026 28258 6043
rect 28275 6042 28281 6043
rect 28665 6042 28668 6048
rect 28275 6028 28668 6042
rect 28275 6026 28281 6028
rect 28252 6023 28281 6026
rect 28665 6022 28668 6028
rect 28694 6022 28697 6048
rect 38141 6042 38144 6048
rect 38121 6028 38144 6042
rect 38141 6022 38144 6028
rect 38170 6022 38173 6048
rect 38932 6046 38946 6062
rect 38924 6043 38953 6046
rect 38924 6026 38930 6043
rect 38947 6042 38953 6043
rect 40119 6042 40122 6048
rect 38947 6028 40122 6042
rect 38947 6026 38953 6028
rect 38924 6023 38953 6026
rect 40119 6022 40122 6028
rect 40148 6022 40151 6048
rect 42005 6042 42008 6048
rect 41985 6028 42008 6042
rect 42005 6022 42008 6028
rect 42034 6022 42037 6048
rect 42327 6022 42330 6048
rect 42356 6042 42359 6048
rect 43155 6042 43158 6048
rect 42356 6028 43158 6042
rect 42356 6022 42359 6028
rect 43155 6022 43158 6028
rect 43184 6022 43187 6048
rect 43386 6043 43415 6046
rect 43386 6026 43392 6043
rect 43409 6042 43415 6043
rect 43753 6042 43756 6048
rect 43409 6028 43756 6042
rect 43409 6026 43415 6028
rect 43386 6023 43415 6026
rect 43753 6022 43756 6028
rect 43782 6022 43785 6048
rect 43800 6043 43829 6046
rect 43800 6026 43806 6043
rect 43823 6042 43829 6043
rect 43891 6042 43894 6048
rect 43823 6028 43894 6042
rect 43823 6026 43829 6028
rect 43800 6023 43829 6026
rect 43891 6022 43894 6028
rect 43920 6022 43923 6048
rect 43983 6022 43986 6048
rect 44012 6042 44015 6048
rect 44030 6043 44059 6046
rect 44030 6042 44036 6043
rect 44012 6028 44036 6042
rect 44012 6022 44015 6028
rect 44030 6026 44036 6028
rect 44053 6042 44059 6043
rect 44351 6042 44354 6048
rect 44053 6028 44354 6042
rect 44053 6026 44059 6028
rect 44030 6023 44059 6026
rect 44351 6022 44354 6028
rect 44380 6022 44383 6048
rect 44406 6042 44420 6062
rect 44843 6062 47272 6076
rect 50357 6062 50380 6076
rect 44843 6042 44857 6062
rect 50377 6056 50380 6062
rect 50406 6056 50409 6082
rect 50424 6077 50453 6080
rect 50424 6060 50430 6077
rect 50447 6076 50453 6077
rect 50515 6076 50518 6082
rect 50447 6062 50518 6076
rect 50447 6060 50453 6062
rect 50424 6057 50453 6060
rect 50515 6056 50518 6062
rect 50544 6056 50547 6082
rect 50975 6076 50978 6082
rect 50955 6062 50978 6076
rect 50975 6056 50978 6062
rect 51004 6056 51007 6082
rect 51067 6056 51070 6082
rect 51096 6076 51099 6082
rect 51904 6076 51918 6091
rect 55943 6090 55946 6116
rect 55972 6110 55975 6116
rect 56634 6111 56663 6114
rect 56634 6110 56640 6111
rect 55972 6096 56640 6110
rect 55972 6090 55975 6096
rect 56634 6094 56640 6096
rect 56657 6094 56663 6111
rect 56634 6091 56663 6094
rect 56956 6111 56985 6114
rect 56956 6094 56962 6111
rect 56979 6110 56985 6111
rect 57139 6110 57142 6116
rect 56979 6096 57142 6110
rect 56979 6094 56985 6096
rect 56956 6091 56985 6094
rect 57139 6090 57142 6096
rect 57168 6090 57171 6116
rect 58390 6110 58404 6130
rect 58888 6128 58894 6145
rect 58911 6144 58917 6145
rect 59439 6144 59442 6150
rect 58911 6130 59442 6144
rect 58911 6128 58917 6130
rect 58888 6125 58917 6128
rect 59439 6124 59442 6130
rect 59468 6124 59471 6150
rect 65198 6144 65212 6164
rect 70985 6158 70988 6164
rect 71014 6158 71017 6184
rect 73791 6158 73794 6184
rect 73820 6178 73823 6184
rect 74206 6179 74235 6182
rect 74206 6178 74212 6179
rect 73820 6164 74212 6178
rect 73820 6158 73823 6164
rect 74206 6162 74212 6164
rect 74229 6162 74235 6179
rect 74206 6159 74235 6162
rect 75815 6158 75818 6184
rect 75844 6178 75847 6184
rect 76367 6178 76370 6184
rect 75844 6164 76370 6178
rect 75844 6158 75847 6164
rect 64554 6130 65212 6144
rect 58796 6111 58825 6114
rect 58390 6096 58634 6110
rect 51096 6062 51918 6076
rect 51096 6056 51099 6062
rect 56909 6056 56912 6082
rect 56938 6076 56941 6082
rect 57324 6077 57353 6080
rect 57324 6076 57330 6077
rect 56938 6062 57330 6076
rect 56938 6056 56941 6062
rect 57324 6060 57330 6062
rect 57347 6060 57353 6077
rect 57324 6057 57353 6060
rect 57378 6062 57569 6076
rect 50193 6042 50196 6048
rect 44406 6028 44857 6042
rect 50173 6028 50196 6042
rect 50193 6022 50196 6028
rect 50222 6022 50225 6048
rect 50984 6042 50998 6056
rect 51159 6042 51162 6048
rect 50984 6028 51162 6042
rect 51159 6022 51162 6028
rect 51188 6022 51191 6048
rect 51297 6042 51300 6048
rect 51277 6028 51300 6042
rect 51297 6022 51300 6028
rect 51326 6022 51329 6048
rect 51527 6042 51530 6048
rect 51507 6028 51530 6042
rect 51527 6022 51530 6028
rect 51556 6022 51559 6048
rect 56955 6022 56958 6048
rect 56984 6042 56987 6048
rect 57378 6042 57392 6062
rect 56984 6028 57392 6042
rect 56984 6022 56987 6028
rect 57829 6022 57832 6048
rect 57858 6042 57861 6048
rect 58060 6043 58089 6046
rect 58060 6042 58066 6043
rect 57858 6028 58066 6042
rect 57858 6022 57861 6028
rect 58060 6026 58066 6028
rect 58083 6026 58089 6043
rect 58060 6023 58089 6026
rect 58197 6022 58200 6048
rect 58226 6042 58229 6048
rect 58566 6043 58595 6046
rect 58566 6042 58572 6043
rect 58226 6028 58572 6042
rect 58226 6022 58229 6028
rect 58566 6026 58572 6028
rect 58589 6026 58595 6043
rect 58620 6042 58634 6096
rect 58796 6094 58802 6111
rect 58819 6110 58825 6111
rect 59025 6110 59028 6116
rect 58819 6096 59028 6110
rect 58819 6094 58825 6096
rect 58796 6091 58825 6094
rect 59025 6090 59028 6096
rect 59054 6090 59057 6116
rect 59163 6110 59166 6116
rect 59143 6096 59166 6110
rect 59163 6090 59166 6096
rect 59192 6090 59195 6116
rect 63073 6090 63076 6116
rect 63102 6110 63105 6116
rect 63948 6111 63977 6114
rect 63948 6110 63954 6111
rect 63102 6096 63954 6110
rect 63102 6090 63105 6096
rect 63948 6094 63954 6096
rect 63971 6094 63977 6111
rect 64315 6110 64318 6116
rect 64295 6096 64318 6110
rect 63948 6091 63977 6094
rect 64315 6090 64318 6096
rect 64344 6090 64347 6116
rect 64554 6114 64568 6130
rect 65511 6124 65514 6150
rect 65540 6144 65543 6150
rect 65926 6145 65955 6148
rect 65926 6144 65932 6145
rect 65540 6130 65932 6144
rect 65540 6124 65543 6130
rect 65926 6128 65932 6130
rect 65949 6144 65955 6145
rect 66615 6144 66618 6150
rect 65949 6130 66618 6144
rect 65949 6128 65955 6130
rect 65926 6125 65955 6128
rect 66615 6124 66618 6130
rect 66644 6124 66647 6150
rect 74527 6124 74530 6150
rect 74556 6144 74559 6150
rect 76046 6145 76075 6148
rect 76046 6144 76052 6145
rect 74556 6130 76052 6144
rect 74556 6124 74559 6130
rect 76046 6128 76052 6130
rect 76069 6128 76075 6145
rect 76046 6125 76075 6128
rect 76092 6145 76121 6148
rect 76092 6128 76098 6145
rect 76115 6128 76121 6145
rect 76092 6125 76121 6128
rect 64546 6111 64575 6114
rect 64546 6094 64552 6111
rect 64569 6094 64575 6111
rect 64546 6091 64575 6094
rect 58750 6077 58779 6080
rect 58750 6060 58756 6077
rect 58773 6076 58779 6077
rect 59117 6076 59120 6082
rect 58773 6062 59120 6076
rect 58773 6060 58779 6062
rect 58750 6057 58779 6060
rect 59117 6056 59120 6062
rect 59146 6056 59149 6082
rect 64554 6076 64568 6091
rect 65235 6090 65238 6116
rect 65264 6090 65267 6116
rect 65834 6111 65863 6114
rect 65834 6094 65840 6111
rect 65857 6110 65863 6111
rect 66201 6110 66204 6116
rect 65857 6096 66204 6110
rect 65857 6094 65863 6096
rect 65834 6091 65863 6094
rect 66201 6090 66204 6096
rect 66230 6090 66233 6116
rect 66293 6110 66296 6116
rect 66273 6096 66296 6110
rect 66293 6090 66296 6096
rect 66322 6090 66325 6116
rect 68869 6110 68872 6116
rect 68849 6096 68872 6110
rect 68869 6090 68872 6096
rect 68898 6090 68901 6116
rect 73746 6111 73775 6114
rect 73746 6094 73752 6111
rect 73769 6110 73775 6111
rect 74021 6110 74024 6116
rect 73769 6096 74024 6110
rect 73769 6094 73775 6096
rect 73746 6091 73775 6094
rect 74021 6090 74024 6096
rect 74050 6090 74053 6116
rect 74160 6111 74189 6114
rect 74160 6094 74166 6111
rect 74183 6110 74189 6111
rect 74665 6110 74668 6116
rect 74183 6096 74668 6110
rect 74183 6094 74189 6096
rect 74160 6091 74189 6094
rect 74665 6090 74668 6096
rect 74694 6090 74697 6116
rect 74711 6090 74714 6116
rect 74740 6110 74743 6116
rect 74740 6096 74762 6110
rect 74740 6090 74743 6096
rect 75677 6090 75680 6116
rect 75706 6110 75709 6116
rect 76100 6110 76114 6125
rect 76238 6114 76252 6164
rect 76367 6158 76370 6164
rect 76396 6158 76399 6184
rect 75706 6096 76114 6110
rect 76230 6111 76259 6114
rect 75706 6090 75709 6096
rect 76230 6094 76236 6111
rect 76253 6094 76259 6111
rect 76230 6091 76259 6094
rect 61403 6062 64568 6076
rect 64684 6077 64713 6080
rect 61403 6042 61417 6062
rect 64684 6060 64690 6077
rect 64707 6060 64713 6077
rect 66247 6076 66250 6082
rect 64684 6057 64713 6060
rect 65658 6062 66250 6076
rect 58620 6028 61417 6042
rect 64224 6043 64253 6046
rect 58566 6023 58595 6026
rect 64224 6026 64230 6043
rect 64247 6042 64253 6043
rect 64692 6042 64706 6057
rect 65658 6046 65672 6062
rect 66247 6056 66250 6062
rect 66276 6056 66279 6082
rect 69007 6076 69010 6082
rect 68987 6062 69010 6076
rect 69007 6056 69010 6062
rect 69036 6076 69039 6082
rect 72918 6077 72947 6080
rect 72918 6076 72924 6077
rect 69036 6062 72924 6076
rect 69036 6056 69039 6062
rect 72918 6060 72924 6062
rect 72941 6060 72947 6077
rect 72918 6057 72947 6060
rect 73102 6077 73131 6080
rect 73102 6060 73108 6077
rect 73125 6076 73131 6077
rect 76422 6076 76436 6198
rect 76644 6179 76673 6182
rect 76644 6162 76650 6179
rect 76667 6162 76673 6179
rect 76698 6178 76712 6198
rect 76873 6192 76876 6218
rect 76902 6212 76905 6218
rect 77058 6213 77087 6216
rect 77058 6212 77064 6213
rect 76902 6198 77064 6212
rect 76902 6192 76905 6198
rect 77058 6196 77064 6198
rect 77081 6196 77087 6213
rect 77058 6193 77087 6196
rect 78621 6192 78624 6218
rect 78650 6212 78653 6218
rect 80461 6212 80464 6218
rect 78650 6198 80464 6212
rect 78650 6192 78653 6198
rect 80461 6192 80464 6198
rect 80490 6192 80493 6218
rect 80783 6192 80786 6218
rect 80812 6212 80815 6218
rect 82670 6213 82699 6216
rect 80812 6198 82462 6212
rect 80812 6192 80815 6198
rect 77517 6178 77520 6184
rect 76698 6164 77520 6178
rect 76644 6159 76673 6162
rect 76652 6110 76666 6159
rect 77517 6158 77520 6164
rect 77546 6158 77549 6184
rect 79449 6158 79452 6184
rect 79478 6178 79481 6184
rect 80002 6179 80031 6182
rect 80002 6178 80008 6179
rect 79478 6164 80008 6178
rect 79478 6158 79481 6164
rect 80002 6162 80008 6164
rect 80025 6162 80031 6179
rect 82448 6178 82462 6198
rect 82670 6196 82676 6213
rect 82693 6212 82699 6213
rect 83221 6212 83224 6218
rect 82693 6198 83224 6212
rect 82693 6196 82699 6198
rect 82670 6193 82699 6196
rect 83221 6192 83224 6198
rect 83250 6192 83253 6218
rect 87960 6213 87989 6216
rect 87960 6196 87966 6213
rect 87983 6212 87989 6213
rect 88235 6212 88238 6218
rect 87983 6198 88238 6212
rect 87983 6196 87989 6198
rect 87960 6193 87989 6196
rect 88235 6192 88238 6198
rect 88264 6192 88267 6218
rect 89753 6192 89756 6218
rect 89782 6212 89785 6218
rect 90674 6213 90703 6216
rect 90674 6212 90680 6213
rect 89782 6198 90680 6212
rect 89782 6192 89785 6198
rect 90674 6196 90680 6198
rect 90697 6196 90703 6213
rect 90674 6193 90703 6196
rect 94262 6213 94291 6216
rect 94262 6196 94268 6213
rect 94285 6212 94291 6213
rect 94583 6212 94586 6218
rect 94285 6198 94586 6212
rect 94285 6196 94291 6198
rect 94262 6193 94291 6196
rect 94583 6192 94586 6198
rect 94612 6192 94615 6218
rect 94813 6192 94816 6218
rect 94842 6212 94845 6218
rect 95090 6213 95119 6216
rect 95090 6212 95096 6213
rect 94842 6198 95096 6212
rect 94842 6192 94845 6198
rect 95090 6196 95096 6198
rect 95113 6196 95119 6213
rect 95090 6193 95119 6196
rect 95411 6192 95414 6218
rect 95440 6212 95443 6218
rect 97021 6212 97024 6218
rect 95440 6198 97024 6212
rect 95440 6192 95443 6198
rect 97021 6192 97024 6198
rect 97050 6192 97053 6218
rect 100840 6213 100869 6216
rect 97076 6198 98792 6212
rect 82715 6178 82718 6184
rect 82448 6164 82718 6178
rect 80002 6159 80031 6162
rect 82715 6158 82718 6164
rect 82744 6158 82747 6184
rect 83037 6178 83040 6184
rect 83017 6164 83040 6178
rect 83037 6158 83040 6164
rect 83066 6158 83069 6184
rect 88879 6178 88882 6184
rect 88520 6164 88882 6178
rect 76966 6145 76995 6148
rect 76966 6128 76972 6145
rect 76989 6144 76995 6145
rect 77057 6144 77060 6150
rect 76989 6130 77060 6144
rect 76989 6128 76995 6130
rect 76966 6125 76995 6128
rect 77057 6124 77060 6130
rect 77086 6124 77089 6150
rect 80185 6124 80188 6150
rect 80214 6144 80217 6150
rect 80646 6145 80675 6148
rect 80646 6144 80652 6145
rect 80214 6130 80652 6144
rect 80214 6124 80217 6130
rect 80646 6128 80652 6130
rect 80669 6128 80675 6145
rect 80646 6125 80675 6128
rect 80737 6124 80740 6150
rect 80766 6144 80769 6150
rect 81243 6144 81246 6150
rect 80766 6130 80788 6144
rect 81223 6130 81246 6144
rect 80766 6124 80769 6130
rect 81243 6124 81246 6130
rect 81272 6124 81275 6150
rect 81335 6144 81338 6150
rect 81315 6130 81338 6144
rect 81335 6124 81338 6130
rect 81364 6124 81367 6150
rect 81795 6144 81798 6150
rect 81775 6130 81798 6144
rect 81795 6124 81798 6130
rect 81824 6124 81827 6150
rect 88520 6148 88534 6164
rect 88879 6158 88882 6164
rect 88908 6158 88911 6184
rect 90443 6178 90446 6184
rect 90423 6164 90446 6178
rect 90443 6158 90446 6164
rect 90472 6158 90475 6184
rect 96285 6178 96288 6184
rect 92798 6164 95250 6178
rect 96265 6164 96288 6178
rect 88512 6145 88541 6148
rect 88512 6128 88518 6145
rect 88535 6128 88541 6145
rect 88512 6125 88541 6128
rect 88557 6124 88560 6150
rect 88586 6144 88589 6150
rect 92798 6144 92812 6164
rect 88586 6130 88608 6144
rect 89578 6130 92812 6144
rect 88586 6124 88589 6130
rect 77150 6111 77179 6114
rect 77150 6110 77156 6111
rect 76652 6096 77156 6110
rect 77150 6094 77156 6096
rect 77173 6094 77179 6111
rect 77150 6091 77179 6094
rect 79403 6090 79406 6116
rect 79432 6110 79435 6116
rect 80094 6111 80123 6114
rect 80094 6110 80100 6111
rect 79432 6096 80100 6110
rect 79432 6090 79435 6096
rect 80094 6094 80100 6096
rect 80117 6094 80123 6111
rect 80094 6091 80123 6094
rect 80600 6111 80629 6114
rect 80600 6094 80606 6111
rect 80623 6110 80629 6111
rect 80875 6110 80878 6116
rect 80623 6096 80878 6110
rect 80623 6094 80629 6096
rect 80600 6091 80629 6094
rect 80875 6090 80878 6096
rect 80904 6110 80907 6116
rect 81252 6110 81266 6124
rect 89578 6116 89592 6130
rect 93985 6124 93988 6150
rect 94014 6144 94017 6150
rect 94014 6130 95204 6144
rect 94014 6124 94017 6130
rect 80904 6096 81266 6110
rect 88052 6111 88081 6114
rect 80904 6090 80907 6096
rect 88052 6094 88058 6111
rect 88075 6110 88081 6111
rect 88466 6111 88495 6114
rect 88466 6110 88472 6111
rect 88075 6096 88472 6110
rect 88075 6094 88081 6096
rect 88052 6091 88081 6094
rect 88466 6094 88472 6096
rect 88489 6110 88495 6111
rect 88925 6110 88928 6116
rect 88489 6096 88928 6110
rect 88489 6094 88495 6096
rect 88466 6091 88495 6094
rect 88925 6090 88928 6096
rect 88954 6090 88957 6116
rect 89569 6110 89572 6116
rect 89549 6096 89572 6110
rect 89569 6090 89572 6096
rect 89598 6090 89601 6116
rect 90351 6090 90354 6116
rect 90380 6110 90383 6116
rect 90766 6111 90795 6114
rect 90766 6110 90772 6111
rect 90380 6096 90772 6110
rect 90380 6090 90383 6096
rect 90766 6094 90772 6096
rect 90789 6094 90795 6111
rect 90766 6091 90795 6094
rect 94354 6111 94383 6114
rect 94354 6094 94360 6111
rect 94377 6094 94383 6111
rect 94767 6110 94770 6116
rect 94747 6096 94770 6110
rect 94354 6091 94383 6094
rect 73125 6062 73837 6076
rect 73125 6060 73131 6062
rect 73102 6057 73131 6060
rect 64247 6028 64706 6042
rect 65650 6043 65679 6046
rect 64247 6026 64253 6028
rect 64224 6023 64253 6026
rect 65650 6026 65656 6043
rect 65673 6026 65679 6043
rect 65650 6023 65679 6026
rect 65787 6022 65790 6048
rect 65816 6042 65819 6048
rect 65880 6043 65909 6046
rect 65880 6042 65886 6043
rect 65816 6028 65886 6042
rect 65816 6022 65819 6028
rect 65880 6026 65886 6028
rect 65903 6026 65909 6043
rect 73823 6042 73837 6062
rect 74720 6062 76436 6076
rect 76828 6077 76857 6080
rect 74720 6042 74734 6062
rect 76828 6060 76834 6077
rect 76851 6076 76857 6077
rect 77931 6076 77934 6082
rect 76851 6062 77934 6076
rect 76851 6060 76857 6062
rect 76828 6057 76857 6060
rect 77931 6056 77934 6062
rect 77960 6056 77963 6082
rect 78207 6056 78210 6082
rect 78236 6076 78239 6082
rect 81289 6076 81292 6082
rect 78236 6062 81292 6076
rect 78236 6056 78239 6062
rect 81289 6056 81292 6062
rect 81318 6056 81321 6082
rect 81335 6056 81338 6082
rect 81364 6076 81367 6082
rect 81934 6077 81963 6080
rect 81934 6076 81940 6077
rect 81364 6062 81940 6076
rect 81364 6056 81367 6062
rect 81934 6060 81940 6062
rect 81957 6060 81963 6077
rect 81934 6057 81963 6060
rect 82163 6056 82166 6082
rect 82192 6056 82195 6082
rect 82945 6076 82948 6082
rect 82925 6062 82948 6076
rect 82945 6056 82948 6062
rect 82974 6056 82977 6082
rect 83267 6056 83270 6082
rect 83296 6076 83299 6082
rect 88972 6077 89001 6080
rect 88972 6076 88978 6077
rect 83296 6062 88978 6076
rect 83296 6056 83299 6062
rect 88972 6060 88978 6062
rect 88995 6076 89001 6077
rect 89707 6076 89710 6082
rect 88995 6062 89638 6076
rect 89687 6062 89710 6076
rect 88995 6060 89001 6062
rect 88972 6057 89001 6060
rect 73823 6028 74734 6042
rect 65880 6023 65909 6026
rect 74757 6022 74760 6048
rect 74786 6042 74789 6048
rect 75356 6043 75385 6046
rect 75356 6042 75362 6043
rect 74786 6028 75362 6042
rect 74786 6022 74789 6028
rect 75356 6026 75362 6028
rect 75379 6026 75385 6043
rect 75815 6042 75818 6048
rect 75795 6028 75818 6042
rect 75356 6023 75385 6026
rect 75815 6022 75818 6028
rect 75844 6022 75847 6048
rect 75861 6022 75864 6048
rect 75890 6042 75893 6048
rect 76000 6043 76029 6046
rect 76000 6042 76006 6043
rect 75890 6028 76006 6042
rect 75890 6022 75893 6028
rect 76000 6026 76006 6028
rect 76023 6026 76029 6043
rect 76000 6023 76029 6026
rect 76091 6022 76094 6048
rect 76120 6042 76123 6048
rect 76275 6042 76278 6048
rect 76120 6028 76278 6042
rect 76120 6022 76123 6028
rect 76275 6022 76278 6028
rect 76304 6042 76307 6048
rect 76874 6043 76903 6046
rect 76874 6042 76880 6043
rect 76304 6028 76880 6042
rect 76304 6022 76307 6028
rect 76874 6026 76880 6028
rect 76897 6026 76903 6043
rect 76874 6023 76903 6026
rect 80416 6043 80445 6046
rect 80416 6026 80422 6043
rect 80439 6042 80445 6043
rect 80553 6042 80556 6048
rect 80439 6028 80556 6042
rect 80439 6026 80445 6028
rect 80416 6023 80445 6026
rect 80553 6022 80556 6028
rect 80582 6022 80585 6048
rect 81014 6043 81043 6046
rect 81014 6026 81020 6043
rect 81037 6042 81043 6043
rect 81105 6042 81108 6048
rect 81037 6028 81108 6042
rect 81037 6026 81043 6028
rect 81014 6023 81043 6026
rect 81105 6022 81108 6028
rect 81134 6022 81137 6048
rect 81198 6043 81227 6046
rect 81198 6026 81204 6043
rect 81221 6042 81227 6043
rect 81427 6042 81430 6048
rect 81221 6028 81430 6042
rect 81221 6026 81227 6028
rect 81198 6023 81227 6026
rect 81427 6022 81430 6028
rect 81456 6022 81459 6048
rect 88282 6043 88311 6046
rect 88282 6026 88288 6043
rect 88305 6042 88311 6043
rect 88327 6042 88330 6048
rect 88305 6028 88330 6042
rect 88305 6026 88311 6028
rect 88282 6023 88311 6026
rect 88327 6022 88330 6028
rect 88356 6022 88359 6048
rect 89017 6042 89020 6048
rect 88997 6028 89020 6042
rect 89017 6022 89020 6028
rect 89046 6022 89049 6048
rect 89624 6042 89638 6062
rect 89707 6056 89710 6062
rect 89736 6056 89739 6082
rect 90719 6076 90722 6082
rect 90321 6062 90722 6076
rect 90719 6056 90722 6062
rect 90748 6056 90751 6082
rect 94362 6076 94376 6091
rect 94767 6090 94770 6096
rect 94796 6090 94799 6116
rect 95190 6114 95204 6130
rect 95182 6111 95211 6114
rect 95182 6094 95188 6111
rect 95205 6094 95211 6111
rect 95236 6110 95250 6164
rect 96285 6158 96288 6164
rect 96314 6158 96317 6184
rect 95412 6145 95441 6148
rect 95412 6128 95418 6145
rect 95435 6144 95441 6145
rect 95917 6144 95920 6150
rect 95435 6130 95920 6144
rect 95435 6128 95441 6130
rect 95412 6125 95441 6128
rect 95420 6110 95434 6125
rect 95917 6124 95920 6130
rect 95946 6124 95949 6150
rect 96331 6124 96334 6150
rect 96360 6144 96363 6150
rect 96838 6145 96867 6148
rect 96838 6144 96844 6145
rect 96360 6130 96844 6144
rect 96360 6124 96363 6130
rect 96838 6128 96844 6130
rect 96861 6144 96867 6145
rect 97076 6144 97090 6198
rect 98723 6178 98726 6184
rect 98226 6164 98726 6178
rect 96861 6130 97090 6144
rect 97214 6130 98010 6144
rect 96861 6128 96867 6130
rect 96838 6125 96867 6128
rect 97214 6116 97228 6130
rect 97205 6110 97208 6116
rect 95236 6096 95434 6110
rect 96202 6096 96906 6110
rect 97185 6096 97208 6110
rect 95182 6091 95211 6094
rect 95411 6076 95414 6082
rect 94362 6062 95414 6076
rect 95411 6056 95414 6062
rect 95440 6056 95443 6082
rect 95549 6076 95552 6082
rect 95529 6062 95552 6076
rect 95549 6056 95552 6062
rect 95578 6056 95581 6082
rect 95595 6056 95598 6082
rect 95624 6076 95627 6082
rect 95624 6062 95795 6076
rect 95624 6056 95627 6062
rect 90075 6042 90078 6048
rect 89624 6028 90078 6042
rect 90075 6022 90078 6028
rect 90104 6022 90107 6048
rect 94814 6043 94843 6046
rect 94814 6026 94820 6043
rect 94837 6042 94843 6043
rect 96202 6042 96216 6096
rect 96699 6076 96702 6082
rect 96679 6062 96702 6076
rect 96699 6056 96702 6062
rect 96728 6056 96731 6082
rect 96515 6042 96518 6048
rect 94837 6028 96216 6042
rect 96495 6028 96518 6042
rect 94837 6026 94843 6028
rect 94814 6023 94843 6026
rect 96515 6022 96518 6028
rect 96544 6022 96547 6048
rect 96746 6043 96775 6046
rect 96746 6026 96752 6043
rect 96769 6042 96775 6043
rect 96837 6042 96840 6048
rect 96769 6028 96840 6042
rect 96769 6026 96775 6028
rect 96746 6023 96775 6026
rect 96837 6022 96840 6028
rect 96866 6022 96869 6048
rect 96892 6042 96906 6096
rect 97205 6090 97208 6096
rect 97234 6090 97237 6116
rect 97343 6076 97346 6082
rect 97323 6062 97346 6076
rect 97343 6056 97346 6062
rect 97372 6056 97375 6082
rect 97996 6076 98010 6130
rect 98226 6114 98240 6164
rect 98723 6158 98726 6164
rect 98752 6158 98755 6184
rect 98778 6148 98792 6198
rect 100840 6196 100846 6213
rect 100863 6212 100869 6213
rect 101207 6212 101210 6218
rect 100863 6198 101210 6212
rect 100863 6196 100869 6198
rect 100840 6193 100869 6196
rect 101207 6192 101210 6198
rect 101236 6192 101239 6218
rect 102817 6212 102820 6218
rect 101814 6198 102820 6212
rect 100564 6179 100593 6182
rect 100564 6162 100570 6179
rect 100587 6178 100593 6179
rect 101814 6178 101828 6198
rect 102817 6192 102820 6198
rect 102846 6192 102849 6218
rect 103232 6213 103261 6216
rect 103232 6196 103238 6213
rect 103255 6212 103261 6213
rect 103829 6212 103832 6218
rect 103255 6198 103832 6212
rect 103255 6196 103261 6198
rect 103232 6193 103261 6196
rect 103829 6192 103832 6198
rect 103858 6192 103861 6218
rect 113898 6213 113927 6216
rect 113898 6196 113904 6213
rect 113921 6212 113927 6213
rect 115053 6212 115056 6218
rect 113921 6198 115056 6212
rect 113921 6196 113927 6198
rect 113898 6193 113927 6196
rect 115053 6192 115056 6198
rect 115082 6192 115085 6218
rect 115927 6192 115930 6218
rect 115956 6212 115959 6218
rect 116112 6213 116141 6216
rect 116112 6212 116118 6213
rect 115956 6198 116118 6212
rect 115956 6192 115959 6198
rect 116112 6196 116118 6198
rect 116135 6196 116141 6213
rect 116112 6193 116141 6196
rect 119515 6192 119518 6218
rect 119544 6212 119547 6218
rect 119976 6213 120005 6216
rect 119976 6212 119982 6213
rect 119544 6198 119982 6212
rect 119544 6192 119547 6198
rect 119976 6196 119982 6198
rect 119999 6196 120005 6213
rect 119976 6193 120005 6196
rect 120067 6192 120070 6218
rect 120096 6212 120099 6218
rect 121770 6213 121799 6216
rect 120096 6198 120596 6212
rect 120096 6192 120099 6198
rect 100587 6164 101828 6178
rect 100587 6162 100593 6164
rect 100564 6159 100593 6162
rect 114409 6158 114412 6184
rect 114438 6178 114441 6184
rect 114870 6179 114899 6182
rect 114870 6178 114876 6179
rect 114438 6164 114876 6178
rect 114438 6158 114441 6164
rect 114870 6162 114876 6164
rect 114893 6162 114899 6179
rect 114870 6159 114899 6162
rect 115559 6158 115562 6184
rect 115588 6178 115591 6184
rect 116249 6178 116252 6184
rect 115588 6164 116252 6178
rect 115588 6158 115591 6164
rect 116249 6158 116252 6164
rect 116278 6158 116281 6184
rect 119378 6179 119407 6182
rect 119378 6162 119384 6179
rect 119401 6178 119407 6179
rect 120582 6178 120596 6198
rect 121180 6198 121562 6212
rect 121125 6178 121128 6184
rect 119401 6164 119860 6178
rect 119401 6162 119407 6164
rect 119378 6159 119407 6162
rect 98770 6145 98799 6148
rect 98272 6130 98424 6144
rect 98218 6111 98247 6114
rect 98218 6094 98224 6111
rect 98241 6094 98247 6111
rect 98218 6091 98247 6094
rect 98272 6076 98286 6130
rect 98356 6111 98385 6114
rect 98356 6110 98362 6111
rect 97398 6062 97589 6076
rect 97996 6062 98286 6076
rect 98318 6096 98362 6110
rect 97398 6042 97412 6062
rect 96892 6028 97412 6042
rect 97481 6022 97484 6048
rect 97510 6042 97513 6048
rect 98318 6042 98332 6096
rect 98356 6094 98362 6096
rect 98379 6094 98385 6111
rect 98356 6091 98385 6094
rect 98410 6076 98424 6130
rect 98770 6128 98776 6145
rect 98793 6128 98799 6145
rect 98770 6125 98799 6128
rect 100241 6124 100244 6150
rect 100270 6144 100273 6150
rect 100270 6130 100954 6144
rect 100270 6124 100273 6130
rect 98723 6110 98726 6116
rect 98679 6096 98726 6110
rect 98723 6090 98726 6096
rect 98752 6110 98755 6116
rect 99183 6110 99186 6116
rect 98752 6096 99186 6110
rect 98752 6090 98755 6096
rect 99183 6090 99186 6096
rect 99212 6090 99215 6116
rect 100287 6090 100290 6116
rect 100316 6110 100319 6116
rect 100517 6110 100520 6116
rect 100316 6096 100520 6110
rect 100316 6090 100319 6096
rect 100517 6090 100520 6096
rect 100546 6090 100549 6116
rect 100940 6114 100954 6130
rect 101023 6124 101026 6150
rect 101052 6144 101055 6150
rect 101759 6144 101762 6150
rect 101052 6130 101762 6144
rect 101052 6124 101055 6130
rect 101759 6124 101762 6130
rect 101788 6124 101791 6150
rect 102358 6145 102387 6148
rect 102358 6128 102364 6145
rect 102381 6144 102387 6145
rect 115790 6145 115819 6148
rect 102381 6130 104887 6144
rect 102381 6128 102387 6130
rect 102358 6125 102387 6128
rect 100932 6111 100961 6114
rect 100932 6094 100938 6111
rect 100955 6094 100961 6111
rect 100932 6091 100961 6094
rect 101622 6111 101651 6114
rect 101622 6094 101628 6111
rect 101645 6110 101651 6111
rect 102265 6110 102268 6116
rect 101645 6096 102268 6110
rect 101645 6094 101651 6096
rect 101622 6091 101651 6094
rect 102265 6090 102268 6096
rect 102294 6090 102297 6116
rect 102366 6076 102380 6125
rect 104873 6110 104887 6130
rect 113774 6130 115720 6144
rect 113774 6114 113788 6130
rect 113766 6111 113795 6114
rect 113766 6110 113772 6111
rect 104873 6096 113772 6110
rect 113766 6094 113772 6096
rect 113789 6094 113795 6111
rect 114961 6110 114964 6116
rect 114917 6096 114964 6110
rect 113766 6091 113795 6094
rect 114961 6090 114964 6096
rect 114990 6110 114993 6116
rect 115651 6110 115654 6116
rect 114990 6096 115654 6110
rect 114990 6090 114993 6096
rect 115651 6090 115654 6096
rect 115680 6090 115683 6116
rect 102495 6076 102498 6082
rect 98410 6062 102380 6076
rect 102475 6062 102498 6076
rect 102495 6056 102498 6062
rect 102524 6056 102527 6082
rect 115421 6076 115424 6082
rect 102550 6062 102741 6076
rect 114517 6062 115424 6076
rect 98401 6042 98404 6048
rect 97510 6028 98332 6042
rect 98381 6028 98404 6042
rect 97510 6022 97513 6028
rect 98401 6022 98404 6028
rect 98430 6022 98433 6048
rect 98493 6042 98496 6048
rect 98473 6028 98496 6042
rect 98493 6022 98496 6028
rect 98522 6022 98525 6048
rect 98677 6042 98680 6048
rect 98657 6028 98680 6042
rect 98677 6022 98680 6028
rect 98706 6022 98709 6048
rect 101438 6043 101467 6046
rect 101438 6026 101444 6043
rect 101461 6042 101467 6043
rect 101529 6042 101532 6048
rect 101461 6028 101532 6042
rect 101461 6026 101467 6028
rect 101438 6023 101467 6026
rect 101529 6022 101532 6028
rect 101558 6022 101561 6048
rect 101668 6043 101697 6046
rect 101668 6026 101674 6043
rect 101691 6042 101697 6043
rect 101713 6042 101716 6048
rect 101691 6028 101716 6042
rect 101691 6026 101697 6028
rect 101668 6023 101697 6026
rect 101713 6022 101716 6028
rect 101742 6022 101745 6048
rect 102127 6022 102130 6048
rect 102156 6042 102159 6048
rect 102550 6042 102564 6062
rect 115421 6056 115424 6062
rect 115450 6056 115453 6082
rect 115559 6056 115562 6082
rect 115588 6076 115591 6082
rect 115706 6076 115720 6130
rect 115790 6128 115796 6145
rect 115813 6144 115819 6145
rect 115835 6144 115838 6150
rect 115813 6130 115838 6144
rect 115813 6128 115819 6130
rect 115790 6125 115819 6128
rect 115835 6124 115838 6130
rect 115864 6124 115867 6150
rect 119423 6124 119426 6150
rect 119452 6144 119455 6150
rect 119653 6144 119656 6150
rect 119452 6130 119656 6144
rect 119452 6124 119455 6130
rect 119653 6124 119656 6130
rect 119682 6124 119685 6150
rect 116065 6110 116068 6116
rect 116021 6096 116068 6110
rect 116065 6090 116068 6096
rect 116094 6110 116097 6116
rect 116525 6110 116528 6116
rect 116094 6096 116528 6110
rect 116094 6090 116097 6096
rect 116525 6090 116528 6096
rect 116554 6090 116557 6116
rect 119009 6110 119012 6116
rect 118989 6096 119012 6110
rect 119009 6090 119012 6096
rect 119038 6090 119041 6116
rect 119193 6090 119196 6116
rect 119222 6110 119225 6116
rect 119561 6110 119564 6116
rect 119222 6096 119564 6110
rect 119222 6090 119225 6096
rect 119561 6090 119564 6096
rect 119590 6090 119593 6116
rect 119608 6111 119637 6114
rect 119608 6094 119614 6111
rect 119631 6110 119637 6111
rect 119745 6110 119748 6116
rect 119631 6096 119748 6110
rect 119631 6094 119637 6096
rect 119608 6091 119637 6094
rect 119745 6090 119748 6096
rect 119774 6090 119777 6116
rect 119846 6110 119860 6164
rect 119984 6164 120504 6178
rect 120582 6164 121128 6178
rect 119984 6150 119998 6164
rect 119975 6124 119978 6150
rect 120004 6124 120007 6150
rect 120490 6144 120504 6164
rect 121125 6158 121128 6164
rect 121154 6158 121157 6184
rect 121180 6182 121194 6198
rect 121172 6179 121201 6182
rect 121172 6162 121178 6179
rect 121195 6162 121201 6179
rect 121493 6178 121496 6184
rect 121172 6159 121201 6162
rect 121364 6164 121496 6178
rect 120712 6145 120741 6148
rect 120712 6144 120718 6145
rect 120490 6130 120718 6144
rect 120712 6128 120718 6130
rect 120735 6144 120741 6145
rect 120735 6130 121148 6144
rect 120735 6128 120741 6130
rect 120712 6125 120741 6128
rect 121134 6118 121148 6130
rect 121217 6124 121220 6150
rect 121246 6144 121249 6150
rect 121364 6144 121378 6164
rect 121493 6158 121496 6164
rect 121522 6158 121525 6184
rect 121402 6145 121431 6148
rect 121402 6144 121408 6145
rect 121246 6130 121408 6144
rect 121246 6124 121249 6130
rect 121402 6128 121408 6130
rect 121425 6128 121431 6145
rect 121402 6125 121431 6128
rect 121447 6124 121450 6150
rect 121476 6144 121479 6150
rect 121476 6130 121522 6144
rect 121476 6124 121479 6130
rect 120068 6111 120097 6114
rect 120068 6110 120074 6111
rect 119846 6096 120074 6110
rect 120068 6094 120074 6096
rect 120091 6094 120097 6111
rect 120068 6091 120097 6094
rect 120620 6111 120649 6114
rect 120620 6094 120626 6111
rect 120643 6110 120649 6111
rect 121079 6110 121082 6116
rect 120643 6096 121082 6110
rect 120643 6094 120649 6096
rect 120620 6091 120649 6094
rect 121079 6090 121082 6096
rect 121108 6090 121111 6116
rect 121134 6110 121194 6118
rect 121134 6108 121424 6110
rect 121456 6108 121470 6124
rect 121134 6104 121470 6108
rect 121180 6096 121470 6104
rect 121548 6110 121562 6198
rect 121770 6196 121776 6213
rect 121793 6212 121799 6213
rect 121815 6212 121818 6218
rect 121793 6198 121818 6212
rect 121793 6196 121799 6198
rect 121770 6193 121799 6196
rect 121815 6192 121818 6198
rect 121844 6192 121847 6218
rect 122091 6212 122094 6218
rect 122071 6198 122094 6212
rect 122091 6192 122094 6198
rect 122120 6192 122123 6218
rect 125542 6213 125571 6216
rect 125542 6196 125548 6213
rect 125565 6212 125571 6213
rect 125679 6212 125682 6218
rect 125565 6198 125682 6212
rect 125565 6196 125571 6198
rect 125542 6193 125571 6196
rect 125679 6192 125682 6198
rect 125708 6192 125711 6218
rect 125955 6192 125958 6218
rect 125984 6212 125987 6218
rect 125984 6198 128140 6212
rect 125984 6192 125987 6198
rect 125725 6158 125728 6184
rect 125754 6178 125757 6184
rect 126047 6178 126050 6184
rect 125754 6164 126050 6178
rect 125754 6158 125757 6164
rect 126047 6158 126050 6164
rect 126076 6158 126079 6184
rect 127151 6178 127154 6184
rect 127107 6164 127154 6178
rect 127151 6158 127154 6164
rect 127180 6178 127183 6184
rect 127611 6178 127614 6184
rect 127180 6164 127614 6178
rect 127180 6158 127183 6164
rect 127611 6158 127614 6164
rect 127640 6158 127643 6184
rect 121585 6124 121588 6150
rect 121614 6144 121617 6150
rect 121614 6130 122206 6144
rect 121614 6124 121617 6130
rect 122192 6114 122206 6130
rect 124161 6124 124164 6150
rect 124190 6144 124193 6150
rect 124621 6144 124624 6150
rect 124190 6130 124624 6144
rect 124190 6124 124193 6130
rect 124621 6124 124624 6130
rect 124650 6124 124653 6150
rect 126278 6145 126307 6148
rect 126278 6144 126284 6145
rect 125573 6130 126284 6144
rect 121862 6111 121891 6114
rect 121862 6110 121868 6111
rect 121548 6096 121868 6110
rect 121410 6094 121470 6096
rect 121862 6094 121868 6096
rect 121885 6094 121891 6111
rect 121862 6091 121891 6094
rect 122184 6111 122213 6114
rect 122184 6094 122190 6111
rect 122207 6094 122213 6111
rect 125573 6110 125587 6130
rect 126278 6128 126284 6130
rect 126301 6144 126307 6145
rect 127658 6145 127687 6148
rect 126301 6130 127634 6144
rect 126301 6128 126307 6130
rect 126278 6125 126307 6128
rect 122184 6091 122213 6094
rect 124193 6096 125587 6110
rect 124193 6076 124207 6096
rect 125633 6090 125636 6116
rect 125662 6110 125665 6116
rect 125955 6110 125958 6116
rect 125662 6096 125684 6110
rect 125935 6096 125958 6110
rect 125662 6090 125665 6096
rect 125955 6090 125958 6096
rect 125984 6090 125987 6116
rect 127565 6110 127568 6116
rect 127545 6096 127568 6110
rect 127565 6090 127568 6096
rect 127594 6090 127597 6116
rect 124529 6076 124532 6082
rect 115588 6062 115674 6076
rect 115706 6062 124207 6076
rect 124509 6062 124532 6076
rect 115588 6056 115591 6062
rect 102156 6028 102564 6042
rect 102156 6022 102159 6028
rect 114409 6022 114412 6048
rect 114438 6042 114441 6048
rect 114640 6043 114669 6046
rect 114640 6042 114646 6043
rect 114438 6028 114646 6042
rect 114438 6022 114441 6028
rect 114640 6026 114646 6028
rect 114663 6026 114669 6043
rect 114640 6023 114669 6026
rect 115468 6043 115497 6046
rect 115468 6026 115474 6043
rect 115491 6042 115497 6043
rect 115605 6042 115608 6048
rect 115491 6028 115608 6042
rect 115491 6026 115497 6028
rect 115468 6023 115497 6026
rect 115605 6022 115608 6028
rect 115634 6022 115637 6048
rect 115660 6046 115674 6062
rect 124529 6056 124532 6062
rect 124558 6056 124561 6082
rect 124621 6056 124624 6082
rect 124650 6076 124653 6082
rect 125964 6076 125978 6090
rect 124650 6062 125978 6076
rect 126416 6077 126445 6080
rect 124650 6056 124653 6062
rect 126416 6060 126422 6077
rect 126439 6076 126445 6077
rect 126553 6076 126556 6082
rect 126439 6062 126556 6076
rect 126439 6060 126445 6062
rect 126416 6057 126445 6060
rect 126553 6056 126556 6062
rect 126582 6056 126585 6082
rect 127620 6076 127634 6130
rect 127658 6128 127664 6145
rect 127681 6144 127687 6145
rect 127795 6144 127798 6150
rect 127681 6130 127798 6144
rect 127681 6128 127687 6130
rect 127658 6125 127687 6128
rect 127795 6124 127798 6130
rect 127824 6124 127827 6150
rect 128126 6144 128140 6198
rect 128255 6192 128258 6218
rect 128284 6212 128287 6218
rect 128440 6213 128469 6216
rect 128440 6212 128446 6213
rect 128284 6198 128446 6212
rect 128284 6192 128287 6198
rect 128440 6196 128446 6198
rect 128463 6196 128469 6213
rect 131245 6212 131248 6218
rect 131225 6198 131248 6212
rect 128440 6193 128469 6196
rect 131245 6192 131248 6198
rect 131274 6192 131277 6218
rect 132304 6213 132333 6216
rect 132304 6196 132310 6213
rect 132327 6212 132333 6213
rect 132763 6212 132766 6218
rect 132327 6198 132766 6212
rect 132327 6196 132333 6198
rect 132304 6193 132333 6196
rect 132763 6192 132766 6198
rect 132792 6192 132795 6218
rect 134005 6212 134008 6218
rect 132956 6198 134008 6212
rect 128164 6179 128193 6182
rect 128164 6162 128170 6179
rect 128187 6178 128193 6179
rect 128485 6178 128488 6184
rect 128187 6164 128488 6178
rect 128187 6162 128193 6164
rect 128164 6159 128193 6162
rect 128485 6158 128488 6164
rect 128514 6158 128517 6184
rect 132028 6179 132057 6182
rect 132028 6162 132034 6179
rect 132051 6178 132057 6179
rect 132487 6178 132490 6184
rect 132051 6164 132490 6178
rect 132051 6162 132057 6164
rect 132028 6159 132057 6162
rect 132487 6158 132490 6164
rect 132516 6158 132519 6184
rect 132956 6178 132970 6198
rect 134005 6192 134008 6198
rect 134034 6192 134037 6218
rect 134189 6192 134192 6218
rect 134218 6212 134221 6218
rect 135523 6212 135526 6218
rect 134218 6198 135040 6212
rect 135503 6198 135526 6212
rect 134218 6192 134221 6198
rect 132542 6164 132970 6178
rect 135026 6178 135040 6198
rect 135523 6192 135526 6198
rect 135552 6192 135555 6218
rect 152727 6212 152730 6218
rect 152707 6198 152730 6212
rect 152727 6192 152730 6198
rect 152756 6192 152759 6218
rect 135846 6179 135875 6182
rect 135846 6178 135852 6179
rect 135026 6164 135852 6178
rect 130923 6144 130926 6150
rect 128126 6130 130926 6144
rect 130923 6124 130926 6130
rect 130952 6124 130955 6150
rect 131199 6124 131202 6150
rect 131228 6144 131231 6150
rect 131228 6130 132004 6144
rect 131228 6124 131231 6130
rect 128117 6110 128120 6116
rect 128097 6096 128120 6110
rect 128117 6090 128120 6096
rect 128146 6090 128149 6116
rect 128163 6090 128166 6116
rect 128192 6110 128195 6116
rect 128532 6111 128561 6114
rect 128532 6110 128538 6111
rect 128192 6096 128538 6110
rect 128192 6090 128195 6096
rect 128532 6094 128538 6096
rect 128555 6094 128561 6111
rect 128532 6091 128561 6094
rect 131338 6111 131367 6114
rect 131338 6094 131344 6111
rect 131361 6110 131367 6111
rect 131521 6110 131524 6116
rect 131361 6096 131524 6110
rect 131361 6094 131367 6096
rect 131338 6091 131367 6094
rect 131521 6090 131524 6096
rect 131550 6090 131553 6116
rect 131990 6114 132004 6130
rect 132073 6124 132076 6150
rect 132102 6144 132105 6150
rect 132542 6144 132556 6164
rect 132102 6130 132556 6144
rect 132102 6124 132105 6130
rect 132579 6124 132582 6150
rect 132608 6144 132611 6150
rect 132608 6130 132694 6144
rect 132608 6124 132611 6130
rect 131982 6111 132011 6114
rect 131982 6094 131988 6111
rect 132005 6110 132011 6111
rect 132165 6110 132168 6116
rect 132005 6096 132168 6110
rect 132005 6094 132011 6096
rect 131982 6091 132011 6094
rect 132165 6090 132168 6096
rect 132194 6090 132197 6116
rect 132396 6111 132425 6114
rect 132396 6094 132402 6111
rect 132419 6110 132425 6111
rect 132680 6110 132694 6130
rect 132809 6124 132812 6150
rect 132838 6144 132841 6150
rect 132956 6148 132970 6164
rect 135846 6162 135852 6164
rect 135869 6162 135875 6179
rect 135846 6159 135875 6162
rect 132856 6145 132885 6148
rect 132856 6144 132862 6145
rect 132838 6130 132862 6144
rect 132838 6124 132841 6130
rect 132856 6128 132862 6130
rect 132879 6128 132885 6145
rect 132856 6125 132885 6128
rect 132948 6145 132977 6148
rect 132948 6128 132954 6145
rect 132971 6128 132977 6145
rect 134374 6145 134403 6148
rect 134374 6144 134380 6145
rect 132948 6125 132977 6128
rect 133278 6130 134380 6144
rect 133278 6114 133292 6130
rect 134374 6128 134380 6130
rect 134397 6144 134403 6145
rect 134557 6144 134560 6150
rect 134397 6130 134560 6144
rect 134397 6128 134403 6130
rect 134374 6125 134403 6128
rect 134557 6124 134560 6130
rect 134586 6124 134589 6150
rect 134833 6124 134836 6150
rect 134862 6144 134865 6150
rect 135569 6144 135572 6150
rect 134862 6130 135572 6144
rect 134862 6124 134865 6130
rect 135569 6124 135572 6130
rect 135598 6124 135601 6150
rect 136121 6144 136124 6150
rect 136101 6130 136124 6144
rect 136121 6124 136124 6130
rect 136150 6144 136153 6150
rect 136397 6144 136400 6150
rect 136150 6130 136400 6144
rect 136150 6124 136153 6130
rect 136397 6124 136400 6130
rect 136426 6124 136429 6150
rect 133270 6111 133299 6114
rect 133270 6110 133276 6111
rect 132419 6096 132648 6110
rect 132680 6096 133276 6110
rect 132419 6094 132425 6096
rect 132396 6091 132425 6094
rect 132579 6076 132582 6082
rect 127029 6062 127542 6076
rect 127620 6062 128232 6076
rect 127528 6048 127542 6062
rect 115652 6043 115681 6046
rect 115652 6026 115658 6043
rect 115675 6026 115681 6043
rect 115652 6023 115681 6026
rect 115697 6022 115700 6048
rect 115726 6042 115729 6048
rect 115881 6042 115884 6048
rect 115726 6028 115884 6042
rect 115726 6022 115729 6028
rect 115881 6022 115884 6028
rect 115910 6022 115913 6048
rect 116525 6022 116528 6048
rect 116554 6042 116557 6048
rect 119102 6043 119131 6046
rect 119102 6042 119108 6043
rect 116554 6028 119108 6042
rect 116554 6022 116557 6028
rect 119102 6026 119108 6028
rect 119125 6026 119131 6043
rect 120435 6042 120438 6048
rect 120415 6028 120438 6042
rect 119102 6023 119131 6026
rect 120435 6022 120438 6028
rect 120464 6022 120467 6048
rect 120666 6043 120695 6046
rect 120666 6026 120672 6043
rect 120689 6042 120695 6043
rect 120757 6042 120760 6048
rect 120689 6028 120760 6042
rect 120689 6026 120695 6028
rect 120666 6023 120695 6026
rect 120757 6022 120760 6028
rect 120786 6042 120789 6048
rect 121263 6042 121266 6048
rect 120786 6028 121266 6042
rect 120786 6022 120789 6028
rect 121263 6022 121266 6028
rect 121292 6022 121295 6048
rect 121356 6043 121385 6046
rect 121356 6026 121362 6043
rect 121379 6042 121385 6043
rect 122045 6042 122048 6048
rect 121379 6028 122048 6042
rect 121379 6026 121385 6028
rect 121356 6023 121385 6026
rect 122045 6022 122048 6028
rect 122074 6022 122077 6048
rect 127197 6022 127200 6048
rect 127226 6042 127229 6048
rect 127382 6043 127411 6046
rect 127382 6042 127388 6043
rect 127226 6028 127388 6042
rect 127226 6022 127229 6028
rect 127382 6026 127388 6028
rect 127405 6026 127411 6043
rect 127382 6023 127411 6026
rect 127519 6022 127522 6048
rect 127548 6022 127551 6048
rect 127611 6022 127614 6048
rect 127640 6042 127643 6048
rect 128163 6042 128166 6048
rect 127640 6028 128166 6042
rect 127640 6022 127643 6028
rect 128163 6022 128166 6028
rect 128192 6022 128195 6048
rect 128218 6042 128232 6062
rect 131783 6062 132582 6076
rect 131783 6042 131797 6062
rect 132579 6056 132582 6062
rect 132608 6056 132611 6082
rect 132634 6046 132648 6096
rect 133270 6094 133276 6096
rect 133293 6094 133299 6111
rect 133270 6091 133299 6094
rect 134051 6090 134054 6116
rect 134080 6110 134083 6116
rect 134327 6110 134330 6116
rect 134080 6096 134330 6110
rect 134080 6090 134083 6096
rect 134327 6090 134330 6096
rect 134356 6090 134359 6116
rect 135478 6111 135507 6114
rect 135478 6110 135484 6111
rect 135164 6096 135484 6110
rect 132810 6077 132839 6080
rect 132810 6060 132816 6077
rect 132833 6076 132839 6077
rect 133407 6076 133410 6082
rect 132833 6062 133338 6076
rect 133387 6062 133410 6076
rect 132833 6060 132839 6062
rect 132810 6057 132839 6060
rect 128218 6028 131797 6042
rect 132626 6043 132655 6046
rect 132626 6026 132632 6043
rect 132649 6026 132655 6043
rect 133324 6042 133338 6062
rect 133407 6056 133410 6062
rect 133436 6056 133439 6082
rect 133637 6056 133640 6082
rect 133666 6056 133669 6082
rect 134097 6056 134100 6082
rect 134126 6076 134129 6082
rect 134512 6077 134541 6080
rect 134512 6076 134518 6077
rect 134126 6062 134518 6076
rect 134126 6056 134129 6062
rect 134512 6060 134518 6062
rect 134535 6060 134541 6077
rect 134512 6057 134541 6060
rect 134741 6056 134744 6082
rect 134770 6056 134773 6082
rect 133499 6042 133502 6048
rect 133324 6028 133502 6042
rect 132626 6023 132655 6026
rect 133499 6022 133502 6028
rect 133528 6022 133531 6048
rect 134144 6043 134173 6046
rect 134144 6026 134150 6043
rect 134167 6042 134173 6043
rect 134235 6042 134238 6048
rect 134167 6028 134238 6042
rect 134167 6026 134173 6028
rect 134144 6023 134173 6026
rect 134235 6022 134238 6028
rect 134264 6022 134267 6048
rect 134327 6022 134330 6048
rect 134356 6042 134359 6048
rect 135164 6042 135178 6096
rect 135478 6094 135484 6096
rect 135501 6110 135507 6111
rect 135661 6110 135664 6116
rect 135501 6096 135664 6110
rect 135501 6094 135507 6096
rect 135478 6091 135507 6094
rect 135661 6090 135664 6096
rect 135690 6090 135693 6116
rect 136030 6111 136059 6114
rect 136030 6094 136036 6111
rect 136053 6110 136059 6111
rect 136443 6110 136446 6116
rect 136053 6096 136446 6110
rect 136053 6094 136059 6096
rect 136030 6091 136059 6094
rect 136443 6090 136446 6096
rect 136472 6090 136475 6116
rect 135256 6062 136098 6076
rect 134356 6028 135178 6042
rect 134356 6022 134359 6028
rect 135201 6022 135204 6048
rect 135230 6042 135233 6048
rect 135256 6046 135270 6062
rect 136084 6046 136098 6062
rect 135248 6043 135277 6046
rect 135248 6042 135254 6043
rect 135230 6028 135254 6042
rect 135230 6022 135233 6028
rect 135248 6026 135254 6028
rect 135271 6026 135277 6043
rect 135248 6023 135277 6026
rect 136076 6043 136105 6046
rect 136076 6026 136082 6043
rect 136099 6042 136105 6043
rect 142377 6042 142380 6048
rect 136099 6028 142380 6042
rect 136099 6026 136105 6028
rect 136076 6023 136105 6026
rect 142377 6022 142380 6028
rect 142406 6022 142409 6048
rect 552 5997 152904 6008
rect 552 5971 38574 5997
rect 38600 5971 38606 5997
rect 38632 5971 38638 5997
rect 38664 5971 38670 5997
rect 38696 5971 38702 5997
rect 38728 5971 76673 5997
rect 76699 5971 76705 5997
rect 76731 5971 76737 5997
rect 76763 5971 76769 5997
rect 76795 5971 76801 5997
rect 76827 5971 114772 5997
rect 114798 5971 114804 5997
rect 114830 5971 114836 5997
rect 114862 5971 114868 5997
rect 114894 5971 114900 5997
rect 114926 5971 152904 5997
rect 552 5960 152904 5971
rect 13900 5941 13929 5944
rect 13900 5924 13906 5941
rect 13923 5940 13929 5941
rect 14543 5940 14546 5946
rect 13923 5926 14546 5940
rect 13923 5924 13929 5926
rect 13900 5921 13929 5924
rect 14543 5920 14546 5926
rect 14572 5920 14575 5946
rect 14727 5920 14730 5946
rect 14756 5940 14759 5946
rect 15463 5940 15466 5946
rect 14756 5926 15466 5940
rect 14756 5920 14759 5926
rect 15463 5920 15466 5926
rect 15492 5920 15495 5946
rect 16107 5920 16110 5946
rect 16136 5940 16139 5946
rect 16292 5941 16321 5944
rect 16292 5940 16298 5941
rect 16136 5926 16298 5940
rect 16136 5920 16139 5926
rect 16292 5924 16298 5926
rect 16315 5924 16321 5941
rect 16889 5940 16892 5946
rect 16869 5926 16892 5940
rect 16292 5921 16321 5924
rect 16889 5920 16892 5926
rect 16918 5920 16921 5946
rect 17211 5940 17214 5946
rect 17191 5926 17214 5940
rect 17211 5920 17214 5926
rect 17240 5920 17243 5946
rect 17488 5941 17517 5944
rect 17488 5924 17494 5941
rect 17511 5924 17517 5941
rect 19189 5940 19192 5946
rect 19169 5926 19192 5940
rect 17488 5921 17517 5924
rect 13853 5886 13856 5912
rect 13882 5906 13885 5912
rect 13882 5892 14060 5906
rect 13882 5886 13885 5892
rect 13992 5873 14021 5876
rect 13992 5856 13998 5873
rect 14015 5856 14021 5873
rect 13992 5853 14021 5856
rect 14000 5804 14014 5853
rect 14046 5838 14060 5892
rect 14359 5886 14362 5912
rect 14388 5906 14391 5912
rect 14406 5907 14435 5910
rect 14406 5906 14412 5907
rect 14388 5892 14412 5906
rect 14388 5886 14391 5892
rect 14406 5890 14412 5892
rect 14429 5890 14435 5907
rect 14406 5887 14435 5890
rect 14497 5886 14500 5912
rect 14526 5906 14529 5912
rect 15003 5906 15006 5912
rect 14526 5892 15006 5906
rect 14526 5886 14529 5892
rect 14451 5838 14454 5844
rect 14046 5824 14454 5838
rect 14451 5818 14454 5824
rect 14480 5818 14483 5844
rect 14552 5842 14566 5892
rect 15003 5886 15006 5892
rect 15032 5886 15035 5912
rect 16015 5886 16018 5912
rect 16044 5906 16047 5912
rect 17496 5906 17510 5921
rect 19189 5920 19192 5926
rect 19218 5920 19221 5946
rect 19512 5941 19541 5944
rect 19512 5924 19518 5941
rect 19535 5940 19541 5941
rect 19787 5940 19790 5946
rect 19535 5926 19790 5940
rect 19535 5924 19541 5926
rect 19512 5921 19541 5924
rect 19787 5920 19790 5926
rect 19816 5920 19819 5946
rect 19834 5941 19863 5944
rect 19834 5924 19840 5941
rect 19857 5924 19863 5941
rect 19834 5921 19863 5924
rect 16044 5892 17510 5906
rect 16044 5886 16047 5892
rect 14773 5852 14776 5878
rect 14802 5872 14805 5878
rect 14820 5873 14849 5876
rect 14820 5872 14826 5873
rect 14802 5858 14826 5872
rect 14802 5852 14805 5858
rect 14820 5856 14826 5858
rect 14843 5856 14849 5873
rect 16199 5872 16202 5878
rect 15525 5858 16202 5872
rect 14820 5853 14849 5856
rect 16199 5852 16202 5858
rect 16228 5852 16231 5878
rect 16246 5873 16275 5876
rect 16246 5856 16252 5873
rect 16269 5872 16275 5873
rect 16844 5873 16873 5876
rect 16269 5858 16406 5872
rect 16269 5856 16275 5858
rect 16246 5853 16275 5856
rect 14544 5839 14573 5842
rect 14544 5822 14550 5839
rect 14567 5822 14573 5839
rect 14957 5838 14960 5844
rect 14937 5824 14960 5838
rect 14544 5819 14573 5822
rect 14957 5818 14960 5824
rect 14986 5818 14989 5844
rect 16254 5838 16268 5853
rect 15472 5824 16268 5838
rect 14000 5790 14888 5804
rect 14221 5770 14224 5776
rect 14201 5756 14224 5770
rect 14221 5750 14224 5756
rect 14250 5750 14253 5776
rect 14874 5770 14888 5790
rect 15472 5770 15486 5824
rect 16291 5818 16294 5844
rect 16320 5838 16323 5844
rect 16338 5839 16367 5842
rect 16338 5838 16344 5839
rect 16320 5824 16344 5838
rect 16320 5818 16323 5824
rect 16338 5822 16344 5824
rect 16361 5822 16367 5839
rect 16392 5838 16406 5858
rect 16844 5856 16850 5873
rect 16867 5872 16873 5873
rect 17166 5873 17195 5876
rect 17166 5872 17172 5873
rect 16867 5858 17172 5872
rect 16867 5856 16873 5858
rect 16844 5853 16873 5856
rect 17166 5856 17172 5858
rect 17189 5872 17195 5873
rect 17349 5872 17352 5878
rect 17189 5858 17352 5872
rect 17189 5856 17195 5858
rect 17166 5853 17195 5856
rect 17349 5852 17352 5858
rect 17378 5852 17381 5878
rect 17580 5873 17609 5876
rect 17580 5856 17586 5873
rect 17603 5856 17609 5873
rect 17580 5853 17609 5856
rect 19282 5873 19311 5876
rect 19282 5856 19288 5873
rect 19305 5856 19311 5873
rect 19282 5853 19311 5856
rect 19604 5873 19633 5876
rect 19604 5856 19610 5873
rect 19627 5872 19633 5873
rect 19842 5872 19856 5921
rect 19971 5920 19974 5946
rect 20000 5940 20003 5946
rect 20064 5941 20093 5944
rect 20064 5940 20070 5941
rect 20000 5926 20070 5940
rect 20000 5920 20003 5926
rect 20064 5924 20070 5926
rect 20087 5924 20093 5941
rect 20064 5921 20093 5924
rect 20570 5941 20599 5944
rect 20570 5924 20576 5941
rect 20593 5940 20599 5941
rect 20707 5940 20710 5946
rect 20593 5926 20710 5940
rect 20593 5924 20599 5926
rect 20570 5921 20599 5924
rect 20707 5920 20710 5926
rect 20736 5920 20739 5946
rect 20846 5941 20875 5944
rect 20846 5924 20852 5941
rect 20869 5940 20875 5941
rect 21443 5940 21446 5946
rect 20869 5926 21446 5940
rect 20869 5924 20875 5926
rect 20846 5921 20875 5924
rect 21443 5920 21446 5926
rect 21472 5920 21475 5946
rect 26319 5920 26322 5946
rect 26348 5940 26351 5946
rect 26412 5941 26441 5944
rect 26412 5940 26418 5941
rect 26348 5926 26418 5940
rect 26348 5920 26351 5926
rect 26412 5924 26418 5926
rect 26435 5924 26441 5941
rect 26825 5940 26828 5946
rect 26805 5926 26828 5940
rect 26412 5921 26441 5924
rect 26825 5920 26828 5926
rect 26854 5920 26857 5946
rect 27193 5940 27196 5946
rect 27173 5926 27196 5940
rect 27193 5920 27196 5926
rect 27222 5920 27225 5946
rect 27653 5940 27656 5946
rect 27633 5926 27656 5940
rect 27653 5920 27656 5926
rect 27682 5920 27685 5946
rect 28252 5941 28281 5944
rect 28252 5924 28258 5941
rect 28275 5940 28281 5941
rect 28297 5940 28300 5946
rect 28275 5926 28300 5940
rect 28275 5924 28281 5926
rect 28252 5921 28281 5924
rect 28297 5920 28300 5926
rect 28326 5920 28329 5946
rect 28574 5941 28603 5944
rect 28574 5924 28580 5941
rect 28597 5940 28603 5941
rect 29309 5940 29312 5946
rect 28597 5926 29312 5940
rect 28597 5924 28603 5926
rect 28574 5921 28603 5924
rect 29309 5920 29312 5926
rect 29338 5920 29341 5946
rect 37727 5920 37730 5946
rect 37756 5940 37759 5946
rect 37774 5941 37803 5944
rect 37774 5940 37780 5941
rect 37756 5926 37780 5940
rect 37756 5920 37759 5926
rect 37774 5924 37780 5926
rect 37797 5924 37803 5941
rect 37774 5921 37803 5924
rect 37819 5920 37822 5946
rect 37848 5940 37851 5946
rect 38004 5941 38033 5944
rect 38004 5940 38010 5941
rect 37848 5926 38010 5940
rect 37848 5920 37851 5926
rect 38004 5924 38010 5926
rect 38027 5924 38033 5941
rect 38004 5921 38033 5924
rect 38233 5920 38236 5946
rect 38262 5940 38265 5946
rect 38464 5941 38493 5944
rect 38464 5940 38470 5941
rect 38262 5926 38470 5940
rect 38262 5920 38265 5926
rect 38464 5924 38470 5926
rect 38487 5924 38493 5941
rect 38923 5940 38926 5946
rect 38903 5926 38926 5940
rect 38464 5921 38493 5924
rect 38923 5920 38926 5926
rect 38952 5920 38955 5946
rect 39245 5940 39248 5946
rect 39225 5926 39248 5940
rect 39245 5920 39248 5926
rect 39274 5920 39277 5946
rect 42143 5920 42146 5946
rect 42172 5940 42175 5946
rect 42190 5941 42219 5944
rect 42190 5940 42196 5941
rect 42172 5926 42196 5940
rect 42172 5920 42175 5926
rect 42190 5924 42196 5926
rect 42213 5924 42219 5941
rect 43017 5940 43020 5946
rect 42190 5921 42219 5924
rect 42520 5926 43020 5940
rect 20018 5907 20047 5910
rect 20018 5890 20024 5907
rect 20041 5906 20047 5907
rect 20339 5906 20342 5912
rect 20041 5892 20342 5906
rect 20041 5890 20047 5892
rect 20018 5887 20047 5890
rect 19627 5858 19856 5872
rect 19627 5856 19633 5858
rect 19604 5853 19633 5856
rect 17027 5838 17030 5844
rect 16392 5824 17030 5838
rect 16338 5819 16367 5822
rect 17027 5818 17030 5824
rect 17056 5818 17059 5844
rect 15555 5784 15558 5810
rect 15584 5804 15587 5810
rect 17588 5804 17602 5853
rect 19290 5838 19304 5853
rect 20026 5838 20040 5887
rect 20339 5886 20342 5892
rect 20368 5906 20371 5912
rect 20615 5906 20618 5912
rect 20368 5892 20618 5906
rect 20368 5886 20371 5892
rect 20615 5886 20618 5892
rect 20644 5886 20647 5912
rect 26871 5886 26874 5912
rect 26900 5906 26903 5912
rect 26900 5892 28228 5906
rect 26900 5886 26903 5892
rect 20155 5852 20158 5878
rect 20184 5872 20187 5878
rect 20524 5873 20553 5876
rect 20524 5872 20530 5873
rect 20184 5858 20530 5872
rect 20184 5852 20187 5858
rect 20524 5856 20530 5858
rect 20547 5872 20553 5873
rect 20938 5873 20967 5876
rect 20547 5858 20707 5872
rect 20547 5856 20553 5858
rect 20524 5853 20553 5856
rect 20693 5844 20707 5858
rect 20938 5856 20944 5873
rect 20961 5872 20967 5873
rect 21397 5872 21400 5878
rect 20961 5858 21400 5872
rect 20961 5856 20967 5858
rect 20938 5853 20967 5856
rect 21397 5852 21400 5858
rect 21426 5852 21429 5878
rect 21444 5873 21473 5876
rect 21444 5856 21450 5873
rect 21467 5872 21473 5873
rect 21489 5872 21492 5878
rect 21467 5858 21492 5872
rect 21467 5856 21473 5858
rect 21444 5853 21473 5856
rect 21489 5852 21492 5858
rect 21518 5872 21521 5878
rect 26503 5872 26506 5878
rect 21518 5858 21742 5872
rect 26483 5858 26506 5872
rect 21518 5852 21521 5858
rect 19290 5824 20040 5838
rect 20110 5839 20139 5842
rect 20110 5822 20116 5839
rect 20133 5838 20139 5839
rect 20477 5838 20480 5844
rect 20133 5824 20480 5838
rect 20133 5822 20139 5824
rect 20110 5819 20139 5822
rect 20477 5818 20480 5824
rect 20506 5818 20509 5844
rect 20693 5824 20710 5844
rect 20707 5818 20710 5824
rect 20736 5838 20739 5844
rect 21536 5839 21565 5842
rect 21536 5838 21542 5839
rect 20736 5824 21542 5838
rect 20736 5818 20739 5824
rect 21536 5822 21542 5824
rect 21559 5822 21565 5839
rect 21536 5819 21565 5822
rect 21728 5808 21742 5858
rect 26503 5852 26506 5858
rect 26532 5852 26535 5878
rect 27156 5876 27170 5892
rect 28214 5876 28228 5892
rect 28711 5886 28714 5912
rect 28740 5906 28743 5912
rect 42465 5906 42468 5912
rect 28740 5892 42468 5906
rect 28740 5886 28743 5892
rect 42465 5886 42468 5892
rect 42494 5886 42497 5912
rect 26918 5873 26947 5876
rect 26918 5856 26924 5873
rect 26941 5856 26947 5873
rect 26918 5853 26947 5856
rect 27148 5873 27177 5876
rect 27148 5856 27154 5873
rect 27171 5856 27177 5873
rect 27148 5853 27177 5856
rect 28206 5873 28235 5876
rect 28206 5856 28212 5873
rect 28229 5872 28235 5873
rect 28528 5873 28557 5876
rect 28528 5872 28534 5873
rect 28229 5858 28534 5872
rect 28229 5856 28235 5858
rect 28206 5853 28235 5856
rect 28528 5856 28534 5858
rect 28551 5856 28557 5873
rect 28528 5853 28557 5856
rect 26926 5838 26940 5853
rect 27331 5838 27334 5844
rect 26926 5824 27334 5838
rect 27331 5818 27334 5824
rect 27360 5838 27363 5844
rect 27700 5839 27729 5842
rect 27700 5838 27706 5839
rect 27360 5824 27706 5838
rect 27360 5818 27363 5824
rect 27700 5822 27706 5824
rect 27723 5822 27729 5839
rect 27791 5838 27794 5844
rect 27771 5824 27794 5838
rect 27700 5819 27729 5822
rect 27791 5818 27794 5824
rect 27820 5818 27823 5844
rect 27929 5818 27932 5844
rect 27958 5838 27961 5844
rect 28720 5838 28734 5886
rect 37958 5873 37987 5876
rect 37958 5856 37964 5873
rect 37981 5872 37987 5873
rect 38003 5872 38006 5878
rect 37981 5858 38006 5872
rect 37981 5856 37987 5858
rect 37958 5853 37987 5856
rect 38003 5852 38006 5858
rect 38032 5852 38035 5878
rect 38141 5852 38144 5878
rect 38170 5872 38173 5878
rect 38556 5873 38585 5876
rect 38556 5872 38562 5873
rect 38170 5858 38562 5872
rect 38170 5852 38173 5858
rect 38556 5856 38562 5858
rect 38579 5856 38585 5873
rect 38556 5853 38585 5856
rect 38878 5873 38907 5876
rect 38878 5856 38884 5873
rect 38901 5872 38907 5873
rect 39291 5872 39294 5878
rect 38901 5858 39294 5872
rect 38901 5856 38907 5858
rect 38878 5853 38907 5856
rect 39291 5852 39294 5858
rect 39320 5852 39323 5878
rect 39338 5873 39367 5876
rect 39338 5856 39344 5873
rect 39361 5872 39367 5873
rect 40717 5872 40720 5878
rect 39361 5858 40720 5872
rect 39361 5856 39367 5858
rect 39338 5853 39367 5856
rect 40717 5852 40720 5858
rect 40746 5852 40749 5878
rect 42282 5873 42311 5876
rect 42282 5856 42288 5873
rect 42305 5872 42311 5873
rect 42520 5872 42534 5926
rect 43017 5920 43020 5926
rect 43046 5920 43049 5946
rect 43063 5920 43066 5946
rect 43092 5940 43095 5946
rect 43570 5941 43599 5944
rect 43570 5940 43576 5941
rect 43092 5926 43576 5940
rect 43092 5920 43095 5926
rect 43570 5924 43576 5926
rect 43593 5924 43599 5941
rect 43937 5940 43940 5946
rect 43917 5926 43940 5940
rect 43570 5921 43599 5924
rect 43937 5920 43940 5926
rect 43966 5920 43969 5946
rect 44444 5941 44473 5944
rect 44444 5924 44450 5941
rect 44467 5940 44473 5941
rect 44765 5940 44768 5946
rect 44467 5926 44768 5940
rect 44467 5924 44473 5926
rect 44444 5921 44473 5924
rect 44765 5920 44768 5926
rect 44794 5920 44797 5946
rect 49825 5920 49828 5946
rect 49854 5940 49857 5946
rect 50102 5941 50131 5944
rect 50102 5940 50108 5941
rect 49854 5926 50108 5940
rect 49854 5920 49857 5926
rect 50102 5924 50108 5926
rect 50125 5924 50131 5941
rect 50469 5940 50472 5946
rect 50449 5926 50472 5940
rect 50102 5921 50131 5924
rect 50469 5920 50472 5926
rect 50498 5920 50501 5946
rect 50930 5941 50959 5944
rect 50930 5924 50936 5941
rect 50953 5940 50959 5941
rect 51527 5940 51530 5946
rect 50953 5926 51530 5940
rect 50953 5924 50959 5926
rect 50930 5921 50959 5924
rect 51527 5920 51530 5926
rect 51556 5920 51559 5946
rect 51757 5920 51760 5946
rect 51786 5940 51789 5946
rect 56909 5940 56912 5946
rect 51786 5926 56587 5940
rect 56889 5926 56912 5940
rect 51786 5920 51789 5926
rect 42649 5886 42652 5912
rect 42678 5906 42681 5912
rect 56573 5906 56587 5926
rect 56909 5920 56912 5926
rect 56938 5920 56941 5946
rect 57139 5920 57142 5946
rect 57168 5940 57171 5946
rect 57508 5941 57537 5944
rect 57508 5940 57514 5941
rect 57168 5926 57514 5940
rect 57168 5920 57171 5926
rect 57508 5924 57514 5926
rect 57531 5940 57537 5941
rect 57829 5940 57832 5946
rect 57531 5926 57832 5940
rect 57531 5924 57537 5926
rect 57508 5921 57537 5924
rect 57829 5920 57832 5926
rect 57858 5920 57861 5946
rect 58106 5941 58135 5944
rect 58106 5924 58112 5941
rect 58129 5940 58135 5941
rect 58381 5940 58384 5946
rect 58129 5926 58384 5940
rect 58129 5924 58135 5926
rect 58106 5921 58135 5924
rect 58381 5920 58384 5926
rect 58410 5920 58413 5946
rect 58474 5941 58503 5944
rect 58474 5924 58480 5941
rect 58497 5940 58503 5941
rect 58657 5940 58660 5946
rect 58497 5926 58660 5940
rect 58497 5924 58503 5926
rect 58474 5921 58503 5924
rect 58657 5920 58660 5926
rect 58686 5920 58689 5946
rect 58796 5941 58825 5944
rect 58796 5924 58802 5941
rect 58819 5940 58825 5941
rect 59393 5940 59396 5946
rect 58819 5926 59396 5940
rect 58819 5924 58825 5926
rect 58796 5921 58825 5924
rect 59393 5920 59396 5926
rect 59422 5920 59425 5946
rect 64683 5940 64686 5946
rect 64663 5926 64686 5940
rect 64683 5920 64686 5926
rect 64712 5920 64715 5946
rect 65143 5920 65146 5946
rect 65172 5940 65175 5946
rect 65236 5941 65265 5944
rect 65236 5940 65242 5941
rect 65172 5926 65242 5940
rect 65172 5920 65175 5926
rect 65236 5924 65242 5926
rect 65259 5924 65265 5941
rect 65465 5940 65468 5946
rect 65445 5926 65468 5940
rect 65236 5921 65265 5924
rect 65465 5920 65468 5926
rect 65494 5920 65497 5946
rect 65557 5920 65560 5946
rect 65586 5940 65589 5946
rect 66202 5941 66231 5944
rect 66202 5940 66208 5941
rect 65586 5926 66208 5940
rect 65586 5920 65589 5926
rect 66202 5924 66208 5926
rect 66225 5924 66231 5941
rect 66202 5921 66231 5924
rect 68869 5920 68872 5946
rect 68898 5940 68901 5946
rect 75539 5940 75542 5946
rect 68898 5926 75470 5940
rect 75519 5926 75542 5940
rect 68898 5920 68901 5926
rect 57277 5906 57280 5912
rect 42678 5892 54126 5906
rect 56573 5892 57280 5906
rect 42678 5886 42681 5892
rect 42305 5858 42534 5872
rect 42604 5873 42633 5876
rect 42305 5856 42311 5858
rect 42282 5853 42311 5856
rect 42604 5856 42610 5873
rect 42627 5856 42633 5873
rect 42604 5853 42633 5856
rect 27958 5824 28734 5838
rect 27958 5818 27961 5824
rect 37497 5818 37500 5844
rect 37526 5838 37529 5844
rect 38096 5839 38125 5842
rect 38096 5838 38102 5839
rect 37526 5824 38102 5838
rect 37526 5818 37529 5824
rect 38096 5822 38102 5824
rect 38119 5838 38125 5839
rect 38463 5838 38466 5844
rect 38119 5824 38466 5838
rect 38119 5822 38125 5824
rect 38096 5819 38125 5822
rect 38463 5818 38466 5824
rect 38492 5818 38495 5844
rect 42005 5818 42008 5844
rect 42034 5838 42037 5844
rect 42612 5838 42626 5853
rect 42879 5852 42882 5878
rect 42908 5872 42911 5878
rect 43064 5873 43093 5876
rect 43064 5872 43070 5873
rect 42908 5858 43070 5872
rect 42908 5852 42911 5858
rect 43064 5856 43070 5858
rect 43087 5856 43093 5873
rect 43064 5853 43093 5856
rect 43477 5852 43480 5878
rect 43506 5872 43509 5878
rect 43892 5873 43921 5876
rect 43506 5858 43528 5872
rect 43506 5852 43509 5858
rect 43892 5856 43898 5873
rect 43915 5872 43921 5873
rect 44398 5873 44427 5876
rect 43915 5858 43960 5872
rect 43915 5856 43921 5858
rect 43892 5853 43921 5856
rect 43155 5838 43158 5844
rect 42034 5824 42626 5838
rect 43135 5824 43158 5838
rect 42034 5818 42037 5824
rect 43155 5818 43158 5824
rect 43184 5818 43187 5844
rect 43946 5838 43960 5858
rect 44398 5856 44404 5873
rect 44421 5872 44427 5873
rect 44581 5872 44584 5878
rect 44421 5858 44584 5872
rect 44421 5856 44427 5858
rect 44398 5853 44427 5856
rect 44581 5852 44584 5858
rect 44610 5852 44613 5878
rect 50193 5872 50196 5878
rect 50173 5858 50196 5872
rect 50193 5852 50196 5858
rect 50222 5852 50225 5878
rect 50424 5873 50453 5876
rect 50424 5856 50430 5873
rect 50447 5872 50453 5873
rect 51067 5872 51070 5878
rect 50447 5858 51070 5872
rect 50447 5856 50453 5858
rect 50424 5853 50453 5856
rect 51067 5852 51070 5858
rect 51096 5852 51099 5878
rect 51574 5873 51603 5876
rect 51574 5856 51580 5873
rect 51597 5872 51603 5873
rect 51803 5872 51806 5878
rect 51597 5858 51806 5872
rect 51597 5856 51603 5858
rect 51574 5853 51603 5856
rect 51803 5852 51806 5858
rect 51832 5852 51835 5878
rect 45225 5838 45228 5844
rect 43210 5824 43477 5838
rect 43946 5824 45228 5838
rect 15584 5790 17602 5804
rect 21720 5805 21749 5808
rect 15584 5784 15587 5790
rect 21720 5788 21726 5805
rect 21743 5804 21749 5805
rect 28021 5804 28024 5810
rect 21743 5790 28024 5804
rect 21743 5788 21749 5790
rect 21720 5785 21749 5788
rect 28021 5784 28024 5790
rect 28050 5804 28053 5810
rect 43210 5804 43224 5824
rect 28050 5790 43224 5804
rect 43463 5804 43477 5824
rect 45225 5818 45228 5824
rect 45254 5818 45257 5844
rect 50377 5818 50380 5844
rect 50406 5838 50409 5844
rect 50976 5839 51005 5842
rect 50976 5838 50982 5839
rect 50406 5824 50982 5838
rect 50406 5818 50409 5824
rect 50976 5822 50982 5824
rect 50999 5822 51005 5839
rect 50976 5819 51005 5822
rect 51021 5818 51024 5844
rect 51050 5838 51053 5844
rect 51050 5824 51072 5838
rect 51050 5818 51053 5824
rect 51159 5818 51162 5844
rect 51188 5838 51191 5844
rect 51757 5838 51760 5844
rect 51188 5824 51760 5838
rect 51188 5818 51191 5824
rect 51757 5818 51760 5824
rect 51786 5818 51789 5844
rect 54112 5838 54126 5892
rect 57277 5886 57280 5892
rect 57306 5886 57309 5912
rect 69007 5906 69010 5912
rect 57470 5892 69010 5906
rect 57001 5872 57004 5878
rect 56981 5858 57004 5872
rect 57001 5852 57004 5858
rect 57030 5852 57033 5878
rect 57470 5838 57484 5892
rect 69007 5886 69010 5892
rect 69036 5886 69039 5912
rect 74987 5906 74990 5912
rect 74911 5892 74990 5906
rect 74987 5886 74990 5892
rect 75016 5886 75019 5912
rect 75456 5906 75470 5926
rect 75539 5920 75542 5926
rect 75568 5920 75571 5946
rect 75999 5940 76002 5946
rect 75979 5926 76002 5940
rect 75999 5920 76002 5926
rect 76028 5920 76031 5946
rect 76368 5941 76397 5944
rect 76368 5924 76374 5941
rect 76391 5940 76397 5941
rect 77103 5940 77106 5946
rect 76391 5926 77106 5940
rect 76391 5924 76397 5926
rect 76368 5921 76397 5924
rect 77103 5920 77106 5926
rect 77132 5920 77135 5946
rect 78653 5926 80990 5940
rect 78653 5906 78667 5926
rect 75456 5892 78667 5906
rect 57507 5852 57510 5878
rect 57536 5872 57539 5878
rect 57554 5873 57583 5876
rect 57554 5872 57560 5873
rect 57536 5858 57560 5872
rect 57536 5852 57539 5858
rect 57554 5856 57560 5858
rect 57577 5856 57583 5873
rect 58197 5872 58200 5878
rect 58177 5858 58200 5872
rect 57554 5853 57583 5856
rect 58197 5852 58200 5858
rect 58226 5852 58229 5878
rect 58428 5873 58457 5876
rect 58428 5856 58434 5873
rect 58451 5872 58457 5873
rect 58750 5873 58779 5876
rect 58750 5872 58756 5873
rect 58451 5858 58756 5872
rect 58451 5856 58457 5858
rect 58428 5853 58457 5856
rect 58750 5856 58756 5858
rect 58773 5872 58779 5873
rect 59163 5872 59166 5878
rect 58773 5858 59166 5872
rect 58773 5856 58779 5858
rect 58750 5853 58779 5856
rect 54112 5824 57484 5838
rect 57646 5839 57675 5842
rect 57646 5822 57652 5839
rect 57669 5838 57675 5839
rect 57829 5838 57832 5844
rect 57669 5824 57832 5838
rect 57669 5822 57675 5824
rect 57646 5819 57675 5822
rect 57829 5818 57832 5824
rect 57858 5818 57861 5844
rect 57875 5818 57878 5844
rect 57904 5838 57907 5844
rect 58436 5838 58450 5853
rect 59163 5852 59166 5858
rect 59192 5852 59195 5878
rect 64177 5852 64180 5878
rect 64206 5872 64209 5878
rect 64638 5873 64667 5876
rect 64638 5872 64644 5873
rect 64206 5858 64644 5872
rect 64206 5852 64209 5858
rect 64638 5856 64644 5858
rect 64661 5872 64667 5873
rect 65143 5872 65146 5878
rect 64661 5858 65146 5872
rect 64661 5856 64667 5858
rect 64638 5853 64667 5856
rect 65143 5852 65146 5858
rect 65172 5852 65175 5878
rect 65420 5873 65449 5876
rect 65420 5856 65426 5873
rect 65443 5872 65449 5873
rect 65787 5872 65790 5878
rect 65443 5858 65790 5872
rect 65443 5856 65449 5858
rect 65420 5853 65449 5856
rect 65787 5852 65790 5858
rect 65816 5852 65819 5878
rect 65834 5873 65863 5876
rect 65834 5856 65840 5873
rect 65857 5856 65863 5873
rect 65834 5853 65863 5856
rect 57904 5824 58450 5838
rect 57904 5818 57907 5824
rect 64867 5818 64870 5844
rect 64896 5838 64899 5844
rect 65511 5838 65514 5844
rect 64896 5824 65514 5838
rect 64896 5818 64899 5824
rect 65511 5818 65514 5824
rect 65540 5818 65543 5844
rect 65842 5838 65856 5853
rect 66247 5852 66250 5878
rect 66276 5872 66279 5878
rect 66294 5873 66323 5876
rect 66294 5872 66300 5873
rect 66276 5858 66300 5872
rect 66276 5852 66279 5858
rect 66294 5856 66300 5858
rect 66317 5856 66323 5873
rect 66294 5853 66323 5856
rect 73837 5852 73840 5878
rect 73866 5872 73869 5878
rect 73884 5873 73913 5876
rect 73884 5872 73890 5873
rect 73866 5858 73890 5872
rect 73866 5852 73869 5858
rect 73884 5856 73890 5858
rect 73907 5856 73913 5873
rect 75631 5872 75634 5878
rect 75611 5858 75634 5872
rect 73884 5853 73913 5856
rect 75631 5852 75634 5858
rect 75660 5852 75663 5878
rect 76091 5872 76094 5878
rect 76071 5858 76094 5872
rect 76091 5852 76094 5858
rect 76120 5852 76123 5878
rect 76322 5873 76351 5876
rect 76322 5856 76328 5873
rect 76345 5872 76351 5873
rect 76367 5872 76370 5878
rect 76345 5858 76370 5872
rect 76345 5856 76351 5858
rect 76322 5853 76351 5856
rect 76367 5852 76370 5858
rect 76396 5852 76399 5878
rect 80553 5872 80556 5878
rect 80533 5858 80556 5872
rect 80553 5852 80556 5858
rect 80582 5852 80585 5878
rect 80875 5872 80878 5878
rect 80855 5858 80878 5872
rect 80875 5852 80878 5858
rect 80904 5852 80907 5878
rect 68869 5838 68872 5844
rect 65842 5824 68872 5838
rect 68869 5818 68872 5824
rect 68898 5818 68901 5844
rect 74159 5838 74162 5844
rect 74139 5824 74162 5838
rect 74159 5818 74162 5824
rect 74188 5818 74191 5844
rect 74297 5838 74300 5844
rect 74277 5824 74300 5838
rect 74297 5818 74300 5824
rect 74326 5818 74329 5844
rect 71629 5804 71632 5810
rect 43463 5790 71632 5804
rect 28050 5784 28053 5790
rect 71629 5784 71632 5790
rect 71658 5784 71661 5810
rect 73009 5784 73012 5810
rect 73038 5804 73041 5810
rect 73792 5805 73821 5808
rect 73792 5804 73798 5805
rect 73038 5790 73798 5804
rect 73038 5784 73041 5790
rect 73792 5788 73798 5790
rect 73815 5788 73821 5805
rect 73792 5785 73821 5788
rect 80462 5805 80491 5808
rect 80462 5788 80468 5805
rect 80485 5804 80491 5805
rect 80599 5804 80602 5810
rect 80485 5790 80602 5804
rect 80485 5788 80491 5790
rect 80462 5785 80491 5788
rect 80599 5784 80602 5790
rect 80628 5784 80631 5810
rect 80645 5784 80648 5810
rect 80674 5804 80677 5810
rect 80784 5805 80813 5808
rect 80784 5804 80790 5805
rect 80674 5790 80790 5804
rect 80674 5784 80677 5790
rect 80784 5788 80790 5790
rect 80807 5788 80813 5805
rect 80976 5804 80990 5926
rect 81013 5920 81016 5946
rect 81042 5940 81045 5946
rect 81152 5941 81181 5944
rect 81152 5940 81158 5941
rect 81042 5926 81158 5940
rect 81042 5920 81045 5926
rect 81152 5924 81158 5926
rect 81175 5924 81181 5941
rect 81152 5921 81181 5924
rect 81381 5920 81384 5946
rect 81410 5940 81413 5946
rect 81474 5941 81503 5944
rect 81474 5940 81480 5941
rect 81410 5926 81480 5940
rect 81410 5920 81413 5926
rect 81474 5924 81480 5926
rect 81497 5924 81503 5941
rect 81474 5921 81503 5924
rect 81750 5941 81779 5944
rect 81750 5924 81756 5941
rect 81773 5940 81779 5941
rect 81887 5940 81890 5946
rect 81773 5926 81890 5940
rect 81773 5924 81779 5926
rect 81750 5921 81779 5924
rect 81887 5920 81890 5926
rect 81916 5920 81919 5946
rect 82118 5941 82147 5944
rect 82118 5924 82124 5941
rect 82141 5940 82147 5941
rect 82163 5940 82166 5946
rect 82141 5926 82166 5940
rect 82141 5924 82147 5926
rect 82118 5921 82147 5924
rect 82163 5920 82166 5926
rect 82192 5920 82195 5946
rect 82439 5940 82442 5946
rect 82419 5926 82442 5940
rect 82439 5920 82442 5926
rect 82468 5920 82471 5946
rect 88236 5941 88265 5944
rect 88236 5924 88242 5941
rect 88259 5940 88265 5941
rect 88373 5940 88376 5946
rect 88259 5926 88376 5940
rect 88259 5924 88265 5926
rect 88236 5921 88265 5924
rect 88373 5920 88376 5926
rect 88402 5920 88405 5946
rect 88695 5920 88698 5946
rect 88724 5940 88727 5946
rect 88788 5941 88817 5944
rect 88788 5940 88794 5941
rect 88724 5926 88794 5940
rect 88724 5920 88727 5926
rect 88788 5924 88794 5926
rect 88811 5924 88817 5941
rect 88788 5921 88817 5924
rect 88925 5920 88928 5946
rect 88954 5940 88957 5946
rect 89018 5941 89047 5944
rect 89018 5940 89024 5941
rect 88954 5926 89024 5940
rect 88954 5920 88957 5926
rect 89018 5924 89024 5926
rect 89041 5924 89047 5941
rect 89018 5921 89047 5924
rect 89570 5941 89599 5944
rect 89570 5924 89576 5941
rect 89593 5940 89599 5941
rect 89937 5940 89940 5946
rect 89593 5926 89940 5940
rect 89593 5924 89599 5926
rect 89570 5921 89599 5924
rect 89937 5920 89940 5926
rect 89966 5920 89969 5946
rect 89983 5920 89986 5946
rect 90012 5940 90015 5946
rect 90030 5941 90059 5944
rect 90030 5940 90036 5941
rect 90012 5926 90036 5940
rect 90012 5920 90015 5926
rect 90030 5924 90036 5926
rect 90053 5924 90059 5941
rect 90030 5921 90059 5924
rect 90075 5920 90078 5946
rect 90104 5940 90107 5946
rect 94169 5940 94172 5946
rect 90104 5926 94172 5940
rect 90104 5920 90107 5926
rect 94169 5920 94172 5926
rect 94198 5920 94201 5946
rect 95412 5941 95441 5944
rect 95412 5924 95418 5941
rect 95435 5940 95441 5941
rect 95871 5940 95874 5946
rect 95435 5926 95874 5940
rect 95435 5924 95441 5926
rect 95412 5921 95441 5924
rect 95871 5920 95874 5926
rect 95900 5920 95903 5946
rect 95917 5920 95920 5946
rect 95946 5940 95949 5946
rect 97205 5940 97208 5946
rect 95946 5926 97208 5940
rect 95946 5920 95949 5926
rect 81289 5886 81292 5912
rect 81318 5906 81321 5912
rect 94767 5906 94770 5912
rect 81318 5892 94770 5906
rect 81318 5886 81321 5892
rect 94767 5886 94770 5892
rect 94796 5886 94799 5912
rect 96929 5906 96932 5912
rect 96669 5892 96932 5906
rect 96929 5886 96932 5892
rect 96958 5886 96961 5912
rect 81106 5873 81135 5876
rect 81106 5856 81112 5873
rect 81129 5872 81135 5873
rect 81428 5873 81457 5876
rect 81428 5872 81434 5873
rect 81129 5858 81434 5872
rect 81129 5856 81135 5858
rect 81106 5853 81135 5856
rect 81428 5856 81434 5858
rect 81451 5856 81457 5873
rect 81841 5872 81844 5878
rect 81821 5858 81844 5872
rect 81428 5853 81457 5856
rect 81436 5838 81450 5853
rect 81841 5852 81844 5858
rect 81870 5852 81873 5878
rect 82072 5873 82101 5876
rect 82072 5856 82078 5873
rect 82095 5872 82101 5873
rect 82394 5873 82423 5876
rect 82394 5872 82400 5873
rect 82095 5858 82400 5872
rect 82095 5856 82101 5858
rect 82072 5853 82101 5856
rect 82394 5856 82400 5858
rect 82417 5872 82423 5873
rect 83313 5872 83316 5878
rect 82417 5858 83316 5872
rect 82417 5856 82423 5858
rect 82394 5853 82423 5856
rect 81749 5838 81752 5844
rect 81436 5824 81752 5838
rect 81749 5818 81752 5824
rect 81778 5838 81781 5844
rect 82080 5838 82094 5853
rect 83313 5852 83316 5858
rect 83342 5852 83345 5878
rect 88327 5872 88330 5878
rect 88307 5858 88330 5872
rect 88327 5852 88330 5858
rect 88356 5852 88359 5878
rect 88972 5873 89001 5876
rect 88972 5856 88978 5873
rect 88995 5872 89001 5873
rect 89616 5873 89645 5876
rect 89616 5872 89622 5873
rect 88995 5858 89622 5872
rect 88995 5856 89001 5858
rect 88972 5853 89001 5856
rect 89616 5856 89622 5858
rect 89639 5872 89645 5873
rect 89937 5872 89940 5878
rect 89639 5858 89940 5872
rect 89639 5856 89645 5858
rect 89616 5853 89645 5856
rect 89937 5852 89940 5858
rect 89966 5852 89969 5878
rect 89984 5873 90013 5876
rect 89984 5856 89990 5873
rect 90007 5856 90013 5873
rect 89984 5853 90013 5856
rect 81778 5824 82094 5838
rect 81778 5818 81781 5824
rect 88557 5818 88560 5844
rect 88586 5838 88589 5844
rect 89064 5839 89093 5842
rect 89064 5838 89070 5839
rect 88586 5824 89070 5838
rect 88586 5818 88589 5824
rect 89064 5822 89070 5824
rect 89087 5838 89093 5839
rect 89662 5839 89691 5842
rect 89662 5838 89668 5839
rect 89087 5824 89668 5838
rect 89087 5822 89093 5824
rect 89064 5819 89093 5822
rect 82945 5804 82948 5810
rect 80976 5790 82948 5804
rect 80784 5785 80813 5788
rect 82945 5784 82948 5790
rect 82974 5784 82977 5810
rect 15693 5770 15696 5776
rect 14874 5756 15486 5770
rect 15673 5756 15696 5770
rect 15693 5750 15696 5756
rect 15722 5750 15725 5776
rect 16062 5771 16091 5774
rect 16062 5754 16068 5771
rect 16085 5770 16091 5771
rect 16475 5770 16478 5776
rect 16085 5756 16478 5770
rect 16085 5754 16091 5756
rect 16062 5751 16091 5754
rect 16475 5750 16478 5756
rect 16504 5750 16507 5776
rect 27470 5771 27499 5774
rect 27470 5754 27476 5771
rect 27493 5770 27499 5771
rect 27745 5770 27748 5776
rect 27493 5756 27748 5770
rect 27493 5754 27499 5756
rect 27470 5751 27499 5754
rect 27745 5750 27748 5756
rect 27774 5750 27777 5776
rect 42419 5750 42422 5776
rect 42448 5770 42451 5776
rect 42512 5771 42541 5774
rect 42512 5770 42518 5771
rect 42448 5756 42518 5770
rect 42448 5750 42451 5756
rect 42512 5754 42518 5756
rect 42535 5754 42541 5771
rect 42512 5751 42541 5754
rect 42834 5771 42863 5774
rect 42834 5754 42840 5771
rect 42857 5770 42863 5771
rect 43201 5770 43204 5776
rect 42857 5756 43204 5770
rect 42857 5754 42863 5756
rect 42834 5751 42863 5754
rect 43201 5750 43204 5756
rect 43230 5750 43233 5776
rect 50746 5771 50775 5774
rect 50746 5754 50752 5771
rect 50769 5770 50775 5771
rect 50929 5770 50932 5776
rect 50769 5756 50932 5770
rect 50769 5754 50775 5756
rect 50746 5751 50775 5754
rect 50929 5750 50932 5756
rect 50958 5750 50961 5776
rect 51482 5771 51511 5774
rect 51482 5754 51488 5771
rect 51505 5770 51511 5771
rect 52033 5770 52036 5776
rect 51505 5756 52036 5770
rect 51505 5754 51511 5756
rect 51482 5751 51511 5754
rect 52033 5750 52036 5756
rect 52062 5750 52065 5776
rect 57001 5750 57004 5776
rect 57030 5770 57033 5776
rect 57324 5771 57353 5774
rect 57324 5770 57330 5771
rect 57030 5756 57330 5770
rect 57030 5750 57033 5756
rect 57324 5754 57330 5756
rect 57347 5754 57353 5771
rect 65925 5770 65928 5776
rect 65905 5756 65928 5770
rect 57324 5751 57353 5754
rect 65925 5750 65928 5756
rect 65954 5750 65957 5776
rect 73653 5750 73656 5776
rect 73682 5770 73685 5776
rect 75034 5771 75063 5774
rect 75034 5770 75040 5771
rect 73682 5756 75040 5770
rect 73682 5750 73685 5756
rect 75034 5754 75040 5756
rect 75057 5770 75063 5771
rect 75861 5770 75864 5776
rect 75057 5756 75864 5770
rect 75057 5754 75063 5756
rect 75034 5751 75063 5754
rect 75861 5750 75864 5756
rect 75890 5750 75893 5776
rect 89348 5770 89362 5824
rect 89662 5822 89668 5824
rect 89685 5822 89691 5839
rect 89992 5838 90006 5853
rect 90029 5852 90032 5878
rect 90058 5872 90061 5878
rect 90305 5872 90308 5878
rect 90058 5858 90308 5872
rect 90058 5852 90061 5858
rect 90305 5852 90308 5858
rect 90334 5852 90337 5878
rect 90397 5838 90400 5844
rect 89992 5824 90400 5838
rect 89662 5819 89691 5822
rect 90397 5818 90400 5824
rect 90426 5838 90429 5844
rect 90765 5838 90768 5844
rect 90426 5824 90768 5838
rect 90426 5818 90429 5824
rect 90765 5818 90768 5824
rect 90794 5818 90797 5844
rect 94776 5838 94790 5886
rect 94813 5852 94816 5878
rect 94842 5872 94845 5878
rect 95044 5873 95073 5876
rect 94842 5858 94864 5872
rect 94842 5852 94845 5858
rect 95044 5856 95050 5873
rect 95067 5872 95073 5873
rect 95366 5873 95395 5876
rect 95366 5872 95372 5873
rect 95067 5858 95372 5872
rect 95067 5856 95073 5858
rect 95044 5853 95073 5856
rect 95366 5856 95372 5858
rect 95389 5872 95395 5873
rect 95411 5872 95414 5878
rect 95389 5858 95414 5872
rect 95389 5856 95395 5858
rect 95366 5853 95395 5856
rect 95052 5838 95066 5853
rect 95411 5852 95414 5858
rect 95440 5852 95443 5878
rect 95917 5872 95920 5878
rect 95897 5858 95920 5872
rect 95917 5852 95920 5858
rect 95946 5852 95949 5878
rect 97030 5876 97044 5926
rect 97205 5920 97208 5926
rect 97234 5920 97237 5946
rect 97343 5920 97346 5946
rect 97372 5940 97375 5946
rect 98126 5941 98155 5944
rect 98126 5940 98132 5941
rect 97372 5926 98132 5940
rect 97372 5920 97375 5926
rect 98126 5924 98132 5926
rect 98149 5924 98155 5941
rect 101437 5940 101440 5946
rect 101417 5926 101440 5940
rect 98126 5921 98155 5924
rect 101437 5920 101440 5926
rect 101466 5920 101469 5946
rect 102036 5941 102065 5944
rect 102036 5924 102042 5941
rect 102059 5940 102065 5941
rect 102265 5940 102268 5946
rect 102059 5926 102268 5940
rect 102059 5924 102065 5926
rect 102036 5921 102065 5924
rect 102265 5920 102268 5926
rect 102294 5920 102297 5946
rect 102588 5941 102617 5944
rect 102588 5924 102594 5941
rect 102611 5940 102617 5941
rect 103277 5940 103280 5946
rect 102611 5926 103280 5940
rect 102611 5924 102617 5926
rect 102588 5921 102617 5924
rect 103277 5920 103280 5926
rect 103306 5920 103309 5946
rect 113903 5920 113906 5946
rect 113932 5940 113935 5946
rect 114134 5941 114163 5944
rect 114134 5940 114140 5941
rect 113932 5926 114140 5940
rect 113932 5920 113935 5926
rect 114134 5924 114140 5926
rect 114157 5940 114163 5941
rect 114409 5940 114412 5946
rect 114157 5926 114412 5940
rect 114157 5924 114163 5926
rect 114134 5921 114163 5924
rect 114409 5920 114412 5926
rect 114438 5940 114441 5946
rect 114732 5941 114761 5944
rect 114438 5926 114547 5940
rect 114438 5920 114441 5926
rect 98401 5906 98404 5912
rect 97773 5892 98404 5906
rect 98401 5886 98404 5892
rect 98430 5886 98433 5912
rect 101162 5907 101191 5910
rect 101162 5890 101168 5907
rect 101185 5906 101191 5907
rect 101575 5906 101578 5912
rect 101185 5892 101578 5906
rect 101185 5890 101191 5892
rect 101162 5887 101191 5890
rect 101575 5886 101578 5892
rect 101604 5886 101607 5912
rect 101990 5907 102019 5910
rect 101990 5890 101996 5907
rect 102013 5906 102019 5907
rect 102634 5907 102663 5910
rect 102634 5906 102640 5907
rect 102013 5892 102640 5906
rect 102013 5890 102019 5892
rect 101990 5887 102019 5890
rect 102634 5890 102640 5892
rect 102657 5906 102663 5907
rect 102771 5906 102774 5912
rect 102657 5892 102774 5906
rect 102657 5890 102663 5892
rect 102634 5887 102663 5890
rect 102771 5886 102774 5892
rect 102800 5886 102803 5912
rect 113857 5886 113860 5912
rect 113886 5906 113889 5912
rect 114180 5907 114209 5910
rect 114180 5906 114186 5907
rect 113886 5892 114186 5906
rect 113886 5886 113889 5892
rect 114180 5890 114186 5892
rect 114203 5890 114209 5907
rect 114533 5906 114547 5926
rect 114732 5924 114738 5941
rect 114755 5940 114761 5941
rect 114961 5940 114964 5946
rect 114755 5926 114964 5940
rect 114755 5924 114761 5926
rect 114732 5921 114761 5924
rect 114961 5920 114964 5926
rect 114990 5920 114993 5946
rect 115191 5940 115194 5946
rect 115171 5926 115194 5940
rect 115191 5920 115194 5926
rect 115220 5920 115223 5946
rect 115513 5920 115516 5946
rect 115542 5940 115545 5946
rect 115790 5941 115819 5944
rect 115790 5940 115796 5941
rect 115542 5926 115796 5940
rect 115542 5920 115545 5926
rect 115790 5924 115796 5926
rect 115813 5924 115819 5941
rect 115790 5921 115819 5924
rect 115835 5920 115838 5946
rect 115864 5940 115867 5946
rect 119378 5941 119407 5944
rect 119378 5940 119384 5941
rect 115864 5926 119384 5940
rect 115864 5920 115867 5926
rect 119378 5924 119384 5926
rect 119401 5924 119407 5941
rect 120159 5940 120162 5946
rect 120139 5926 120162 5940
rect 119378 5921 119407 5924
rect 120159 5920 120162 5926
rect 120188 5920 120191 5946
rect 120527 5940 120530 5946
rect 120507 5926 120530 5940
rect 120527 5920 120530 5926
rect 120556 5920 120559 5946
rect 120895 5940 120898 5946
rect 120875 5926 120898 5940
rect 120895 5920 120898 5926
rect 120924 5920 120927 5946
rect 125910 5941 125939 5944
rect 125910 5924 125916 5941
rect 125933 5940 125939 5941
rect 126461 5940 126464 5946
rect 125933 5926 126464 5940
rect 125933 5924 125939 5926
rect 125910 5921 125939 5924
rect 126461 5920 126464 5926
rect 126490 5920 126493 5946
rect 127060 5941 127089 5944
rect 127060 5924 127066 5941
rect 127083 5940 127089 5941
rect 127335 5940 127338 5946
rect 127083 5926 127338 5940
rect 127083 5924 127089 5926
rect 127060 5921 127089 5924
rect 127335 5920 127338 5926
rect 127364 5920 127367 5946
rect 127381 5920 127384 5946
rect 127410 5940 127413 5946
rect 127474 5941 127503 5944
rect 127474 5940 127480 5941
rect 127410 5926 127480 5940
rect 127410 5920 127413 5926
rect 127474 5924 127480 5926
rect 127497 5924 127503 5941
rect 127474 5921 127503 5924
rect 127519 5920 127522 5946
rect 127548 5940 127551 5946
rect 127796 5941 127825 5944
rect 127796 5940 127802 5941
rect 127548 5926 127802 5940
rect 127548 5920 127551 5926
rect 127796 5924 127802 5926
rect 127819 5924 127825 5941
rect 127796 5921 127825 5924
rect 132488 5941 132517 5944
rect 132488 5924 132494 5941
rect 132511 5940 132517 5941
rect 133407 5940 133410 5946
rect 132511 5926 133410 5940
rect 132511 5924 132517 5926
rect 132488 5921 132517 5924
rect 133407 5920 133410 5926
rect 133436 5920 133439 5946
rect 133684 5941 133713 5944
rect 133684 5924 133690 5941
rect 133707 5940 133713 5941
rect 134098 5941 134127 5944
rect 133707 5926 133867 5940
rect 133707 5924 133713 5926
rect 133684 5921 133713 5924
rect 114778 5907 114807 5910
rect 114778 5906 114784 5907
rect 114533 5892 114784 5906
rect 114180 5887 114209 5890
rect 114778 5890 114784 5892
rect 114801 5890 114807 5907
rect 114778 5887 114807 5890
rect 97022 5873 97051 5876
rect 97022 5856 97028 5873
rect 97045 5856 97051 5873
rect 97022 5853 97051 5856
rect 98218 5873 98247 5876
rect 98218 5856 98224 5873
rect 98241 5872 98247 5873
rect 98953 5872 98956 5878
rect 98241 5858 98956 5872
rect 98241 5856 98247 5858
rect 98218 5853 98247 5856
rect 98953 5852 98956 5858
rect 98982 5852 98985 5878
rect 100517 5852 100520 5878
rect 100546 5872 100549 5878
rect 101116 5873 101145 5876
rect 101116 5872 101122 5873
rect 100546 5858 101122 5872
rect 100546 5852 100549 5858
rect 101116 5856 101122 5858
rect 101139 5856 101145 5873
rect 101529 5872 101532 5878
rect 101509 5858 101532 5872
rect 101116 5853 101145 5856
rect 101529 5852 101532 5858
rect 101558 5852 101561 5878
rect 103185 5872 103188 5878
rect 101584 5858 103188 5872
rect 96055 5838 96058 5844
rect 94776 5824 95066 5838
rect 96035 5824 96058 5838
rect 96055 5818 96058 5824
rect 96084 5818 96087 5844
rect 97159 5838 97162 5844
rect 97139 5824 97162 5838
rect 97159 5818 97162 5824
rect 97188 5818 97191 5844
rect 97205 5818 97208 5844
rect 97234 5838 97237 5844
rect 97896 5839 97925 5842
rect 97234 5824 97688 5838
rect 97234 5818 97237 5824
rect 89386 5805 89415 5808
rect 89386 5788 89392 5805
rect 89409 5804 89415 5805
rect 90167 5804 90170 5810
rect 89409 5790 90170 5804
rect 89409 5788 89415 5790
rect 89386 5785 89415 5788
rect 90167 5784 90170 5790
rect 90196 5784 90199 5810
rect 95090 5805 95119 5808
rect 95090 5788 95096 5805
rect 95113 5804 95119 5805
rect 97674 5804 97688 5824
rect 97896 5822 97902 5839
rect 97919 5838 97925 5839
rect 98677 5838 98680 5844
rect 97919 5824 98680 5838
rect 97919 5822 97925 5824
rect 97896 5819 97925 5822
rect 98677 5818 98680 5824
rect 98706 5838 98709 5844
rect 100655 5838 100658 5844
rect 98706 5824 100658 5838
rect 98706 5818 98709 5824
rect 100655 5818 100658 5824
rect 100684 5818 100687 5844
rect 101437 5818 101440 5844
rect 101466 5838 101469 5844
rect 101584 5838 101598 5858
rect 103185 5852 103188 5858
rect 103214 5852 103217 5878
rect 114188 5872 114202 5887
rect 115421 5886 115424 5912
rect 115450 5906 115453 5912
rect 119332 5907 119361 5910
rect 115450 5892 115536 5906
rect 115450 5886 115453 5892
rect 114685 5872 114688 5878
rect 114188 5858 114688 5872
rect 114685 5852 114688 5858
rect 114714 5852 114717 5878
rect 115522 5876 115536 5892
rect 119332 5890 119338 5907
rect 119355 5906 119361 5907
rect 120067 5906 120070 5912
rect 119355 5892 120070 5906
rect 119355 5890 119361 5892
rect 119332 5887 119361 5890
rect 120067 5886 120070 5892
rect 120096 5886 120099 5912
rect 120757 5906 120760 5912
rect 120122 5892 120760 5906
rect 115146 5873 115175 5876
rect 115146 5856 115152 5873
rect 115169 5872 115175 5873
rect 115468 5873 115497 5876
rect 115468 5872 115474 5873
rect 115169 5858 115474 5872
rect 115169 5856 115175 5858
rect 115146 5853 115175 5856
rect 115468 5856 115474 5858
rect 115491 5856 115497 5873
rect 115468 5853 115497 5856
rect 115514 5873 115543 5876
rect 115514 5856 115520 5873
rect 115537 5856 115543 5873
rect 115514 5853 115543 5856
rect 101466 5824 101598 5838
rect 101466 5818 101469 5824
rect 101759 5818 101762 5844
rect 101788 5838 101791 5844
rect 102128 5839 102157 5842
rect 102128 5838 102134 5839
rect 101788 5824 102134 5838
rect 101788 5818 101791 5824
rect 102128 5822 102134 5824
rect 102151 5838 102157 5839
rect 102726 5839 102755 5842
rect 102726 5838 102732 5839
rect 102151 5824 102732 5838
rect 102151 5822 102157 5824
rect 102128 5819 102157 5822
rect 102726 5822 102732 5824
rect 102749 5838 102755 5839
rect 103921 5838 103924 5844
rect 102749 5824 103924 5838
rect 102749 5822 102755 5824
rect 102726 5819 102755 5822
rect 103921 5818 103924 5824
rect 103950 5818 103953 5844
rect 113627 5818 113630 5844
rect 113656 5838 113659 5844
rect 114226 5839 114255 5842
rect 114226 5838 114232 5839
rect 113656 5824 114232 5838
rect 113656 5818 113659 5824
rect 114226 5822 114232 5824
rect 114249 5838 114255 5839
rect 114870 5839 114899 5842
rect 114870 5838 114876 5839
rect 114249 5824 114876 5838
rect 114249 5822 114255 5824
rect 114226 5819 114255 5822
rect 114870 5822 114876 5824
rect 114893 5838 114899 5839
rect 114893 5824 115444 5838
rect 114893 5822 114899 5824
rect 114870 5819 114899 5822
rect 98723 5804 98726 5810
rect 95113 5790 95986 5804
rect 97674 5790 98726 5804
rect 95113 5788 95119 5790
rect 95090 5785 95119 5788
rect 90259 5770 90262 5776
rect 89348 5756 90262 5770
rect 90259 5750 90262 5756
rect 90288 5750 90291 5776
rect 94721 5770 94724 5776
rect 94701 5756 94724 5770
rect 94721 5750 94724 5756
rect 94750 5750 94753 5776
rect 95972 5770 95986 5790
rect 98723 5784 98726 5790
rect 98752 5784 98755 5810
rect 101713 5784 101716 5810
rect 101742 5804 101745 5810
rect 102449 5804 102452 5810
rect 101742 5790 102452 5804
rect 101742 5784 101745 5790
rect 102449 5784 102452 5790
rect 102478 5784 102481 5810
rect 113950 5805 113979 5808
rect 113950 5788 113956 5805
rect 113973 5804 113979 5805
rect 115145 5804 115148 5810
rect 113973 5790 115148 5804
rect 113973 5788 113979 5790
rect 113950 5785 113979 5788
rect 115145 5784 115148 5790
rect 115174 5784 115177 5810
rect 96653 5770 96656 5776
rect 95972 5756 96656 5770
rect 96653 5750 96656 5756
rect 96682 5750 96685 5776
rect 96745 5750 96748 5776
rect 96774 5770 96777 5776
rect 96792 5771 96821 5774
rect 96792 5770 96798 5771
rect 96774 5756 96798 5770
rect 96774 5750 96777 5756
rect 96792 5754 96798 5756
rect 96815 5770 96821 5771
rect 97895 5770 97898 5776
rect 96815 5756 97898 5770
rect 96815 5754 96821 5756
rect 96792 5751 96821 5754
rect 97895 5750 97898 5756
rect 97924 5750 97927 5776
rect 97941 5750 97944 5776
rect 97970 5770 97973 5776
rect 98493 5770 98496 5776
rect 97970 5756 98496 5770
rect 97970 5750 97973 5756
rect 98493 5750 98496 5756
rect 98522 5750 98525 5776
rect 100747 5750 100750 5776
rect 100776 5770 100779 5776
rect 101806 5771 101835 5774
rect 101806 5770 101812 5771
rect 100776 5756 101812 5770
rect 100776 5750 100779 5756
rect 101806 5754 101812 5756
rect 101829 5754 101835 5771
rect 102403 5770 102406 5776
rect 102383 5756 102406 5770
rect 101806 5751 101835 5754
rect 102403 5750 102406 5756
rect 102432 5750 102435 5776
rect 114548 5771 114577 5774
rect 114548 5754 114554 5771
rect 114571 5770 114577 5771
rect 114685 5770 114688 5776
rect 114571 5756 114688 5770
rect 114571 5754 114577 5756
rect 114548 5751 114577 5754
rect 114685 5750 114688 5756
rect 114714 5750 114717 5776
rect 115430 5770 115444 5824
rect 115476 5804 115490 5853
rect 115605 5852 115608 5878
rect 115634 5872 115637 5878
rect 120122 5876 120136 5892
rect 120757 5886 120760 5892
rect 120786 5886 120789 5912
rect 122413 5906 122416 5912
rect 121318 5892 122416 5906
rect 115882 5873 115911 5876
rect 115882 5872 115888 5873
rect 115634 5858 115888 5872
rect 115634 5852 115637 5858
rect 115882 5856 115888 5858
rect 115905 5856 115911 5873
rect 115882 5853 115911 5856
rect 120114 5873 120143 5876
rect 120114 5856 120120 5873
rect 120137 5856 120143 5873
rect 120620 5873 120649 5876
rect 120620 5872 120626 5873
rect 120114 5853 120143 5856
rect 120306 5858 120626 5872
rect 119653 5818 119656 5844
rect 119682 5838 119685 5844
rect 119975 5838 119978 5844
rect 119682 5824 119978 5838
rect 119682 5818 119685 5824
rect 119975 5818 119978 5824
rect 120004 5838 120007 5844
rect 120206 5839 120235 5842
rect 120206 5838 120212 5839
rect 120004 5824 120212 5838
rect 120004 5818 120007 5824
rect 120206 5822 120212 5824
rect 120229 5822 120235 5839
rect 120206 5819 120235 5822
rect 116065 5804 116068 5810
rect 115476 5790 116068 5804
rect 116065 5784 116068 5790
rect 116094 5784 116097 5810
rect 119930 5805 119959 5808
rect 119930 5788 119936 5805
rect 119953 5804 119959 5805
rect 120306 5804 120320 5858
rect 120620 5856 120626 5858
rect 120643 5856 120649 5873
rect 120620 5853 120649 5856
rect 120850 5873 120879 5876
rect 120850 5856 120856 5873
rect 120873 5856 120879 5873
rect 121263 5872 121266 5878
rect 121243 5858 121266 5872
rect 120850 5853 120879 5856
rect 120858 5838 120872 5853
rect 121263 5852 121266 5858
rect 121292 5852 121295 5878
rect 120987 5838 120990 5844
rect 120858 5824 120990 5838
rect 120987 5818 120990 5824
rect 121016 5838 121019 5844
rect 121318 5838 121332 5892
rect 122413 5886 122416 5892
rect 122442 5886 122445 5912
rect 127014 5907 127043 5910
rect 127014 5890 127020 5907
rect 127037 5906 127043 5907
rect 127151 5906 127154 5912
rect 127037 5892 127154 5906
rect 127037 5890 127043 5892
rect 127014 5887 127043 5890
rect 127151 5886 127154 5892
rect 127180 5886 127183 5912
rect 132212 5907 132241 5910
rect 132212 5890 132218 5907
rect 132235 5906 132241 5907
rect 133853 5906 133867 5926
rect 134098 5924 134104 5941
rect 134121 5940 134127 5941
rect 135339 5940 135342 5946
rect 134121 5926 135342 5940
rect 134121 5924 134127 5926
rect 134098 5921 134127 5924
rect 135339 5920 135342 5926
rect 135368 5920 135371 5946
rect 135385 5920 135388 5946
rect 135414 5940 135417 5946
rect 135708 5941 135737 5944
rect 135708 5940 135714 5941
rect 135414 5926 135714 5940
rect 135414 5920 135417 5926
rect 135708 5924 135714 5926
rect 135731 5924 135737 5941
rect 135708 5921 135737 5924
rect 134143 5906 134146 5912
rect 132235 5892 133193 5906
rect 133853 5892 134146 5906
rect 132235 5890 132241 5892
rect 132212 5887 132241 5890
rect 134143 5886 134146 5892
rect 134172 5886 134175 5912
rect 134925 5886 134928 5912
rect 134954 5886 134957 5912
rect 126001 5872 126004 5878
rect 125981 5858 126004 5872
rect 126001 5852 126004 5858
rect 126030 5852 126033 5878
rect 126186 5873 126215 5876
rect 126186 5856 126192 5873
rect 126209 5872 126215 5873
rect 126369 5872 126372 5878
rect 126209 5858 126372 5872
rect 126209 5856 126215 5858
rect 126186 5853 126215 5856
rect 126369 5852 126372 5858
rect 126398 5852 126401 5878
rect 126507 5852 126510 5878
rect 126536 5872 126539 5878
rect 127428 5873 127457 5876
rect 127428 5872 127434 5873
rect 126536 5858 127434 5872
rect 126536 5852 126539 5858
rect 127428 5856 127434 5858
rect 127451 5872 127457 5873
rect 127750 5873 127779 5876
rect 127750 5872 127756 5873
rect 127451 5858 127756 5872
rect 127451 5856 127457 5858
rect 127428 5853 127457 5856
rect 127750 5856 127756 5858
rect 127773 5872 127779 5873
rect 128117 5872 128120 5878
rect 127773 5858 128120 5872
rect 127773 5856 127779 5858
rect 127750 5853 127779 5856
rect 128117 5852 128120 5858
rect 128146 5872 128149 5878
rect 128623 5872 128626 5878
rect 128146 5858 128626 5872
rect 128146 5852 128149 5858
rect 128623 5852 128626 5858
rect 128652 5852 128655 5878
rect 132165 5872 132168 5878
rect 132145 5858 132168 5872
rect 132165 5852 132168 5858
rect 132194 5852 132197 5878
rect 132579 5872 132582 5878
rect 132559 5858 132582 5872
rect 132579 5852 132582 5858
rect 132608 5852 132611 5878
rect 132625 5852 132628 5878
rect 132654 5872 132657 5878
rect 132810 5873 132839 5876
rect 132810 5872 132816 5873
rect 132654 5858 132816 5872
rect 132654 5852 132657 5858
rect 132810 5856 132816 5858
rect 132833 5856 132839 5873
rect 134235 5872 134238 5878
rect 132810 5853 132839 5856
rect 134152 5858 134238 5872
rect 121016 5824 121332 5838
rect 121016 5818 121019 5824
rect 121355 5818 121358 5844
rect 121384 5838 121387 5844
rect 122275 5838 122278 5844
rect 121384 5824 122278 5838
rect 121384 5818 121387 5824
rect 122275 5818 122278 5824
rect 122304 5818 122307 5844
rect 126047 5818 126050 5844
rect 126076 5838 126079 5844
rect 127106 5839 127135 5842
rect 127106 5838 127112 5839
rect 126076 5824 127112 5838
rect 126076 5818 126079 5824
rect 127106 5822 127112 5824
rect 127129 5838 127135 5839
rect 127795 5838 127798 5844
rect 127129 5824 127798 5838
rect 127129 5822 127135 5824
rect 127106 5819 127135 5822
rect 127795 5818 127798 5824
rect 127824 5838 127827 5844
rect 128209 5838 128212 5844
rect 127824 5824 128212 5838
rect 127824 5818 127827 5824
rect 128209 5818 128212 5824
rect 128238 5818 128241 5844
rect 131981 5818 131984 5844
rect 132010 5838 132013 5844
rect 134152 5842 134166 5858
rect 134235 5852 134238 5858
rect 134264 5852 134267 5878
rect 134557 5872 134560 5878
rect 134537 5858 134560 5872
rect 134557 5852 134560 5858
rect 134586 5852 134589 5878
rect 135661 5872 135664 5878
rect 135641 5858 135664 5872
rect 135661 5852 135664 5858
rect 135690 5852 135693 5878
rect 132948 5839 132977 5842
rect 132948 5838 132954 5839
rect 132010 5824 132954 5838
rect 132010 5818 132013 5824
rect 132948 5822 132954 5824
rect 132971 5822 132977 5839
rect 132948 5819 132977 5822
rect 134144 5839 134173 5842
rect 134144 5822 134150 5839
rect 134167 5822 134173 5839
rect 134144 5819 134173 5822
rect 134190 5839 134219 5842
rect 134190 5822 134196 5839
rect 134213 5822 134219 5839
rect 134190 5819 134219 5822
rect 119953 5790 120320 5804
rect 120352 5790 124207 5804
rect 119953 5788 119959 5790
rect 119930 5785 119959 5788
rect 115835 5770 115838 5776
rect 115430 5756 115838 5770
rect 115835 5750 115838 5756
rect 115864 5750 115867 5776
rect 119699 5750 119702 5776
rect 119728 5770 119731 5776
rect 120352 5770 120366 5790
rect 119728 5756 120366 5770
rect 119728 5750 119731 5756
rect 120619 5750 120622 5776
rect 120648 5770 120651 5776
rect 121172 5771 121201 5774
rect 121172 5770 121178 5771
rect 120648 5756 121178 5770
rect 120648 5750 120651 5756
rect 121172 5754 121178 5756
rect 121195 5754 121201 5771
rect 124193 5770 124207 5790
rect 125817 5784 125820 5810
rect 125846 5804 125849 5810
rect 126462 5805 126491 5808
rect 126462 5804 126468 5805
rect 125846 5790 126468 5804
rect 125846 5784 125849 5790
rect 126462 5788 126468 5790
rect 126485 5804 126491 5805
rect 126485 5790 130417 5804
rect 126485 5788 126491 5790
rect 126462 5785 126491 5788
rect 124529 5770 124532 5776
rect 124193 5756 124532 5770
rect 121172 5751 121201 5754
rect 124529 5750 124532 5756
rect 124558 5750 124561 5776
rect 126645 5750 126648 5776
rect 126674 5770 126677 5776
rect 126830 5771 126859 5774
rect 126830 5770 126836 5771
rect 126674 5756 126836 5770
rect 126674 5750 126677 5756
rect 126830 5754 126836 5756
rect 126853 5754 126859 5771
rect 130403 5770 130417 5790
rect 134005 5784 134008 5810
rect 134034 5804 134037 5810
rect 134198 5804 134212 5819
rect 134034 5790 134212 5804
rect 134034 5784 134037 5790
rect 130877 5770 130880 5776
rect 130403 5756 130880 5770
rect 126830 5751 126859 5754
rect 130877 5750 130880 5756
rect 130906 5750 130909 5776
rect 131337 5750 131340 5776
rect 131366 5770 131369 5776
rect 133131 5770 133134 5776
rect 131366 5756 133134 5770
rect 131366 5750 131369 5756
rect 133131 5750 133134 5756
rect 133160 5750 133163 5776
rect 133177 5750 133180 5776
rect 133206 5770 133209 5776
rect 133914 5771 133943 5774
rect 133914 5770 133920 5771
rect 133206 5756 133920 5770
rect 133206 5750 133209 5756
rect 133914 5754 133920 5756
rect 133937 5754 133943 5771
rect 134244 5770 134258 5852
rect 134695 5838 134698 5844
rect 134675 5824 134698 5838
rect 134695 5818 134698 5824
rect 134724 5818 134727 5844
rect 134971 5818 134974 5844
rect 135000 5838 135003 5844
rect 135432 5839 135461 5842
rect 135432 5838 135438 5839
rect 135000 5824 135438 5838
rect 135000 5818 135003 5824
rect 135432 5822 135438 5824
rect 135455 5838 135461 5839
rect 136581 5838 136584 5844
rect 135455 5824 136584 5838
rect 135455 5822 135461 5824
rect 135432 5819 135461 5822
rect 136581 5818 136584 5824
rect 136610 5818 136613 5844
rect 137547 5770 137550 5776
rect 134244 5756 137550 5770
rect 133914 5751 133943 5754
rect 137547 5750 137550 5756
rect 137576 5750 137579 5776
rect 552 5725 152904 5736
rect 552 5699 19524 5725
rect 19550 5699 19556 5725
rect 19582 5699 19588 5725
rect 19614 5699 19620 5725
rect 19646 5699 19652 5725
rect 19678 5699 57623 5725
rect 57649 5699 57655 5725
rect 57681 5699 57687 5725
rect 57713 5699 57719 5725
rect 57745 5699 57751 5725
rect 57777 5699 95722 5725
rect 95748 5699 95754 5725
rect 95780 5699 95786 5725
rect 95812 5699 95818 5725
rect 95844 5699 95850 5725
rect 95876 5699 133821 5725
rect 133847 5699 133853 5725
rect 133879 5699 133885 5725
rect 133911 5699 133917 5725
rect 133943 5699 133949 5725
rect 133975 5699 152904 5725
rect 552 5688 152904 5699
rect 14406 5669 14435 5672
rect 14406 5652 14412 5669
rect 14429 5668 14435 5669
rect 14957 5668 14960 5674
rect 14429 5654 14960 5668
rect 14429 5652 14435 5654
rect 14406 5649 14435 5652
rect 14957 5648 14960 5654
rect 14986 5648 14989 5674
rect 15003 5648 15006 5674
rect 15032 5668 15035 5674
rect 15032 5654 15877 5668
rect 15032 5648 15035 5654
rect 14451 5614 14454 5640
rect 14480 5634 14483 5640
rect 15863 5634 15877 5654
rect 16199 5648 16202 5674
rect 16228 5668 16231 5674
rect 16659 5668 16662 5674
rect 16228 5654 16662 5668
rect 16228 5648 16231 5654
rect 16659 5648 16662 5654
rect 16688 5648 16691 5674
rect 16797 5668 16800 5674
rect 16777 5654 16800 5668
rect 16797 5648 16800 5654
rect 16826 5648 16829 5674
rect 20156 5669 20185 5672
rect 20156 5652 20162 5669
rect 20179 5668 20185 5669
rect 20201 5668 20204 5674
rect 20179 5654 20204 5668
rect 20179 5652 20185 5654
rect 20156 5649 20185 5652
rect 20201 5648 20204 5654
rect 20230 5648 20233 5674
rect 20523 5668 20526 5674
rect 20503 5654 20526 5668
rect 20523 5648 20526 5654
rect 20552 5648 20555 5674
rect 20799 5668 20802 5674
rect 20779 5654 20802 5668
rect 20799 5648 20802 5654
rect 20828 5648 20831 5674
rect 27515 5648 27518 5674
rect 27544 5668 27547 5674
rect 27654 5669 27683 5672
rect 27654 5668 27660 5669
rect 27544 5654 27660 5668
rect 27544 5648 27547 5654
rect 27654 5652 27660 5654
rect 27677 5652 27683 5669
rect 27654 5649 27683 5652
rect 28114 5669 28143 5672
rect 28114 5652 28120 5669
rect 28137 5668 28143 5669
rect 28849 5668 28852 5674
rect 28137 5654 28852 5668
rect 28137 5652 28143 5654
rect 28114 5649 28143 5652
rect 28849 5648 28852 5654
rect 28878 5648 28881 5674
rect 38187 5648 38190 5674
rect 38216 5668 38219 5674
rect 38234 5669 38263 5672
rect 38234 5668 38240 5669
rect 38216 5654 38240 5668
rect 38216 5648 38219 5654
rect 38234 5652 38240 5654
rect 38257 5652 38263 5669
rect 38234 5649 38263 5652
rect 39108 5669 39137 5672
rect 39108 5652 39114 5669
rect 39131 5668 39137 5669
rect 39383 5668 39386 5674
rect 39131 5654 39386 5668
rect 39131 5652 39137 5654
rect 39108 5649 39137 5652
rect 39383 5648 39386 5654
rect 39412 5648 39415 5674
rect 42235 5648 42238 5674
rect 42264 5668 42267 5674
rect 43110 5669 43139 5672
rect 43110 5668 43116 5669
rect 42264 5654 43116 5668
rect 42264 5648 42267 5654
rect 43110 5652 43116 5654
rect 43133 5652 43139 5669
rect 43110 5649 43139 5652
rect 43478 5669 43507 5672
rect 43478 5652 43484 5669
rect 43501 5668 43507 5669
rect 43569 5668 43572 5674
rect 43501 5654 43572 5668
rect 43501 5652 43507 5654
rect 43478 5649 43507 5652
rect 43569 5648 43572 5654
rect 43598 5648 43601 5674
rect 44122 5669 44151 5672
rect 44122 5652 44128 5669
rect 44145 5668 44151 5669
rect 44535 5668 44538 5674
rect 44145 5654 44538 5668
rect 44145 5652 44151 5654
rect 44122 5649 44151 5652
rect 44535 5648 44538 5654
rect 44564 5648 44567 5674
rect 51435 5668 51438 5674
rect 51415 5654 51438 5668
rect 51435 5648 51438 5654
rect 51464 5648 51467 5674
rect 57553 5648 57556 5674
rect 57582 5668 57585 5674
rect 58014 5669 58043 5672
rect 58014 5668 58020 5669
rect 57582 5654 58020 5668
rect 57582 5648 57585 5654
rect 58014 5652 58020 5654
rect 58037 5652 58043 5669
rect 58014 5649 58043 5652
rect 58566 5669 58595 5672
rect 58566 5652 58572 5669
rect 58589 5668 58595 5669
rect 58841 5668 58844 5674
rect 58589 5654 58844 5668
rect 58589 5652 58595 5654
rect 58566 5649 58595 5652
rect 58841 5648 58844 5654
rect 58870 5648 58873 5674
rect 65189 5648 65192 5674
rect 65218 5668 65221 5674
rect 65236 5669 65265 5672
rect 65236 5668 65242 5669
rect 65218 5654 65242 5668
rect 65218 5648 65221 5654
rect 65236 5652 65242 5654
rect 65259 5652 65265 5669
rect 65603 5668 65606 5674
rect 65583 5654 65606 5668
rect 65236 5649 65265 5652
rect 65603 5648 65606 5654
rect 65632 5648 65635 5674
rect 65880 5669 65909 5672
rect 65880 5652 65886 5669
rect 65903 5668 65909 5669
rect 66431 5668 66434 5674
rect 65903 5654 66434 5668
rect 65903 5652 65909 5654
rect 65880 5649 65909 5652
rect 66431 5648 66434 5654
rect 66460 5648 66463 5674
rect 74021 5668 74024 5674
rect 74001 5654 74024 5668
rect 74021 5648 74024 5654
rect 74050 5648 74053 5674
rect 75401 5668 75404 5674
rect 75381 5654 75404 5668
rect 75401 5648 75404 5654
rect 75430 5648 75433 5674
rect 78621 5648 78624 5674
rect 78650 5668 78653 5674
rect 78668 5669 78697 5672
rect 78668 5668 78674 5669
rect 78650 5654 78674 5668
rect 78650 5648 78653 5654
rect 78668 5652 78674 5654
rect 78691 5652 78697 5669
rect 78668 5649 78697 5652
rect 81014 5669 81043 5672
rect 81014 5652 81020 5669
rect 81037 5668 81043 5669
rect 81059 5668 81062 5674
rect 81037 5654 81062 5668
rect 81037 5652 81043 5654
rect 81014 5649 81043 5652
rect 81059 5648 81062 5654
rect 81088 5648 81091 5674
rect 81335 5668 81338 5674
rect 81315 5654 81338 5668
rect 81335 5648 81338 5654
rect 81364 5648 81367 5674
rect 81703 5648 81706 5674
rect 81732 5668 81735 5674
rect 81796 5669 81825 5672
rect 81796 5668 81802 5669
rect 81732 5654 81802 5668
rect 81732 5648 81735 5654
rect 81796 5652 81802 5654
rect 81819 5652 81825 5669
rect 81796 5649 81825 5652
rect 82945 5648 82948 5674
rect 82974 5668 82977 5674
rect 119699 5668 119702 5674
rect 82974 5654 119702 5668
rect 82974 5648 82977 5654
rect 119699 5648 119702 5654
rect 119728 5648 119731 5674
rect 119883 5648 119886 5674
rect 119912 5668 119915 5674
rect 119976 5669 120005 5672
rect 119976 5668 119982 5669
rect 119912 5654 119982 5668
rect 119912 5648 119915 5654
rect 119976 5652 119982 5654
rect 119999 5652 120005 5669
rect 119976 5649 120005 5652
rect 120021 5648 120024 5674
rect 120050 5668 120053 5674
rect 120436 5669 120465 5672
rect 120436 5668 120442 5669
rect 120050 5654 120442 5668
rect 120050 5648 120053 5654
rect 120436 5652 120442 5654
rect 120459 5652 120465 5669
rect 120436 5649 120465 5652
rect 120481 5648 120484 5674
rect 120510 5668 120513 5674
rect 120712 5669 120741 5672
rect 120712 5668 120718 5669
rect 120510 5654 120718 5668
rect 120510 5648 120513 5654
rect 120712 5652 120718 5654
rect 120735 5652 120741 5669
rect 120712 5649 120741 5652
rect 121033 5648 121036 5674
rect 121062 5668 121065 5674
rect 121080 5669 121109 5672
rect 121080 5668 121086 5669
rect 121062 5654 121086 5668
rect 121062 5648 121065 5654
rect 121080 5652 121086 5654
rect 121103 5652 121109 5669
rect 121080 5649 121109 5652
rect 126231 5648 126234 5674
rect 126260 5668 126263 5674
rect 126278 5669 126307 5672
rect 126278 5668 126284 5669
rect 126260 5654 126284 5668
rect 126260 5648 126263 5654
rect 126278 5652 126284 5654
rect 126301 5652 126307 5669
rect 126553 5668 126556 5674
rect 126533 5654 126556 5668
rect 126278 5649 126307 5652
rect 126553 5648 126556 5654
rect 126582 5648 126585 5674
rect 126876 5669 126905 5672
rect 126876 5652 126882 5669
rect 126899 5668 126905 5669
rect 127013 5668 127016 5674
rect 126899 5654 127016 5668
rect 126899 5652 126905 5654
rect 126876 5649 126905 5652
rect 127013 5648 127016 5654
rect 127042 5648 127045 5674
rect 132717 5648 132720 5674
rect 132746 5668 132749 5674
rect 132764 5669 132793 5672
rect 132764 5668 132770 5669
rect 132746 5654 132770 5668
rect 132746 5648 132749 5654
rect 132764 5652 132770 5654
rect 132787 5652 132793 5669
rect 132764 5649 132793 5652
rect 133131 5648 133134 5674
rect 133160 5668 133163 5674
rect 134006 5669 134035 5672
rect 133160 5654 133982 5668
rect 133160 5648 133163 5654
rect 18223 5634 18226 5640
rect 14480 5620 14888 5634
rect 15863 5620 18226 5634
rect 14480 5614 14483 5620
rect 13531 5580 13534 5606
rect 13560 5600 13563 5606
rect 14727 5600 14730 5606
rect 13560 5586 14730 5600
rect 13560 5580 13563 5586
rect 14727 5580 14730 5586
rect 14756 5580 14759 5606
rect 14773 5580 14776 5606
rect 14802 5600 14805 5606
rect 14820 5601 14849 5604
rect 14820 5600 14826 5601
rect 14802 5586 14826 5600
rect 14802 5580 14805 5586
rect 14820 5584 14826 5586
rect 14843 5584 14849 5601
rect 14874 5600 14888 5620
rect 18223 5614 18226 5620
rect 18252 5614 18255 5640
rect 20661 5614 20664 5640
rect 20690 5634 20693 5640
rect 21122 5635 21151 5638
rect 21122 5634 21128 5635
rect 20690 5620 21128 5634
rect 20690 5614 20693 5620
rect 21122 5618 21128 5620
rect 21145 5618 21151 5635
rect 21122 5615 21151 5618
rect 43385 5614 43388 5640
rect 43414 5634 43417 5640
rect 43800 5635 43829 5638
rect 43800 5634 43806 5635
rect 43414 5620 43806 5634
rect 43414 5614 43417 5620
rect 43800 5618 43806 5620
rect 43823 5618 43829 5635
rect 43800 5615 43829 5618
rect 51113 5614 51116 5640
rect 51142 5634 51145 5640
rect 51758 5635 51787 5638
rect 51758 5634 51764 5635
rect 51142 5620 51764 5634
rect 51142 5614 51145 5620
rect 51758 5618 51764 5620
rect 51781 5618 51787 5635
rect 51758 5615 51787 5618
rect 57093 5614 57096 5640
rect 57122 5634 57125 5640
rect 57692 5635 57721 5638
rect 57692 5634 57698 5635
rect 57122 5620 57698 5634
rect 57122 5614 57125 5620
rect 57692 5618 57698 5620
rect 57715 5618 57721 5635
rect 57692 5615 57721 5618
rect 73699 5614 73702 5640
rect 73728 5634 73731 5640
rect 74942 5635 74971 5638
rect 73728 5620 74366 5634
rect 73728 5614 73731 5620
rect 15693 5600 15696 5606
rect 14874 5586 15696 5600
rect 14820 5581 14849 5584
rect 15693 5580 15696 5586
rect 15722 5580 15725 5606
rect 16153 5600 16156 5606
rect 16133 5586 16156 5600
rect 16153 5580 16156 5586
rect 16182 5580 16185 5606
rect 16246 5601 16275 5604
rect 16246 5584 16252 5601
rect 16269 5600 16275 5601
rect 16291 5600 16294 5606
rect 16269 5586 16294 5600
rect 16269 5584 16275 5586
rect 16246 5581 16275 5584
rect 13807 5546 13810 5572
rect 13836 5566 13839 5572
rect 14498 5567 14527 5570
rect 14498 5566 14504 5567
rect 13836 5552 14504 5566
rect 13836 5546 13839 5552
rect 14498 5550 14504 5552
rect 14521 5550 14527 5567
rect 16107 5566 16110 5572
rect 16087 5552 16110 5566
rect 14498 5547 14527 5550
rect 16107 5546 16110 5552
rect 16136 5546 16139 5572
rect 13991 5512 13994 5538
rect 14020 5532 14023 5538
rect 14957 5532 14960 5538
rect 14020 5518 14888 5532
rect 14937 5518 14960 5532
rect 14020 5512 14023 5518
rect 14874 5498 14888 5518
rect 14957 5512 14960 5518
rect 14986 5512 14989 5538
rect 15831 5532 15834 5538
rect 15571 5518 15834 5532
rect 15831 5512 15834 5518
rect 15860 5512 15863 5538
rect 15877 5512 15880 5538
rect 15906 5532 15909 5538
rect 16254 5532 16268 5581
rect 16291 5580 16294 5586
rect 16320 5580 16323 5606
rect 22501 5600 22504 5606
rect 20900 5586 22504 5600
rect 16752 5567 16781 5570
rect 16752 5550 16758 5567
rect 16775 5566 16781 5567
rect 17349 5566 17352 5572
rect 16775 5552 17352 5566
rect 16775 5550 16781 5552
rect 16752 5547 16781 5550
rect 17349 5546 17352 5552
rect 17378 5546 17381 5572
rect 20247 5566 20250 5572
rect 20227 5552 20250 5566
rect 20247 5546 20250 5552
rect 20276 5546 20279 5572
rect 20478 5567 20507 5570
rect 20478 5550 20484 5567
rect 20501 5566 20507 5567
rect 20707 5566 20710 5572
rect 20501 5552 20710 5566
rect 20501 5550 20507 5552
rect 20478 5547 20507 5550
rect 20707 5546 20710 5552
rect 20736 5546 20739 5572
rect 20900 5570 20914 5586
rect 22501 5580 22504 5586
rect 22530 5580 22533 5606
rect 42741 5580 42744 5606
rect 42770 5600 42773 5606
rect 44581 5600 44584 5606
rect 42770 5586 44584 5600
rect 42770 5580 42773 5586
rect 20892 5567 20921 5570
rect 20892 5550 20898 5567
rect 20915 5550 20921 5567
rect 21213 5566 21216 5572
rect 21193 5552 21216 5566
rect 20892 5547 20921 5550
rect 21213 5546 21216 5552
rect 21242 5546 21245 5572
rect 27745 5566 27748 5572
rect 27725 5552 27748 5566
rect 27745 5546 27748 5552
rect 27774 5546 27777 5572
rect 28206 5567 28235 5570
rect 28206 5550 28212 5567
rect 28229 5566 28235 5567
rect 28619 5566 28622 5572
rect 28229 5552 28622 5566
rect 28229 5550 28235 5552
rect 28206 5547 28235 5550
rect 28619 5546 28622 5552
rect 28648 5546 28651 5572
rect 37359 5546 37362 5572
rect 37388 5566 37391 5572
rect 38326 5567 38355 5570
rect 38326 5566 38332 5567
rect 37388 5552 38332 5566
rect 37388 5546 37391 5552
rect 38326 5550 38332 5552
rect 38349 5550 38355 5567
rect 39199 5566 39202 5572
rect 39179 5552 39202 5566
rect 38326 5547 38355 5550
rect 39199 5546 39202 5552
rect 39228 5546 39231 5572
rect 43201 5566 43204 5572
rect 43181 5552 43204 5566
rect 43201 5546 43204 5552
rect 43230 5546 43233 5572
rect 43440 5570 43454 5586
rect 44581 5580 44584 5586
rect 44610 5580 44613 5606
rect 51021 5580 51024 5606
rect 51050 5600 51053 5606
rect 51160 5601 51189 5604
rect 51160 5600 51166 5601
rect 51050 5586 51166 5600
rect 51050 5580 51053 5586
rect 51160 5584 51166 5586
rect 51183 5584 51189 5601
rect 51160 5581 51189 5584
rect 51297 5580 51300 5606
rect 51326 5600 51329 5606
rect 51326 5586 51757 5600
rect 51326 5580 51329 5586
rect 43432 5567 43461 5570
rect 43432 5550 43438 5567
rect 43455 5550 43461 5567
rect 43891 5566 43894 5572
rect 43871 5552 43894 5566
rect 43432 5547 43461 5550
rect 43891 5546 43894 5552
rect 43920 5546 43923 5572
rect 44213 5566 44216 5572
rect 44193 5552 44216 5566
rect 44213 5546 44216 5552
rect 44242 5546 44245 5572
rect 51068 5567 51097 5570
rect 51068 5550 51074 5567
rect 51091 5566 51097 5567
rect 51205 5566 51208 5572
rect 51091 5552 51208 5566
rect 51091 5550 51097 5552
rect 51068 5547 51097 5550
rect 51205 5546 51208 5552
rect 51234 5546 51237 5572
rect 51527 5566 51530 5572
rect 51507 5552 51530 5566
rect 51527 5546 51530 5552
rect 51556 5546 51559 5572
rect 51743 5566 51757 5586
rect 65143 5580 65146 5606
rect 65172 5600 65175 5606
rect 66293 5600 66296 5606
rect 65172 5586 66296 5600
rect 65172 5580 65175 5586
rect 51850 5567 51879 5570
rect 51850 5566 51856 5567
rect 51743 5552 51856 5566
rect 51850 5550 51856 5552
rect 51873 5550 51879 5567
rect 51850 5547 51879 5550
rect 57369 5546 57372 5572
rect 57398 5566 57401 5572
rect 57646 5567 57675 5570
rect 57646 5566 57652 5567
rect 57398 5552 57652 5566
rect 57398 5546 57401 5552
rect 57646 5550 57652 5552
rect 57669 5566 57675 5567
rect 57875 5566 57878 5572
rect 57669 5552 57878 5566
rect 57669 5550 57675 5552
rect 57646 5547 57675 5550
rect 57875 5546 57878 5552
rect 57904 5546 57907 5572
rect 57921 5546 57924 5572
rect 57950 5566 57953 5572
rect 58106 5567 58135 5570
rect 58106 5566 58112 5567
rect 57950 5552 58112 5566
rect 57950 5546 57953 5552
rect 58106 5550 58112 5552
rect 58129 5550 58135 5567
rect 58106 5547 58135 5550
rect 58658 5567 58687 5570
rect 58658 5550 58664 5567
rect 58681 5566 58687 5567
rect 59853 5566 59856 5572
rect 58681 5552 59856 5566
rect 58681 5550 58687 5552
rect 58658 5547 58687 5550
rect 59853 5546 59856 5552
rect 59882 5546 59885 5572
rect 65328 5567 65357 5570
rect 65328 5550 65334 5567
rect 65351 5566 65357 5567
rect 65465 5566 65468 5572
rect 65351 5552 65468 5566
rect 65351 5550 65357 5552
rect 65328 5547 65357 5550
rect 65465 5546 65468 5552
rect 65494 5546 65497 5572
rect 65566 5570 65580 5586
rect 66293 5580 66296 5586
rect 66322 5580 66325 5606
rect 71629 5580 71632 5606
rect 71658 5600 71661 5606
rect 71658 5586 72940 5600
rect 71658 5580 71661 5586
rect 65558 5567 65587 5570
rect 65558 5550 65564 5567
rect 65581 5550 65587 5567
rect 65558 5547 65587 5550
rect 65972 5567 66001 5570
rect 65972 5550 65978 5567
rect 65995 5566 66001 5567
rect 66569 5566 66572 5572
rect 65995 5552 66572 5566
rect 65995 5550 66001 5552
rect 65972 5547 66001 5550
rect 66569 5546 66572 5552
rect 66598 5546 66601 5572
rect 71031 5566 71034 5572
rect 70987 5552 71034 5566
rect 71031 5546 71034 5552
rect 71060 5566 71063 5572
rect 72871 5566 72874 5572
rect 71060 5552 72874 5566
rect 71060 5546 71063 5552
rect 72871 5546 72874 5552
rect 72900 5546 72903 5572
rect 72926 5566 72940 5586
rect 73745 5580 73748 5606
rect 73774 5600 73777 5606
rect 74352 5604 74366 5620
rect 74942 5618 74948 5635
rect 74965 5634 74971 5635
rect 78207 5634 78210 5640
rect 74965 5620 78210 5634
rect 74965 5618 74971 5620
rect 74942 5615 74971 5618
rect 78207 5614 78210 5620
rect 78236 5614 78239 5640
rect 82715 5614 82718 5640
rect 82744 5634 82747 5640
rect 126369 5634 126372 5640
rect 82744 5620 96078 5634
rect 82744 5614 82747 5620
rect 74252 5601 74281 5604
rect 74252 5600 74258 5601
rect 73774 5586 74258 5600
rect 73774 5580 73777 5586
rect 74252 5584 74258 5586
rect 74275 5584 74281 5601
rect 74252 5581 74281 5584
rect 74344 5601 74373 5604
rect 74344 5584 74350 5601
rect 74367 5600 74373 5601
rect 75677 5600 75680 5606
rect 74367 5586 75680 5600
rect 74367 5584 74373 5586
rect 74344 5581 74373 5584
rect 75677 5580 75680 5586
rect 75706 5580 75709 5606
rect 82669 5600 82672 5606
rect 81436 5586 82672 5600
rect 75494 5567 75523 5570
rect 72926 5552 74780 5566
rect 15906 5518 16268 5532
rect 15906 5512 15909 5518
rect 40809 5512 40812 5538
rect 40838 5532 40841 5538
rect 43937 5532 43940 5538
rect 40838 5518 43940 5532
rect 40838 5512 40841 5518
rect 43937 5512 43940 5518
rect 43966 5512 43969 5538
rect 51214 5532 51228 5546
rect 56863 5532 56866 5538
rect 51214 5518 56866 5532
rect 56863 5512 56866 5518
rect 56892 5512 56895 5538
rect 70204 5533 70233 5536
rect 70204 5516 70210 5533
rect 70227 5532 70233 5533
rect 70341 5532 70344 5538
rect 70227 5518 70344 5532
rect 70227 5516 70233 5518
rect 70204 5513 70233 5516
rect 70341 5512 70344 5518
rect 70370 5532 70373 5538
rect 74766 5532 74780 5552
rect 75494 5550 75500 5567
rect 75517 5566 75523 5567
rect 76551 5566 76554 5572
rect 75517 5552 76554 5566
rect 75517 5550 75523 5552
rect 75494 5547 75523 5550
rect 76551 5546 76554 5552
rect 76580 5546 76583 5572
rect 81105 5566 81108 5572
rect 81085 5552 81108 5566
rect 81105 5546 81108 5552
rect 81134 5546 81137 5572
rect 81436 5570 81450 5586
rect 82669 5580 82672 5586
rect 82698 5580 82701 5606
rect 88788 5601 88817 5604
rect 88788 5584 88794 5601
rect 88811 5600 88817 5601
rect 88833 5600 88836 5606
rect 88811 5586 88836 5600
rect 88811 5584 88817 5586
rect 88788 5581 88817 5584
rect 88833 5580 88836 5586
rect 88862 5580 88865 5606
rect 88971 5580 88974 5606
rect 89000 5600 89003 5606
rect 89110 5601 89139 5604
rect 89110 5600 89116 5601
rect 89000 5586 89116 5600
rect 89000 5580 89003 5586
rect 89110 5584 89116 5586
rect 89133 5584 89139 5601
rect 90397 5600 90400 5606
rect 89110 5581 89139 5584
rect 89302 5586 90400 5600
rect 81428 5567 81457 5570
rect 81428 5550 81434 5567
rect 81451 5550 81457 5567
rect 81749 5566 81752 5572
rect 81729 5552 81752 5566
rect 81428 5547 81457 5550
rect 81749 5546 81752 5552
rect 81778 5546 81781 5572
rect 88742 5567 88771 5570
rect 88742 5550 88748 5567
rect 88765 5566 88771 5567
rect 89017 5566 89020 5572
rect 88765 5552 89020 5566
rect 88765 5550 88771 5552
rect 88742 5547 88771 5550
rect 89017 5546 89020 5552
rect 89046 5566 89049 5572
rect 89064 5567 89093 5570
rect 89064 5566 89070 5567
rect 89046 5552 89070 5566
rect 89046 5546 89049 5552
rect 89064 5550 89070 5552
rect 89087 5566 89093 5567
rect 89302 5566 89316 5586
rect 90397 5580 90400 5586
rect 90426 5580 90429 5606
rect 95136 5601 95165 5604
rect 95136 5584 95142 5601
rect 95159 5600 95165 5601
rect 95595 5600 95598 5606
rect 95159 5586 95598 5600
rect 95159 5584 95165 5586
rect 95136 5581 95165 5584
rect 95595 5580 95598 5586
rect 95624 5580 95627 5606
rect 95917 5580 95920 5606
rect 95946 5600 95949 5606
rect 96010 5601 96039 5604
rect 96010 5600 96016 5601
rect 95946 5586 96016 5600
rect 95946 5580 95949 5586
rect 96010 5584 96016 5586
rect 96033 5584 96039 5601
rect 96064 5600 96078 5620
rect 96662 5620 126372 5634
rect 96662 5600 96676 5620
rect 126369 5614 126372 5620
rect 126398 5614 126401 5640
rect 126599 5614 126602 5640
rect 126628 5634 126631 5640
rect 127198 5635 127227 5638
rect 127198 5634 127204 5635
rect 126628 5620 127204 5634
rect 126628 5614 126631 5620
rect 127198 5618 127204 5620
rect 127221 5618 127227 5635
rect 127198 5615 127227 5618
rect 132579 5614 132582 5640
rect 132608 5634 132611 5640
rect 133408 5635 133437 5638
rect 133408 5634 133414 5635
rect 132608 5620 133414 5634
rect 132608 5614 132611 5620
rect 133408 5618 133414 5620
rect 133431 5618 133437 5635
rect 133968 5634 133982 5654
rect 134006 5652 134012 5669
rect 134029 5668 134035 5669
rect 134649 5668 134652 5674
rect 134029 5654 134652 5668
rect 134029 5652 134035 5654
rect 134006 5649 134035 5652
rect 134649 5648 134652 5654
rect 134678 5648 134681 5674
rect 133968 5620 134718 5634
rect 133408 5615 133437 5618
rect 96064 5586 96676 5600
rect 96010 5581 96039 5584
rect 96745 5580 96748 5606
rect 96774 5600 96777 5606
rect 96884 5601 96913 5604
rect 96884 5600 96890 5601
rect 96774 5586 96890 5600
rect 96774 5580 96777 5586
rect 96884 5584 96890 5586
rect 96907 5600 96913 5601
rect 97205 5600 97208 5606
rect 96907 5586 97208 5600
rect 96907 5584 96913 5586
rect 96884 5581 96913 5584
rect 97205 5580 97208 5586
rect 97234 5580 97237 5606
rect 97297 5580 97300 5606
rect 97326 5600 97329 5606
rect 97482 5601 97511 5604
rect 97482 5600 97488 5601
rect 97326 5586 97488 5600
rect 97326 5580 97329 5586
rect 97482 5584 97488 5586
rect 97505 5584 97511 5601
rect 98217 5600 98220 5606
rect 97482 5581 97511 5584
rect 97720 5586 98220 5600
rect 89087 5552 89316 5566
rect 89570 5567 89599 5570
rect 89087 5550 89093 5552
rect 89064 5547 89093 5550
rect 89570 5550 89576 5567
rect 89593 5566 89599 5567
rect 90213 5566 90216 5572
rect 89593 5552 90216 5566
rect 89593 5550 89599 5552
rect 89570 5547 89599 5550
rect 90213 5546 90216 5552
rect 90242 5546 90245 5572
rect 94491 5546 94494 5572
rect 94520 5566 94523 5572
rect 95090 5567 95119 5570
rect 95090 5566 95096 5567
rect 94520 5552 95096 5566
rect 94520 5546 94523 5552
rect 95090 5550 95096 5552
rect 95113 5566 95119 5567
rect 95319 5566 95322 5572
rect 95113 5552 95322 5566
rect 95113 5550 95119 5552
rect 95090 5547 95119 5550
rect 95319 5546 95322 5552
rect 95348 5546 95351 5572
rect 95411 5566 95414 5572
rect 95391 5552 95414 5566
rect 95411 5546 95414 5552
rect 95440 5546 95443 5572
rect 95458 5567 95487 5570
rect 95458 5550 95464 5567
rect 95481 5566 95487 5567
rect 95963 5566 95966 5572
rect 95481 5552 95966 5566
rect 95481 5550 95487 5552
rect 95458 5547 95487 5550
rect 95963 5546 95966 5552
rect 95992 5546 95995 5572
rect 97390 5567 97419 5570
rect 97390 5550 97396 5567
rect 97413 5566 97419 5567
rect 97435 5566 97438 5572
rect 97413 5552 97438 5566
rect 97413 5550 97419 5552
rect 97390 5547 97419 5550
rect 97435 5546 97438 5552
rect 97464 5546 97467 5572
rect 97720 5566 97734 5586
rect 98217 5580 98220 5586
rect 98246 5580 98249 5606
rect 100517 5580 100520 5606
rect 100546 5600 100549 5606
rect 101438 5601 101467 5604
rect 100546 5586 101414 5600
rect 100546 5580 100549 5586
rect 97895 5566 97898 5572
rect 97582 5552 97734 5566
rect 97875 5552 97898 5566
rect 74804 5533 74833 5536
rect 74804 5532 74810 5533
rect 70370 5518 74734 5532
rect 74766 5518 74810 5532
rect 70370 5512 70373 5518
rect 15694 5499 15723 5502
rect 15694 5498 15700 5499
rect 14874 5484 15700 5498
rect 15694 5482 15700 5484
rect 15717 5482 15723 5499
rect 15923 5498 15926 5504
rect 15903 5484 15926 5498
rect 15694 5479 15723 5482
rect 15923 5478 15926 5484
rect 15952 5478 15955 5504
rect 74206 5499 74235 5502
rect 74206 5482 74212 5499
rect 74229 5498 74235 5499
rect 74527 5498 74530 5504
rect 74229 5484 74530 5498
rect 74229 5482 74235 5484
rect 74206 5479 74235 5482
rect 74527 5478 74530 5484
rect 74556 5478 74559 5504
rect 74720 5498 74734 5518
rect 74804 5516 74810 5518
rect 74827 5516 74833 5533
rect 78024 5533 78053 5536
rect 78024 5532 78030 5533
rect 74804 5513 74833 5516
rect 74858 5518 78030 5532
rect 74757 5498 74760 5504
rect 74720 5484 74760 5498
rect 74757 5478 74760 5484
rect 74786 5498 74789 5504
rect 74858 5498 74872 5518
rect 78024 5516 78030 5518
rect 78047 5532 78053 5533
rect 78069 5532 78072 5538
rect 78047 5518 78072 5532
rect 78047 5516 78053 5518
rect 78024 5513 78053 5516
rect 78069 5512 78072 5518
rect 78098 5512 78101 5538
rect 89707 5532 89710 5538
rect 89486 5518 89710 5532
rect 89486 5502 89500 5518
rect 89707 5512 89710 5518
rect 89736 5512 89739 5538
rect 94721 5512 94724 5538
rect 94750 5532 94753 5538
rect 96148 5533 96177 5536
rect 96148 5532 96154 5533
rect 94750 5518 96154 5532
rect 94750 5512 94753 5518
rect 96148 5516 96154 5518
rect 96171 5516 96177 5533
rect 96148 5513 96177 5516
rect 96653 5512 96656 5538
rect 96682 5512 96685 5538
rect 97582 5532 97596 5552
rect 97895 5546 97898 5552
rect 97924 5546 97927 5572
rect 101162 5567 101191 5570
rect 101162 5550 101168 5567
rect 101185 5566 101191 5567
rect 101345 5566 101348 5572
rect 101185 5552 101348 5566
rect 101185 5550 101191 5552
rect 101162 5547 101191 5550
rect 101345 5546 101348 5552
rect 101374 5546 101377 5572
rect 101400 5570 101414 5586
rect 101438 5584 101444 5601
rect 101461 5600 101467 5601
rect 101667 5600 101670 5606
rect 101461 5586 101670 5600
rect 101461 5584 101467 5586
rect 101438 5581 101467 5584
rect 101667 5580 101670 5586
rect 101696 5580 101699 5606
rect 102495 5600 102498 5606
rect 101768 5586 102498 5600
rect 101392 5567 101421 5570
rect 101392 5550 101398 5567
rect 101415 5566 101421 5567
rect 101714 5567 101743 5570
rect 101714 5566 101720 5567
rect 101415 5552 101720 5566
rect 101415 5550 101421 5552
rect 101392 5547 101421 5550
rect 101714 5550 101720 5552
rect 101737 5550 101743 5567
rect 101714 5547 101743 5550
rect 97444 5518 97596 5532
rect 74786 5484 74872 5498
rect 89478 5499 89507 5502
rect 74786 5478 74789 5484
rect 89478 5482 89484 5499
rect 89501 5482 89507 5499
rect 97205 5498 97208 5504
rect 97185 5484 97208 5498
rect 89478 5479 89507 5482
rect 97205 5478 97208 5484
rect 97234 5478 97237 5504
rect 97444 5502 97458 5518
rect 97619 5512 97622 5538
rect 97648 5532 97651 5538
rect 101768 5532 101782 5586
rect 102495 5580 102498 5586
rect 102524 5580 102527 5606
rect 119009 5580 119012 5606
rect 119038 5600 119041 5606
rect 121355 5600 121358 5606
rect 119038 5586 121358 5600
rect 119038 5580 119041 5586
rect 121355 5580 121358 5586
rect 121384 5580 121387 5606
rect 132488 5601 132517 5604
rect 132488 5584 132494 5601
rect 132511 5600 132517 5601
rect 133637 5600 133640 5606
rect 132511 5586 133640 5600
rect 132511 5584 132517 5586
rect 132488 5581 132517 5584
rect 133637 5580 133640 5586
rect 133666 5580 133669 5606
rect 133730 5601 133759 5604
rect 133730 5584 133736 5601
rect 133753 5600 133759 5601
rect 134005 5600 134008 5606
rect 133753 5586 134008 5600
rect 133753 5584 133759 5586
rect 133730 5581 133759 5584
rect 134005 5580 134008 5586
rect 134034 5580 134037 5606
rect 134235 5600 134238 5606
rect 134060 5586 134238 5600
rect 97648 5518 97826 5532
rect 97648 5512 97651 5518
rect 97812 5502 97826 5518
rect 101078 5518 101782 5532
rect 101814 5552 102426 5566
rect 101078 5502 101092 5518
rect 97436 5499 97465 5502
rect 97436 5482 97442 5499
rect 97459 5482 97465 5499
rect 97436 5479 97465 5482
rect 97804 5499 97833 5502
rect 97804 5482 97810 5499
rect 97827 5482 97833 5499
rect 97804 5479 97833 5482
rect 101070 5499 101099 5502
rect 101070 5482 101076 5499
rect 101093 5482 101099 5499
rect 101070 5479 101099 5482
rect 101760 5499 101789 5502
rect 101760 5482 101766 5499
rect 101783 5498 101789 5499
rect 101814 5498 101828 5552
rect 102035 5512 102038 5538
rect 102064 5532 102067 5538
rect 102412 5532 102426 5552
rect 102449 5546 102452 5572
rect 102478 5566 102481 5572
rect 114685 5566 114688 5572
rect 102478 5552 102500 5566
rect 114665 5552 114688 5566
rect 102478 5546 102481 5552
rect 114685 5546 114688 5552
rect 114714 5546 114717 5572
rect 119930 5567 119959 5570
rect 119930 5550 119936 5567
rect 119953 5566 119959 5567
rect 120390 5567 120419 5570
rect 120390 5566 120396 5567
rect 119953 5552 120396 5566
rect 119953 5550 119959 5552
rect 119930 5547 119959 5550
rect 120390 5550 120396 5552
rect 120413 5550 120419 5567
rect 120390 5547 120419 5550
rect 102725 5532 102728 5538
rect 102064 5518 102380 5532
rect 102412 5518 102728 5532
rect 102064 5512 102067 5518
rect 102366 5502 102380 5518
rect 102725 5512 102728 5518
rect 102754 5512 102757 5538
rect 115375 5532 115378 5538
rect 114602 5518 115378 5532
rect 114602 5502 114616 5518
rect 115375 5512 115378 5518
rect 115404 5512 115407 5538
rect 120398 5532 120412 5547
rect 120435 5546 120438 5572
rect 120464 5566 120467 5572
rect 120804 5567 120833 5570
rect 120804 5566 120810 5567
rect 120464 5552 120810 5566
rect 120464 5546 120467 5552
rect 120804 5550 120810 5552
rect 120827 5550 120833 5567
rect 120804 5547 120833 5550
rect 120987 5546 120990 5572
rect 121016 5566 121019 5572
rect 121034 5567 121063 5570
rect 121034 5566 121040 5567
rect 121016 5552 121040 5566
rect 121016 5546 121019 5552
rect 121034 5550 121040 5552
rect 121057 5550 121063 5567
rect 121034 5547 121063 5550
rect 125771 5546 125774 5572
rect 125800 5566 125803 5572
rect 126232 5567 126261 5570
rect 126232 5566 126238 5567
rect 125800 5552 126238 5566
rect 125800 5546 125803 5552
rect 126232 5550 126238 5552
rect 126255 5566 126261 5567
rect 126507 5566 126510 5572
rect 126255 5552 126510 5566
rect 126255 5550 126261 5552
rect 126232 5547 126261 5550
rect 126507 5546 126510 5552
rect 126536 5546 126539 5572
rect 126645 5566 126648 5572
rect 126625 5552 126648 5566
rect 126645 5546 126648 5552
rect 126674 5546 126677 5572
rect 126968 5567 126997 5570
rect 126968 5550 126974 5567
rect 126991 5566 126997 5567
rect 127197 5566 127200 5572
rect 126991 5552 127200 5566
rect 126991 5550 126997 5552
rect 126968 5547 126997 5550
rect 127197 5546 127200 5552
rect 127226 5546 127229 5572
rect 127290 5567 127319 5570
rect 127290 5550 127296 5567
rect 127313 5566 127319 5567
rect 127335 5566 127338 5572
rect 127313 5552 127338 5566
rect 127313 5550 127319 5552
rect 127290 5547 127319 5550
rect 127335 5546 127338 5552
rect 127364 5546 127367 5572
rect 132165 5546 132168 5572
rect 132194 5566 132197 5572
rect 132441 5566 132444 5572
rect 132194 5552 132444 5566
rect 132194 5546 132197 5552
rect 132441 5546 132444 5552
rect 132470 5546 132473 5572
rect 132809 5546 132812 5572
rect 132838 5566 132841 5572
rect 132856 5567 132885 5570
rect 132856 5566 132862 5567
rect 132838 5552 132862 5566
rect 132838 5546 132841 5552
rect 132856 5550 132862 5552
rect 132879 5550 132885 5567
rect 132856 5547 132885 5550
rect 133592 5567 133621 5570
rect 133592 5550 133598 5567
rect 133615 5566 133621 5567
rect 134060 5566 134074 5586
rect 134235 5580 134238 5586
rect 134264 5580 134267 5606
rect 134282 5601 134311 5604
rect 134282 5584 134288 5601
rect 134305 5600 134311 5601
rect 134465 5600 134468 5606
rect 134305 5586 134468 5600
rect 134305 5584 134311 5586
rect 134282 5581 134311 5584
rect 134465 5580 134468 5586
rect 134494 5580 134497 5606
rect 134704 5604 134718 5620
rect 134696 5601 134725 5604
rect 134696 5584 134702 5601
rect 134719 5600 134725 5601
rect 135294 5601 135323 5604
rect 135294 5600 135300 5601
rect 134719 5586 135300 5600
rect 134719 5584 134725 5586
rect 134696 5581 134725 5584
rect 135294 5584 135300 5586
rect 135317 5600 135323 5601
rect 136121 5600 136124 5606
rect 135317 5586 136124 5600
rect 135317 5584 135323 5586
rect 135294 5581 135323 5584
rect 136121 5580 136124 5586
rect 136150 5580 136153 5606
rect 133615 5552 134074 5566
rect 134098 5567 134127 5570
rect 133615 5550 133621 5552
rect 133592 5547 133621 5550
rect 134098 5550 134104 5567
rect 134121 5566 134127 5567
rect 134833 5566 134836 5572
rect 134121 5552 134836 5566
rect 134121 5550 134127 5552
rect 134098 5547 134127 5550
rect 134833 5546 134836 5552
rect 134862 5546 134865 5572
rect 135201 5566 135204 5572
rect 135181 5552 135204 5566
rect 135201 5546 135204 5552
rect 135230 5546 135233 5572
rect 135248 5567 135277 5570
rect 135248 5550 135254 5567
rect 135271 5566 135277 5567
rect 135431 5566 135434 5572
rect 135271 5552 135434 5566
rect 135271 5550 135277 5552
rect 135248 5547 135277 5550
rect 135431 5546 135434 5552
rect 135460 5546 135463 5572
rect 120996 5532 121010 5546
rect 120398 5518 121010 5532
rect 133638 5533 133667 5536
rect 133638 5516 133644 5533
rect 133661 5532 133667 5533
rect 134143 5532 134146 5538
rect 133661 5518 134146 5532
rect 133661 5516 133667 5518
rect 133638 5513 133667 5516
rect 134143 5512 134146 5518
rect 134172 5512 134175 5538
rect 134465 5512 134468 5538
rect 134494 5532 134497 5538
rect 134604 5533 134633 5536
rect 134604 5532 134610 5533
rect 134494 5518 134610 5532
rect 134494 5512 134497 5518
rect 134604 5516 134610 5518
rect 134627 5516 134633 5533
rect 134604 5513 134633 5516
rect 134650 5533 134679 5536
rect 134650 5516 134656 5533
rect 134673 5532 134679 5533
rect 134971 5532 134974 5538
rect 134673 5518 134974 5532
rect 134673 5516 134679 5518
rect 134650 5513 134679 5516
rect 134971 5512 134974 5518
rect 135000 5512 135003 5538
rect 101783 5484 101828 5498
rect 102358 5499 102387 5502
rect 101783 5482 101789 5484
rect 101760 5479 101789 5482
rect 102358 5482 102364 5499
rect 102381 5482 102387 5499
rect 102358 5479 102387 5482
rect 114594 5499 114623 5502
rect 114594 5482 114600 5499
rect 114617 5482 114623 5499
rect 134419 5498 134422 5504
rect 134399 5484 134422 5498
rect 114594 5479 114623 5482
rect 134419 5478 134422 5484
rect 134448 5478 134451 5504
rect 135017 5498 135020 5504
rect 134997 5484 135020 5498
rect 135017 5478 135020 5484
rect 135046 5478 135049 5504
rect 552 5453 152904 5464
rect 552 5427 38574 5453
rect 38600 5427 38606 5453
rect 38632 5427 38638 5453
rect 38664 5427 38670 5453
rect 38696 5427 38702 5453
rect 38728 5427 76673 5453
rect 76699 5427 76705 5453
rect 76731 5427 76737 5453
rect 76763 5427 76769 5453
rect 76795 5427 76801 5453
rect 76827 5427 114772 5453
rect 114798 5427 114804 5453
rect 114830 5427 114836 5453
rect 114862 5427 114868 5453
rect 114894 5427 114900 5453
rect 114926 5427 152904 5453
rect 552 5416 152904 5427
rect 14820 5397 14849 5400
rect 14820 5380 14826 5397
rect 14843 5396 14849 5397
rect 14911 5396 14914 5402
rect 14843 5382 14914 5396
rect 14843 5380 14849 5382
rect 14820 5377 14849 5380
rect 14911 5376 14914 5382
rect 14940 5376 14943 5402
rect 15233 5376 15236 5402
rect 15262 5396 15265 5402
rect 15326 5397 15355 5400
rect 15326 5396 15332 5397
rect 15262 5382 15332 5396
rect 15262 5376 15265 5382
rect 15326 5380 15332 5382
rect 15349 5380 15355 5397
rect 15326 5377 15355 5380
rect 15371 5376 15374 5402
rect 15400 5396 15403 5402
rect 16062 5397 16091 5400
rect 16062 5396 16068 5397
rect 15400 5382 15422 5396
rect 15472 5382 16068 5396
rect 15400 5376 15403 5382
rect 14865 5342 14868 5368
rect 14894 5362 14897 5368
rect 14894 5348 15072 5362
rect 14894 5342 14897 5348
rect 14221 5308 14224 5334
rect 14250 5328 14253 5334
rect 14912 5329 14941 5332
rect 14912 5328 14918 5329
rect 14250 5314 14918 5328
rect 14250 5308 14253 5314
rect 14912 5312 14918 5314
rect 14935 5312 14941 5329
rect 15058 5328 15072 5348
rect 15095 5342 15098 5368
rect 15124 5362 15127 5368
rect 15472 5362 15486 5382
rect 16062 5380 16068 5382
rect 16085 5380 16091 5397
rect 16062 5377 16091 5380
rect 16337 5376 16340 5402
rect 16366 5396 16369 5402
rect 16384 5397 16413 5400
rect 16384 5396 16390 5397
rect 16366 5382 16390 5396
rect 16366 5376 16369 5382
rect 16384 5380 16390 5382
rect 16407 5380 16413 5397
rect 16384 5377 16413 5380
rect 16521 5376 16524 5402
rect 16550 5396 16553 5402
rect 16706 5397 16735 5400
rect 16706 5396 16712 5397
rect 16550 5382 16712 5396
rect 16550 5376 16553 5382
rect 16706 5380 16712 5382
rect 16729 5380 16735 5397
rect 50837 5396 50840 5402
rect 50817 5382 50840 5396
rect 16706 5377 16735 5380
rect 50837 5376 50840 5382
rect 50866 5376 50869 5402
rect 65235 5396 65238 5402
rect 65215 5382 65238 5396
rect 65235 5376 65238 5382
rect 65264 5376 65267 5402
rect 70985 5396 70988 5402
rect 70965 5382 70988 5396
rect 70985 5376 70988 5382
rect 71014 5376 71017 5402
rect 74297 5376 74300 5402
rect 74326 5396 74329 5402
rect 74436 5397 74465 5400
rect 74436 5396 74442 5397
rect 74326 5382 74442 5396
rect 74326 5376 74329 5382
rect 74436 5380 74442 5382
rect 74459 5380 74465 5397
rect 74436 5377 74465 5380
rect 74481 5376 74484 5402
rect 74510 5396 74513 5402
rect 75356 5397 75385 5400
rect 75356 5396 75362 5397
rect 74510 5382 75362 5396
rect 74510 5376 74513 5382
rect 75356 5380 75362 5382
rect 75379 5380 75385 5397
rect 75356 5377 75385 5380
rect 95549 5376 95552 5402
rect 95578 5396 95581 5402
rect 95918 5397 95947 5400
rect 95918 5396 95924 5397
rect 95578 5382 95924 5396
rect 95578 5376 95581 5382
rect 95918 5380 95924 5382
rect 95941 5380 95947 5397
rect 95918 5377 95947 5380
rect 96064 5382 96906 5396
rect 15877 5362 15880 5368
rect 15124 5348 15486 5362
rect 15518 5348 15880 5362
rect 15124 5342 15127 5348
rect 15518 5328 15532 5348
rect 15877 5342 15880 5348
rect 15906 5342 15909 5368
rect 15923 5342 15926 5368
rect 15952 5362 15955 5368
rect 70341 5362 70344 5368
rect 15952 5348 16820 5362
rect 70321 5348 70344 5362
rect 15952 5342 15955 5348
rect 16154 5329 16183 5332
rect 16154 5328 16160 5329
rect 15058 5314 15532 5328
rect 15863 5314 16160 5328
rect 14912 5309 14941 5312
rect 15426 5298 15440 5314
rect 15418 5295 15447 5298
rect 15418 5278 15424 5295
rect 15441 5278 15447 5295
rect 15418 5275 15447 5278
rect 15142 5261 15171 5264
rect 15142 5244 15148 5261
rect 15165 5260 15171 5261
rect 15863 5260 15877 5314
rect 16154 5312 16160 5314
rect 16177 5312 16183 5329
rect 16475 5328 16478 5334
rect 16455 5314 16478 5328
rect 16154 5309 16183 5312
rect 16475 5308 16478 5314
rect 16504 5308 16507 5334
rect 16806 5332 16820 5348
rect 70341 5342 70344 5348
rect 70370 5342 70373 5368
rect 75815 5362 75818 5368
rect 74536 5348 75818 5362
rect 16798 5329 16827 5332
rect 16798 5312 16804 5329
rect 16821 5312 16827 5329
rect 50929 5328 50932 5334
rect 50909 5314 50932 5328
rect 16798 5309 16827 5312
rect 50929 5308 50932 5314
rect 50958 5308 50961 5334
rect 65143 5308 65146 5334
rect 65172 5328 65175 5334
rect 74536 5332 74550 5348
rect 75815 5342 75818 5348
rect 75844 5342 75847 5368
rect 78069 5362 78072 5368
rect 78049 5348 78072 5362
rect 78069 5342 78072 5348
rect 78098 5342 78101 5368
rect 96064 5362 96078 5382
rect 93626 5348 96078 5362
rect 65190 5329 65219 5332
rect 65190 5328 65196 5329
rect 65172 5314 65196 5328
rect 65172 5308 65175 5314
rect 65190 5312 65196 5314
rect 65213 5312 65219 5329
rect 65190 5309 65219 5312
rect 74528 5329 74557 5332
rect 74528 5312 74534 5329
rect 74551 5312 74557 5329
rect 74528 5309 74557 5312
rect 75171 5308 75174 5334
rect 75200 5328 75203 5334
rect 93626 5332 93640 5348
rect 96101 5342 96104 5368
rect 96130 5362 96133 5368
rect 96130 5348 96354 5362
rect 96130 5342 96133 5348
rect 75310 5329 75339 5332
rect 75310 5328 75316 5329
rect 75200 5314 75316 5328
rect 75200 5308 75203 5314
rect 75310 5312 75316 5314
rect 75333 5312 75339 5329
rect 75310 5309 75339 5312
rect 93618 5329 93647 5332
rect 93618 5312 93624 5329
rect 93641 5312 93647 5329
rect 93618 5309 93647 5312
rect 95273 5308 95276 5334
rect 95302 5328 95305 5334
rect 95642 5329 95671 5332
rect 95642 5328 95648 5329
rect 95302 5314 95648 5328
rect 95302 5308 95305 5314
rect 95642 5312 95648 5314
rect 95665 5312 95671 5329
rect 95642 5309 95671 5312
rect 96010 5329 96039 5332
rect 96010 5312 96016 5329
rect 96033 5328 96039 5329
rect 96147 5328 96150 5334
rect 96033 5314 96150 5328
rect 96033 5312 96039 5314
rect 96010 5309 96039 5312
rect 96147 5308 96150 5314
rect 96176 5308 96179 5334
rect 96340 5332 96354 5348
rect 96607 5342 96610 5368
rect 96636 5362 96639 5368
rect 96746 5363 96775 5366
rect 96746 5362 96752 5363
rect 96636 5348 96752 5362
rect 96636 5342 96639 5348
rect 96746 5346 96752 5348
rect 96769 5346 96775 5363
rect 96892 5362 96906 5382
rect 96929 5376 96932 5402
rect 96958 5396 96961 5402
rect 97114 5397 97143 5400
rect 97114 5396 97120 5397
rect 96958 5382 97120 5396
rect 96958 5376 96961 5382
rect 97114 5380 97120 5382
rect 97137 5380 97143 5397
rect 97114 5377 97143 5380
rect 101438 5397 101467 5400
rect 101438 5380 101444 5397
rect 101461 5396 101467 5397
rect 102541 5396 102544 5402
rect 101461 5382 102544 5396
rect 101461 5380 101467 5382
rect 101438 5377 101467 5380
rect 102541 5376 102544 5382
rect 102570 5376 102573 5402
rect 126830 5397 126859 5400
rect 126830 5380 126836 5397
rect 126853 5396 126859 5397
rect 127611 5396 127614 5402
rect 126853 5382 127614 5396
rect 126853 5380 126859 5382
rect 126830 5377 126859 5380
rect 127611 5376 127614 5382
rect 127640 5376 127643 5402
rect 133269 5396 133272 5402
rect 133249 5382 133272 5396
rect 133269 5376 133272 5382
rect 133298 5376 133301 5402
rect 133868 5397 133897 5400
rect 133868 5380 133874 5397
rect 133891 5396 133897 5397
rect 134097 5396 134100 5402
rect 133891 5382 134100 5396
rect 133891 5380 133897 5382
rect 133868 5377 133897 5380
rect 134097 5376 134100 5382
rect 134126 5376 134129 5402
rect 134190 5397 134219 5400
rect 134190 5380 134196 5397
rect 134213 5396 134219 5397
rect 134695 5396 134698 5402
rect 134213 5382 134698 5396
rect 134213 5380 134219 5382
rect 134190 5377 134219 5380
rect 134695 5376 134698 5382
rect 134724 5376 134727 5402
rect 97527 5362 97530 5368
rect 96892 5348 97530 5362
rect 96746 5343 96775 5346
rect 97527 5342 97530 5348
rect 97556 5342 97559 5368
rect 132441 5342 132444 5368
rect 132470 5362 132473 5368
rect 135017 5362 135020 5368
rect 132470 5348 133246 5362
rect 132470 5342 132473 5348
rect 96332 5329 96361 5332
rect 96332 5312 96338 5329
rect 96355 5312 96361 5329
rect 97067 5328 97070 5334
rect 97047 5314 97070 5328
rect 96332 5309 96361 5312
rect 97067 5308 97070 5314
rect 97096 5328 97099 5334
rect 97481 5328 97484 5334
rect 97096 5314 97484 5328
rect 97096 5308 97099 5314
rect 97481 5308 97484 5314
rect 97510 5308 97513 5334
rect 101530 5329 101559 5332
rect 101530 5312 101536 5329
rect 101553 5328 101559 5329
rect 102403 5328 102406 5334
rect 101553 5314 102406 5328
rect 101553 5312 101559 5314
rect 101530 5309 101559 5312
rect 102403 5308 102406 5314
rect 102432 5308 102435 5334
rect 126922 5329 126951 5332
rect 126922 5312 126928 5329
rect 126945 5328 126951 5329
rect 127473 5328 127476 5334
rect 126945 5314 127476 5328
rect 126945 5312 126951 5314
rect 126922 5309 126951 5312
rect 127473 5308 127476 5314
rect 127502 5308 127505 5334
rect 132994 5329 133023 5332
rect 132994 5312 133000 5329
rect 133017 5328 133023 5329
rect 133177 5328 133180 5334
rect 133017 5314 133180 5328
rect 133017 5312 133023 5314
rect 132994 5309 133023 5312
rect 133177 5308 133180 5314
rect 133206 5308 133209 5334
rect 133232 5332 133246 5348
rect 133968 5348 135020 5362
rect 133968 5332 133982 5348
rect 135017 5342 135020 5348
rect 135046 5342 135049 5368
rect 133224 5329 133253 5332
rect 133224 5312 133230 5329
rect 133247 5328 133253 5329
rect 133546 5329 133575 5332
rect 133546 5328 133552 5329
rect 133247 5314 133552 5328
rect 133247 5312 133253 5314
rect 133224 5309 133253 5312
rect 133546 5312 133552 5314
rect 133569 5312 133575 5329
rect 133546 5309 133575 5312
rect 133960 5329 133989 5332
rect 133960 5312 133966 5329
rect 133983 5312 133989 5329
rect 133960 5309 133989 5312
rect 134282 5329 134311 5332
rect 134282 5312 134288 5329
rect 134305 5312 134311 5329
rect 134282 5309 134311 5312
rect 93755 5294 93758 5300
rect 93735 5280 93758 5294
rect 93755 5274 93758 5280
rect 93784 5274 93787 5300
rect 100517 5294 100520 5300
rect 96432 5280 100520 5294
rect 15165 5246 15877 5260
rect 95550 5261 95579 5264
rect 15165 5244 15171 5246
rect 15142 5241 15171 5244
rect 95550 5244 95556 5261
rect 95573 5260 95579 5261
rect 96055 5260 96058 5266
rect 95573 5246 96058 5260
rect 95573 5244 95579 5246
rect 95550 5241 95579 5244
rect 96055 5240 96058 5246
rect 96084 5240 96087 5266
rect 96432 5264 96446 5280
rect 100517 5274 100520 5280
rect 100546 5274 100549 5300
rect 134290 5294 134304 5309
rect 134511 5308 134514 5334
rect 134540 5328 134543 5334
rect 134558 5329 134587 5332
rect 134558 5328 134564 5329
rect 134540 5314 134564 5328
rect 134540 5308 134543 5314
rect 134558 5312 134564 5314
rect 134581 5312 134587 5329
rect 134558 5309 134587 5312
rect 134604 5329 134633 5332
rect 134604 5312 134610 5329
rect 134627 5328 134633 5329
rect 135155 5328 135158 5334
rect 134627 5314 135158 5328
rect 134627 5312 134633 5314
rect 134604 5309 134633 5312
rect 135155 5308 135158 5314
rect 135184 5308 135187 5334
rect 136259 5294 136262 5300
rect 134290 5280 136262 5294
rect 136259 5274 136262 5280
rect 136288 5274 136291 5300
rect 96424 5261 96453 5264
rect 96424 5244 96430 5261
rect 96447 5244 96453 5261
rect 96424 5241 96453 5244
rect 96838 5261 96867 5264
rect 96838 5244 96844 5261
rect 96861 5260 96867 5261
rect 133592 5261 133621 5264
rect 96861 5246 98424 5260
rect 96861 5244 96867 5246
rect 96838 5241 96867 5244
rect 78806 5227 78835 5230
rect 78806 5210 78812 5227
rect 78829 5226 78835 5227
rect 89569 5226 89572 5232
rect 78829 5212 89572 5226
rect 78829 5210 78835 5212
rect 78806 5207 78835 5210
rect 89569 5206 89572 5212
rect 89598 5206 89601 5232
rect 98410 5226 98424 5246
rect 133592 5244 133598 5261
rect 133615 5260 133621 5261
rect 134373 5260 134376 5266
rect 133615 5246 134376 5260
rect 133615 5244 133621 5246
rect 133592 5241 133621 5244
rect 134373 5240 134376 5246
rect 134402 5240 134405 5266
rect 101759 5226 101762 5232
rect 98410 5212 101762 5226
rect 101759 5206 101762 5212
rect 101788 5206 101791 5232
rect 132902 5227 132931 5230
rect 132902 5210 132908 5227
rect 132925 5226 132931 5227
rect 134787 5226 134790 5232
rect 132925 5212 134790 5226
rect 132925 5210 132931 5212
rect 132902 5207 132931 5210
rect 134787 5206 134790 5212
rect 134816 5206 134819 5232
rect 552 5181 152904 5192
rect 552 5155 19524 5181
rect 19550 5155 19556 5181
rect 19582 5155 19588 5181
rect 19614 5155 19620 5181
rect 19646 5155 19652 5181
rect 19678 5155 57623 5181
rect 57649 5155 57655 5181
rect 57681 5155 57687 5181
rect 57713 5155 57719 5181
rect 57745 5155 57751 5181
rect 57777 5155 95722 5181
rect 95748 5155 95754 5181
rect 95780 5155 95786 5181
rect 95812 5155 95818 5181
rect 95844 5155 95850 5181
rect 95876 5155 133821 5181
rect 133847 5155 133853 5181
rect 133879 5155 133885 5181
rect 133911 5155 133917 5181
rect 133943 5155 133949 5181
rect 133975 5155 152904 5181
rect 552 5144 152904 5155
rect 15049 5104 15052 5130
rect 15078 5124 15081 5130
rect 15464 5125 15493 5128
rect 15464 5124 15470 5125
rect 15078 5110 15470 5124
rect 15078 5104 15081 5110
rect 15464 5108 15470 5110
rect 15487 5108 15493 5125
rect 15831 5124 15834 5130
rect 15811 5110 15834 5124
rect 15464 5105 15493 5108
rect 15831 5104 15834 5110
rect 15860 5104 15863 5130
rect 16061 5104 16064 5130
rect 16090 5124 16093 5130
rect 16430 5125 16459 5128
rect 16430 5124 16436 5125
rect 16090 5110 16436 5124
rect 16090 5104 16093 5110
rect 16430 5108 16436 5110
rect 16453 5108 16459 5125
rect 16430 5105 16459 5108
rect 16659 5104 16662 5130
rect 16688 5124 16691 5130
rect 16798 5125 16827 5128
rect 16798 5124 16804 5125
rect 16688 5110 16804 5124
rect 16688 5104 16691 5110
rect 16798 5108 16804 5110
rect 16821 5108 16827 5125
rect 16798 5105 16827 5108
rect 95641 5104 95644 5130
rect 95670 5124 95673 5130
rect 95918 5125 95947 5128
rect 95918 5124 95924 5125
rect 95670 5110 95924 5124
rect 95670 5104 95673 5110
rect 95918 5108 95924 5110
rect 95941 5108 95947 5125
rect 95918 5105 95947 5108
rect 96239 5104 96242 5130
rect 96268 5124 96271 5130
rect 96562 5125 96591 5128
rect 96562 5124 96568 5125
rect 96268 5110 96568 5124
rect 96268 5104 96271 5110
rect 96562 5108 96568 5110
rect 96585 5108 96591 5125
rect 96562 5105 96591 5108
rect 133453 5104 133456 5130
rect 133482 5124 133485 5130
rect 133868 5125 133897 5128
rect 133868 5124 133874 5125
rect 133482 5110 133874 5124
rect 133482 5104 133485 5110
rect 133868 5108 133874 5110
rect 133891 5108 133897 5125
rect 133868 5105 133897 5108
rect 134281 5104 134284 5130
rect 134310 5124 134313 5130
rect 134512 5125 134541 5128
rect 134512 5124 134518 5125
rect 134310 5110 134518 5124
rect 134310 5104 134313 5110
rect 134512 5108 134518 5110
rect 134535 5108 134541 5125
rect 134512 5105 134541 5108
rect 13761 5070 13764 5096
rect 13790 5090 13793 5096
rect 15142 5091 15171 5094
rect 15142 5090 15148 5091
rect 13790 5076 15148 5090
rect 13790 5070 13793 5076
rect 15142 5074 15148 5076
rect 15165 5074 15171 5091
rect 15142 5071 15171 5074
rect 15785 5070 15788 5096
rect 15814 5090 15817 5096
rect 16154 5091 16183 5094
rect 16154 5090 16160 5091
rect 15814 5076 16160 5090
rect 15814 5070 15817 5076
rect 16154 5074 16160 5076
rect 16177 5074 16183 5091
rect 16154 5071 16183 5074
rect 133546 5091 133575 5094
rect 133546 5074 133552 5091
rect 133569 5090 133575 5091
rect 134189 5090 134192 5096
rect 133569 5076 133867 5090
rect 133569 5074 133575 5076
rect 133546 5071 133575 5074
rect 133853 5062 133867 5076
rect 133922 5076 134192 5090
rect 78898 5057 78927 5060
rect 78898 5040 78904 5057
rect 78921 5056 78927 5057
rect 81795 5056 81798 5062
rect 78921 5042 81798 5056
rect 78921 5040 78927 5042
rect 78898 5037 78927 5040
rect 81795 5036 81798 5042
rect 81824 5036 81827 5062
rect 97941 5056 97944 5062
rect 96340 5042 97944 5056
rect 14727 5002 14730 5028
rect 14756 5022 14759 5028
rect 15234 5023 15263 5026
rect 15234 5022 15240 5023
rect 14756 5008 15240 5022
rect 14756 5002 14759 5008
rect 15234 5006 15240 5008
rect 15257 5006 15263 5023
rect 15234 5003 15263 5006
rect 15463 5002 15466 5028
rect 15492 5022 15495 5028
rect 15556 5023 15585 5026
rect 15556 5022 15562 5023
rect 15492 5008 15562 5022
rect 15492 5002 15495 5008
rect 15556 5006 15562 5008
rect 15579 5006 15585 5023
rect 15556 5003 15585 5006
rect 15786 5023 15815 5026
rect 15786 5006 15792 5023
rect 15809 5022 15815 5023
rect 16108 5023 16137 5026
rect 16108 5022 16114 5023
rect 15809 5008 16114 5022
rect 15809 5006 15815 5008
rect 15786 5003 15815 5006
rect 16108 5006 16114 5008
rect 16131 5006 16137 5023
rect 16108 5003 16137 5006
rect 16522 5023 16551 5026
rect 16522 5006 16528 5023
rect 16545 5022 16551 5023
rect 16705 5022 16708 5028
rect 16545 5008 16708 5022
rect 16545 5006 16551 5008
rect 16522 5003 16551 5006
rect 16116 4988 16130 5003
rect 16705 5002 16708 5008
rect 16734 5002 16737 5028
rect 16752 5023 16781 5026
rect 16752 5006 16758 5023
rect 16775 5022 16781 5023
rect 16843 5022 16846 5028
rect 16775 5008 16846 5022
rect 16775 5006 16781 5008
rect 16752 5003 16781 5006
rect 16760 4988 16774 5003
rect 16843 5002 16846 5008
rect 16872 5002 16875 5028
rect 70204 5023 70233 5026
rect 70204 5006 70210 5023
rect 70227 5022 70233 5023
rect 70341 5022 70344 5028
rect 70227 5008 70344 5022
rect 70227 5006 70233 5008
rect 70204 5003 70233 5006
rect 70341 5002 70344 5008
rect 70370 5002 70373 5028
rect 78024 5023 78053 5026
rect 78024 5006 78030 5023
rect 78047 5022 78053 5023
rect 78069 5022 78072 5028
rect 78047 5008 78072 5022
rect 78047 5006 78053 5008
rect 78024 5003 78053 5006
rect 78069 5002 78072 5008
rect 78098 5002 78101 5028
rect 96010 5023 96039 5026
rect 96010 5006 96016 5023
rect 96033 5022 96039 5023
rect 96285 5022 96288 5028
rect 96033 5008 96288 5022
rect 96033 5006 96039 5008
rect 96010 5003 96039 5006
rect 96285 5002 96288 5008
rect 96314 5002 96317 5028
rect 96340 5026 96354 5042
rect 97941 5036 97944 5042
rect 97970 5036 97973 5062
rect 133853 5042 133870 5062
rect 133867 5036 133870 5042
rect 133896 5036 133899 5062
rect 96332 5023 96361 5026
rect 96332 5006 96338 5023
rect 96355 5006 96361 5023
rect 96332 5003 96361 5006
rect 96654 5023 96683 5026
rect 96654 5006 96660 5023
rect 96677 5022 96683 5023
rect 97205 5022 97208 5028
rect 96677 5008 97208 5022
rect 96677 5006 96683 5008
rect 96654 5003 96683 5006
rect 97205 5002 97208 5008
rect 97234 5002 97237 5028
rect 133638 5023 133667 5026
rect 133638 5006 133644 5023
rect 133661 5022 133667 5023
rect 133922 5022 133936 5076
rect 134189 5070 134192 5076
rect 134218 5070 134221 5096
rect 134236 5091 134265 5094
rect 134236 5074 134242 5091
rect 134259 5090 134265 5091
rect 134741 5090 134744 5096
rect 134259 5076 134744 5090
rect 134259 5074 134265 5076
rect 134236 5071 134265 5074
rect 134741 5070 134744 5076
rect 134770 5070 134773 5096
rect 134419 5056 134422 5062
rect 133968 5042 134422 5056
rect 133968 5026 133982 5042
rect 134419 5036 134422 5042
rect 134448 5036 134451 5062
rect 133661 5008 133936 5022
rect 133960 5023 133989 5026
rect 133661 5006 133667 5008
rect 133638 5003 133667 5006
rect 133960 5006 133966 5023
rect 133983 5006 133989 5023
rect 133960 5003 133989 5006
rect 134051 5002 134054 5028
rect 134080 5022 134083 5028
rect 134190 5023 134219 5026
rect 134190 5022 134196 5023
rect 134080 5008 134196 5022
rect 134080 5002 134083 5008
rect 134190 5006 134196 5008
rect 134213 5022 134219 5023
rect 134511 5022 134514 5028
rect 134213 5008 134514 5022
rect 134213 5006 134219 5008
rect 134190 5003 134219 5006
rect 134511 5002 134514 5008
rect 134540 5002 134543 5028
rect 134603 5022 134606 5028
rect 134583 5008 134606 5022
rect 134603 5002 134606 5008
rect 134632 5002 134635 5028
rect 152221 5022 152224 5028
rect 152201 5008 152224 5022
rect 152221 5002 152224 5008
rect 152250 5002 152253 5028
rect 16116 4974 16774 4988
rect 126369 4968 126372 4994
rect 126398 4988 126401 4994
rect 152406 4989 152435 4992
rect 152406 4988 152412 4989
rect 126398 4974 152412 4988
rect 126398 4968 126401 4974
rect 152406 4972 152412 4974
rect 152429 4972 152435 4989
rect 152406 4969 152435 4972
rect 58703 4934 58706 4960
rect 58732 4954 58735 4960
rect 70848 4955 70877 4958
rect 70848 4954 70854 4955
rect 58732 4940 70854 4954
rect 58732 4934 58735 4940
rect 70848 4938 70854 4940
rect 70871 4938 70877 4955
rect 70848 4935 70877 4938
rect 96240 4955 96269 4958
rect 96240 4938 96246 4955
rect 96263 4954 96269 4955
rect 97159 4954 97162 4960
rect 96263 4940 97162 4954
rect 96263 4938 96269 4940
rect 96240 4935 96269 4938
rect 97159 4934 97162 4940
rect 97188 4934 97191 4960
rect 133867 4934 133870 4960
rect 133896 4954 133899 4960
rect 135477 4954 135480 4960
rect 133896 4940 135480 4954
rect 133896 4934 133899 4940
rect 135477 4934 135480 4940
rect 135506 4934 135509 4960
rect 552 4909 152904 4920
rect 552 4883 38574 4909
rect 38600 4883 38606 4909
rect 38632 4883 38638 4909
rect 38664 4883 38670 4909
rect 38696 4883 38702 4909
rect 38728 4883 76673 4909
rect 76699 4883 76705 4909
rect 76731 4883 76737 4909
rect 76763 4883 76769 4909
rect 76795 4883 76801 4909
rect 76827 4883 114772 4909
rect 114798 4883 114804 4909
rect 114830 4883 114836 4909
rect 114862 4883 114868 4909
rect 114894 4883 114900 4909
rect 114926 4883 152904 4909
rect 552 4872 152904 4883
rect 15601 4798 15604 4824
rect 15630 4818 15633 4824
rect 16430 4819 16459 4822
rect 16430 4818 16436 4819
rect 15630 4804 16436 4818
rect 15630 4798 15633 4804
rect 16430 4802 16436 4804
rect 16453 4802 16459 4819
rect 70341 4818 70344 4824
rect 70321 4804 70344 4818
rect 16430 4799 16459 4802
rect 70341 4798 70344 4804
rect 70370 4798 70373 4824
rect 78069 4818 78072 4824
rect 78049 4804 78072 4818
rect 78069 4798 78072 4804
rect 78098 4798 78101 4824
rect 78944 4819 78973 4822
rect 78944 4802 78950 4819
rect 78967 4818 78973 4819
rect 79311 4818 79314 4824
rect 78967 4804 79314 4818
rect 78967 4802 78973 4804
rect 78944 4799 78973 4802
rect 79311 4798 79314 4804
rect 79340 4798 79343 4824
rect 95319 4798 95322 4824
rect 95348 4818 95351 4824
rect 96516 4819 96545 4822
rect 95348 4804 96492 4818
rect 95348 4798 95351 4804
rect 13669 4764 13672 4790
rect 13698 4784 13701 4790
rect 15648 4785 15677 4788
rect 15648 4784 15654 4785
rect 13698 4770 15654 4784
rect 13698 4764 13701 4770
rect 15648 4768 15654 4770
rect 15671 4768 15677 4785
rect 15648 4765 15677 4768
rect 16062 4785 16091 4788
rect 16062 4768 16068 4785
rect 16085 4784 16091 4785
rect 16384 4785 16413 4788
rect 16384 4784 16390 4785
rect 16085 4770 16390 4784
rect 16085 4768 16091 4770
rect 16062 4765 16091 4768
rect 16384 4768 16390 4770
rect 16407 4784 16413 4785
rect 16843 4784 16846 4790
rect 16407 4770 16846 4784
rect 16407 4768 16413 4770
rect 16384 4765 16413 4768
rect 16843 4764 16846 4770
rect 16872 4764 16875 4790
rect 96478 4788 96492 4804
rect 96516 4802 96522 4819
rect 96539 4818 96545 4819
rect 96653 4818 96656 4824
rect 96539 4804 96656 4818
rect 96539 4802 96545 4804
rect 96516 4799 96545 4802
rect 96653 4798 96656 4804
rect 96682 4798 96685 4824
rect 133960 4819 133989 4822
rect 133960 4802 133966 4819
rect 133983 4818 133989 4819
rect 134925 4818 134928 4824
rect 133983 4804 134928 4818
rect 133983 4802 133989 4804
rect 133960 4799 133989 4802
rect 134925 4798 134928 4804
rect 134954 4798 134957 4824
rect 96240 4785 96269 4788
rect 96240 4768 96246 4785
rect 96263 4768 96269 4785
rect 96240 4765 96269 4768
rect 96470 4785 96499 4788
rect 96470 4768 96476 4785
rect 96493 4784 96499 4785
rect 97067 4784 97070 4790
rect 96493 4770 97070 4784
rect 96493 4768 96499 4770
rect 96470 4765 96499 4768
rect 15279 4730 15282 4756
rect 15308 4750 15311 4756
rect 16108 4751 16137 4754
rect 16108 4750 16114 4751
rect 15308 4736 16114 4750
rect 15308 4730 15311 4736
rect 16108 4734 16114 4736
rect 16131 4734 16137 4751
rect 96248 4750 96262 4765
rect 97067 4764 97070 4770
rect 97096 4764 97099 4790
rect 133914 4785 133943 4788
rect 133914 4768 133920 4785
rect 133937 4784 133943 4785
rect 134051 4784 134054 4790
rect 133937 4770 134054 4784
rect 133937 4768 133943 4770
rect 133914 4765 133943 4768
rect 134051 4764 134054 4770
rect 134080 4764 134083 4790
rect 97987 4750 97990 4756
rect 96248 4736 97990 4750
rect 16108 4731 16137 4734
rect 97987 4730 97990 4736
rect 98016 4730 98019 4756
rect 14957 4696 14960 4722
rect 14986 4716 14989 4722
rect 15556 4717 15585 4720
rect 15556 4716 15562 4717
rect 14986 4702 15562 4716
rect 14986 4696 14989 4702
rect 15556 4700 15562 4702
rect 15579 4700 15585 4717
rect 15556 4697 15585 4700
rect 96148 4717 96177 4720
rect 96148 4700 96154 4717
rect 96171 4716 96177 4717
rect 97251 4716 97254 4722
rect 96171 4702 97254 4716
rect 96171 4700 96177 4702
rect 96148 4697 96177 4700
rect 97251 4696 97254 4702
rect 97280 4696 97283 4722
rect 52125 4662 52128 4688
rect 52154 4682 52157 4688
rect 70986 4683 71015 4686
rect 70986 4682 70992 4683
rect 52154 4668 70992 4682
rect 52154 4662 52157 4668
rect 70986 4666 70992 4668
rect 71009 4682 71015 4683
rect 74159 4682 74162 4688
rect 71009 4668 74162 4682
rect 71009 4666 71015 4668
rect 70986 4663 71015 4666
rect 74159 4662 74162 4668
rect 74188 4662 74191 4688
rect 552 4637 152904 4648
rect 552 4611 19524 4637
rect 19550 4611 19556 4637
rect 19582 4611 19588 4637
rect 19614 4611 19620 4637
rect 19646 4611 19652 4637
rect 19678 4611 57623 4637
rect 57649 4611 57655 4637
rect 57681 4611 57687 4637
rect 57713 4611 57719 4637
rect 57745 4611 57751 4637
rect 57777 4611 95722 4637
rect 95748 4611 95754 4637
rect 95780 4611 95786 4637
rect 95812 4611 95818 4637
rect 95844 4611 95850 4637
rect 95876 4611 133821 4637
rect 133847 4611 133853 4637
rect 133879 4611 133885 4637
rect 133911 4611 133917 4637
rect 133943 4611 133949 4637
rect 133975 4611 152904 4637
rect 552 4600 152904 4611
rect 552 4365 152904 4376
rect 552 4339 38574 4365
rect 38600 4339 38606 4365
rect 38632 4339 38638 4365
rect 38664 4339 38670 4365
rect 38696 4339 38702 4365
rect 38728 4339 76673 4365
rect 76699 4339 76705 4365
rect 76731 4339 76737 4365
rect 76763 4339 76769 4365
rect 76795 4339 76801 4365
rect 76827 4339 114772 4365
rect 114798 4339 114804 4365
rect 114830 4339 114836 4365
rect 114862 4339 114868 4365
rect 114894 4339 114900 4365
rect 114926 4339 152904 4365
rect 552 4328 152904 4339
rect 790 4241 819 4244
rect 790 4224 796 4241
rect 813 4240 819 4241
rect 813 4226 996 4240
rect 813 4224 819 4226
rect 790 4221 819 4224
rect 697 4172 700 4178
rect 677 4158 700 4172
rect 697 4152 700 4158
rect 726 4152 729 4178
rect 982 4176 996 4226
rect 974 4173 1003 4176
rect 974 4156 980 4173
rect 997 4172 1003 4173
rect 1158 4173 1187 4176
rect 1158 4172 1164 4173
rect 997 4158 1164 4172
rect 997 4156 1003 4158
rect 974 4153 1003 4156
rect 1158 4156 1164 4158
rect 1181 4172 1187 4173
rect 1342 4173 1371 4176
rect 1342 4172 1348 4173
rect 1181 4158 1348 4172
rect 1181 4156 1187 4158
rect 1158 4153 1187 4156
rect 1342 4156 1348 4158
rect 1365 4172 1371 4173
rect 1526 4173 1555 4176
rect 1526 4172 1532 4173
rect 1365 4158 1532 4172
rect 1365 4156 1371 4158
rect 1342 4153 1371 4156
rect 1526 4156 1532 4158
rect 1549 4172 1555 4173
rect 93755 4172 93758 4178
rect 1549 4158 93758 4172
rect 1549 4156 1555 4158
rect 1526 4153 1555 4156
rect 93755 4152 93758 4158
rect 93784 4152 93787 4178
rect 552 4093 152904 4104
rect 552 4067 19524 4093
rect 19550 4067 19556 4093
rect 19582 4067 19588 4093
rect 19614 4067 19620 4093
rect 19646 4067 19652 4093
rect 19678 4067 57623 4093
rect 57649 4067 57655 4093
rect 57681 4067 57687 4093
rect 57713 4067 57719 4093
rect 57745 4067 57751 4093
rect 57777 4067 95722 4093
rect 95748 4067 95754 4093
rect 95780 4067 95786 4093
rect 95812 4067 95818 4093
rect 95844 4067 95850 4093
rect 95876 4067 133821 4093
rect 133847 4067 133853 4093
rect 133879 4067 133885 4093
rect 133911 4067 133917 4093
rect 133943 4067 133949 4093
rect 133975 4067 152904 4093
rect 552 4056 152904 4067
rect 552 3821 152904 3832
rect 552 3795 38574 3821
rect 38600 3795 38606 3821
rect 38632 3795 38638 3821
rect 38664 3795 38670 3821
rect 38696 3795 38702 3821
rect 38728 3795 76673 3821
rect 76699 3795 76705 3821
rect 76731 3795 76737 3821
rect 76763 3795 76769 3821
rect 76795 3795 76801 3821
rect 76827 3795 114772 3821
rect 114798 3795 114804 3821
rect 114830 3795 114836 3821
rect 114862 3795 114868 3821
rect 114894 3795 114900 3821
rect 114926 3795 152904 3821
rect 552 3784 152904 3795
rect 552 3549 152904 3560
rect 552 3523 19524 3549
rect 19550 3523 19556 3549
rect 19582 3523 19588 3549
rect 19614 3523 19620 3549
rect 19646 3523 19652 3549
rect 19678 3523 57623 3549
rect 57649 3523 57655 3549
rect 57681 3523 57687 3549
rect 57713 3523 57719 3549
rect 57745 3523 57751 3549
rect 57777 3523 95722 3549
rect 95748 3523 95754 3549
rect 95780 3523 95786 3549
rect 95812 3523 95818 3549
rect 95844 3523 95850 3549
rect 95876 3523 133821 3549
rect 133847 3523 133853 3549
rect 133879 3523 133885 3549
rect 133911 3523 133917 3549
rect 133943 3523 133949 3549
rect 133975 3523 152904 3549
rect 552 3512 152904 3523
rect 552 3277 152904 3288
rect 552 3251 38574 3277
rect 38600 3251 38606 3277
rect 38632 3251 38638 3277
rect 38664 3251 38670 3277
rect 38696 3251 38702 3277
rect 38728 3251 76673 3277
rect 76699 3251 76705 3277
rect 76731 3251 76737 3277
rect 76763 3251 76769 3277
rect 76795 3251 76801 3277
rect 76827 3251 114772 3277
rect 114798 3251 114804 3277
rect 114830 3251 114836 3277
rect 114862 3251 114868 3277
rect 114894 3251 114900 3277
rect 114926 3251 152904 3277
rect 552 3240 152904 3251
rect 151991 3152 151994 3158
rect 151971 3138 151994 3152
rect 151991 3132 151994 3138
rect 152020 3132 152023 3158
rect 124529 3098 124532 3124
rect 124558 3118 124561 3124
rect 152130 3119 152159 3122
rect 152130 3118 152136 3119
rect 124558 3104 152136 3118
rect 124558 3098 124561 3104
rect 152130 3102 152136 3104
rect 152153 3102 152159 3119
rect 152130 3099 152159 3102
rect 552 3005 152904 3016
rect 552 2979 19524 3005
rect 19550 2979 19556 3005
rect 19582 2979 19588 3005
rect 19614 2979 19620 3005
rect 19646 2979 19652 3005
rect 19678 2979 57623 3005
rect 57649 2979 57655 3005
rect 57681 2979 57687 3005
rect 57713 2979 57719 3005
rect 57745 2979 57751 3005
rect 57777 2979 95722 3005
rect 95748 2979 95754 3005
rect 95780 2979 95786 3005
rect 95812 2979 95818 3005
rect 95844 2979 95850 3005
rect 95876 2979 133821 3005
rect 133847 2979 133853 3005
rect 133879 2979 133885 3005
rect 133911 2979 133917 3005
rect 133943 2979 133949 3005
rect 133975 2979 152904 3005
rect 552 2968 152904 2979
rect 552 2733 152904 2744
rect 552 2707 38574 2733
rect 38600 2707 38606 2733
rect 38632 2707 38638 2733
rect 38664 2707 38670 2733
rect 38696 2707 38702 2733
rect 38728 2707 76673 2733
rect 76699 2707 76705 2733
rect 76731 2707 76737 2733
rect 76763 2707 76769 2733
rect 76795 2707 76801 2733
rect 76827 2707 114772 2733
rect 114798 2707 114804 2733
rect 114830 2707 114836 2733
rect 114862 2707 114868 2733
rect 114894 2707 114900 2733
rect 114926 2707 152904 2733
rect 552 2696 152904 2707
rect 552 2461 152904 2472
rect 552 2435 19524 2461
rect 19550 2435 19556 2461
rect 19582 2435 19588 2461
rect 19614 2435 19620 2461
rect 19646 2435 19652 2461
rect 19678 2435 57623 2461
rect 57649 2435 57655 2461
rect 57681 2435 57687 2461
rect 57713 2435 57719 2461
rect 57745 2435 57751 2461
rect 57777 2435 95722 2461
rect 95748 2435 95754 2461
rect 95780 2435 95786 2461
rect 95812 2435 95818 2461
rect 95844 2435 95850 2461
rect 95876 2435 133821 2461
rect 133847 2435 133853 2461
rect 133879 2435 133885 2461
rect 133911 2435 133917 2461
rect 133943 2435 133949 2461
rect 133975 2435 152904 2461
rect 552 2424 152904 2435
rect 552 2189 152904 2200
rect 552 2163 38574 2189
rect 38600 2163 38606 2189
rect 38632 2163 38638 2189
rect 38664 2163 38670 2189
rect 38696 2163 38702 2189
rect 38728 2163 76673 2189
rect 76699 2163 76705 2189
rect 76731 2163 76737 2189
rect 76763 2163 76769 2189
rect 76795 2163 76801 2189
rect 76827 2163 114772 2189
rect 114798 2163 114804 2189
rect 114830 2163 114836 2189
rect 114862 2163 114868 2189
rect 114894 2163 114900 2189
rect 114926 2163 152904 2189
rect 552 2152 152904 2163
rect 552 1917 152904 1928
rect 552 1891 19524 1917
rect 19550 1891 19556 1917
rect 19582 1891 19588 1917
rect 19614 1891 19620 1917
rect 19646 1891 19652 1917
rect 19678 1891 57623 1917
rect 57649 1891 57655 1917
rect 57681 1891 57687 1917
rect 57713 1891 57719 1917
rect 57745 1891 57751 1917
rect 57777 1891 95722 1917
rect 95748 1891 95754 1917
rect 95780 1891 95786 1917
rect 95812 1891 95818 1917
rect 95844 1891 95850 1917
rect 95876 1891 133821 1917
rect 133847 1891 133853 1917
rect 133879 1891 133885 1917
rect 133911 1891 133917 1917
rect 133943 1891 133949 1917
rect 133975 1891 152904 1917
rect 552 1880 152904 1891
rect 552 1645 152904 1656
rect 552 1619 38574 1645
rect 38600 1619 38606 1645
rect 38632 1619 38638 1645
rect 38664 1619 38670 1645
rect 38696 1619 38702 1645
rect 38728 1619 76673 1645
rect 76699 1619 76705 1645
rect 76731 1619 76737 1645
rect 76763 1619 76769 1645
rect 76795 1619 76801 1645
rect 76827 1619 114772 1645
rect 114798 1619 114804 1645
rect 114830 1619 114836 1645
rect 114862 1619 114868 1645
rect 114894 1619 114900 1645
rect 114926 1619 152904 1645
rect 552 1608 152904 1619
rect 552 1373 152904 1384
rect 552 1347 19524 1373
rect 19550 1347 19556 1373
rect 19582 1347 19588 1373
rect 19614 1347 19620 1373
rect 19646 1347 19652 1373
rect 19678 1347 57623 1373
rect 57649 1347 57655 1373
rect 57681 1347 57687 1373
rect 57713 1347 57719 1373
rect 57745 1347 57751 1373
rect 57777 1347 95722 1373
rect 95748 1347 95754 1373
rect 95780 1347 95786 1373
rect 95812 1347 95818 1373
rect 95844 1347 95850 1373
rect 95876 1347 133821 1373
rect 133847 1347 133853 1373
rect 133879 1347 133885 1373
rect 133911 1347 133917 1373
rect 133943 1347 133949 1373
rect 133975 1347 152904 1373
rect 552 1336 152904 1347
rect 74711 1296 74714 1322
rect 74740 1316 74743 1322
rect 151117 1316 151120 1322
rect 74740 1302 151120 1316
rect 74740 1296 74743 1302
rect 151117 1296 151120 1302
rect 151146 1296 151149 1322
rect 552 1101 152904 1112
rect 552 1075 38574 1101
rect 38600 1075 38606 1101
rect 38632 1075 38638 1101
rect 38664 1075 38670 1101
rect 38696 1075 38702 1101
rect 38728 1075 76673 1101
rect 76699 1075 76705 1101
rect 76731 1075 76737 1101
rect 76763 1075 76769 1101
rect 76795 1075 76801 1101
rect 76827 1075 114772 1101
rect 114798 1075 114804 1101
rect 114830 1075 114836 1101
rect 114862 1075 114868 1101
rect 114894 1075 114900 1101
rect 114926 1075 152904 1101
rect 552 1064 152904 1075
<< via1 >>
rect 14500 6872 14526 6898
rect 16478 6872 16504 6898
rect 23102 6872 23128 6898
rect 31704 6872 31730 6898
rect 34648 6872 34674 6898
rect 37684 6872 37710 6898
rect 38006 6872 38032 6898
rect 45320 6872 45346 6898
rect 51208 6872 51234 6898
rect 56912 6872 56938 6898
rect 62754 6872 62780 6898
rect 65928 6872 65954 6898
rect 80832 6872 80858 6898
rect 83040 6872 83066 6898
rect 83684 6872 83710 6898
rect 87088 6872 87114 6898
rect 88882 6872 88908 6898
rect 90952 6872 90978 6898
rect 94954 6906 94980 6932
rect 94678 6872 94704 6898
rect 96610 6872 96636 6898
rect 97990 6872 98016 6898
rect 151396 6872 151422 6898
rect 13580 6838 13606 6864
rect 18272 6838 18298 6864
rect 21262 6838 21288 6864
rect 23930 6838 23956 6864
rect 25816 6838 25842 6864
rect 27058 6838 27084 6864
rect 33084 6838 33110 6864
rect 36212 6838 36238 6864
rect 36948 6838 36974 6864
rect 38190 6838 38216 6864
rect 41548 6838 41574 6864
rect 43204 6838 43230 6864
rect 45918 6838 45944 6864
rect 50978 6838 51004 6864
rect 57326 6838 57352 6864
rect 63720 6838 63746 6864
rect 63766 6838 63792 6864
rect 64870 6838 64896 6864
rect 66802 6838 66828 6864
rect 68412 6838 68438 6864
rect 74070 6838 74096 6864
rect 75220 6838 75246 6864
rect 78578 6838 78604 6864
rect 150706 6838 150732 6864
rect 19524 6787 19550 6813
rect 19556 6787 19582 6813
rect 19588 6787 19614 6813
rect 19620 6787 19646 6813
rect 19652 6787 19678 6813
rect 57623 6787 57649 6813
rect 57655 6787 57681 6813
rect 57687 6787 57713 6813
rect 57719 6787 57745 6813
rect 57751 6787 57777 6813
rect 95722 6787 95748 6813
rect 95754 6787 95780 6813
rect 95786 6787 95812 6813
rect 95818 6787 95844 6813
rect 95850 6787 95876 6813
rect 133821 6787 133847 6813
rect 133853 6787 133879 6813
rect 133885 6787 133911 6813
rect 133917 6787 133943 6813
rect 133949 6787 133975 6813
rect 792 6757 818 6762
rect 792 6740 796 6757
rect 796 6740 813 6757
rect 813 6740 818 6757
rect 792 6736 818 6740
rect 2310 6757 2336 6762
rect 2310 6740 2314 6757
rect 2314 6740 2331 6757
rect 2331 6740 2336 6757
rect 2310 6736 2336 6740
rect 3828 6757 3854 6762
rect 3828 6740 3832 6757
rect 3832 6740 3849 6757
rect 3849 6740 3854 6757
rect 3828 6736 3854 6740
rect 5392 6757 5418 6762
rect 5392 6740 5396 6757
rect 5396 6740 5413 6757
rect 5413 6740 5418 6757
rect 5392 6736 5418 6740
rect 6910 6736 6936 6762
rect 8428 6757 8454 6762
rect 8428 6740 8432 6757
rect 8432 6740 8449 6757
rect 8449 6740 8454 6757
rect 8428 6736 8454 6740
rect 9992 6757 10018 6762
rect 9992 6740 9996 6757
rect 9996 6740 10013 6757
rect 10013 6740 10018 6757
rect 9992 6736 10018 6740
rect 11510 6757 11536 6762
rect 11510 6740 11514 6757
rect 11514 6740 11531 6757
rect 11531 6740 11536 6757
rect 11510 6736 11536 6740
rect 13810 6736 13836 6762
rect 13856 6736 13882 6762
rect 15236 6736 15262 6762
rect 18272 6736 18298 6762
rect 23102 6736 23128 6762
rect 23792 6757 23818 6762
rect 23792 6740 23796 6757
rect 23796 6740 23813 6757
rect 23813 6740 23818 6757
rect 23792 6736 23818 6740
rect 25264 6736 25290 6762
rect 26506 6736 26532 6762
rect 27794 6736 27820 6762
rect 28944 6736 28970 6762
rect 30876 6736 30902 6762
rect 31704 6736 31730 6762
rect 71448 6757 71474 6762
rect 13580 6702 13606 6728
rect 22090 6702 22116 6728
rect 2402 6655 2428 6660
rect 2402 6638 2406 6655
rect 2406 6638 2423 6655
rect 2423 6638 2428 6655
rect 2402 6634 2428 6638
rect 7140 6655 7166 6660
rect 7140 6638 7144 6655
rect 7144 6638 7161 6655
rect 7161 6638 7166 6655
rect 7140 6634 7166 6638
rect 8520 6655 8546 6660
rect 8520 6638 8524 6655
rect 8524 6638 8541 6655
rect 8541 6638 8546 6655
rect 8520 6634 8546 6638
rect 10084 6655 10110 6660
rect 10084 6638 10088 6655
rect 10088 6638 10105 6655
rect 10105 6638 10110 6655
rect 10084 6634 10110 6638
rect 11602 6655 11628 6660
rect 11602 6638 11606 6655
rect 11606 6638 11623 6655
rect 11623 6638 11628 6655
rect 11602 6634 11628 6638
rect 13488 6668 13514 6694
rect 14914 6655 14940 6660
rect 14914 6638 14918 6655
rect 14918 6638 14935 6655
rect 14935 6638 14940 6655
rect 14914 6634 14940 6638
rect 16202 6655 16228 6660
rect 16202 6638 16206 6655
rect 16206 6638 16223 6655
rect 16223 6638 16228 6655
rect 16202 6634 16228 6638
rect 16892 6634 16918 6660
rect 22182 6702 22208 6728
rect 22780 6689 22806 6694
rect 22780 6672 22784 6689
rect 22784 6672 22801 6689
rect 22801 6672 22806 6689
rect 25816 6689 25842 6694
rect 22780 6668 22806 6672
rect 25816 6672 25820 6689
rect 25820 6672 25837 6689
rect 25837 6672 25842 6689
rect 25816 6668 25842 6672
rect 29910 6702 29936 6728
rect 31520 6723 31546 6728
rect 31520 6706 31524 6723
rect 31524 6706 31541 6723
rect 31541 6706 31546 6723
rect 31520 6702 31546 6706
rect 37684 6723 37710 6728
rect 36350 6689 36376 6694
rect 13764 6621 13790 6626
rect 13626 6566 13652 6592
rect 13764 6604 13768 6621
rect 13768 6604 13785 6621
rect 13785 6604 13790 6621
rect 13764 6600 13790 6604
rect 13856 6566 13882 6592
rect 15098 6600 15124 6626
rect 16340 6621 16366 6626
rect 15236 6566 15262 6592
rect 16340 6604 16344 6621
rect 16344 6604 16361 6621
rect 16361 6604 16366 6621
rect 16340 6600 16366 6604
rect 17260 6600 17286 6626
rect 17996 6600 18022 6626
rect 16800 6566 16826 6592
rect 17076 6587 17102 6592
rect 17076 6570 17080 6587
rect 17080 6570 17097 6587
rect 17097 6570 17102 6587
rect 17076 6566 17102 6570
rect 17168 6566 17194 6592
rect 18732 6566 18758 6592
rect 19468 6634 19494 6660
rect 18916 6621 18942 6626
rect 18916 6604 18920 6621
rect 18920 6604 18937 6621
rect 18937 6604 18942 6621
rect 18916 6600 18942 6604
rect 21262 6655 21288 6660
rect 19652 6587 19678 6592
rect 19652 6570 19656 6587
rect 19656 6570 19673 6587
rect 19673 6570 19678 6587
rect 19652 6566 19678 6570
rect 19974 6566 20000 6592
rect 21262 6638 21266 6655
rect 21266 6638 21283 6655
rect 21283 6638 21288 6655
rect 21262 6634 21288 6638
rect 22136 6634 22162 6660
rect 25678 6655 25704 6660
rect 20204 6621 20230 6626
rect 20204 6604 20208 6621
rect 20208 6604 20225 6621
rect 20225 6604 20230 6621
rect 20204 6600 20230 6604
rect 20710 6600 20736 6626
rect 21446 6600 21472 6626
rect 21630 6600 21656 6626
rect 21216 6566 21242 6592
rect 22504 6587 22530 6592
rect 22504 6570 22508 6587
rect 22508 6570 22525 6587
rect 22525 6570 22530 6587
rect 22504 6566 22530 6570
rect 22688 6587 22714 6592
rect 22688 6570 22692 6587
rect 22692 6570 22709 6587
rect 22709 6570 22714 6587
rect 22688 6566 22714 6570
rect 25678 6638 25682 6655
rect 25682 6638 25699 6655
rect 25699 6638 25704 6655
rect 25678 6634 25704 6638
rect 23930 6600 23956 6626
rect 27196 6634 27222 6660
rect 27380 6634 27406 6660
rect 27794 6655 27820 6660
rect 27794 6638 27798 6655
rect 27798 6638 27815 6655
rect 27815 6638 27820 6655
rect 27794 6634 27820 6638
rect 28944 6655 28970 6660
rect 28944 6638 28948 6655
rect 28948 6638 28965 6655
rect 28965 6638 28970 6655
rect 28944 6634 28970 6638
rect 30324 6655 30350 6660
rect 30324 6638 30328 6655
rect 30328 6638 30345 6655
rect 30345 6638 30350 6655
rect 30324 6634 30350 6638
rect 26644 6621 26670 6626
rect 26644 6604 26648 6621
rect 26648 6604 26665 6621
rect 26665 6604 26670 6621
rect 26644 6600 26670 6604
rect 27932 6621 27958 6626
rect 27334 6566 27360 6592
rect 27932 6604 27936 6621
rect 27936 6604 27953 6621
rect 27953 6604 27958 6621
rect 27932 6600 27958 6604
rect 28300 6600 28326 6626
rect 28668 6587 28694 6592
rect 28668 6570 28672 6587
rect 28672 6570 28689 6587
rect 28689 6570 28694 6587
rect 28668 6566 28694 6570
rect 28852 6600 28878 6626
rect 29312 6600 29338 6626
rect 30738 6600 30764 6626
rect 29818 6587 29844 6592
rect 29818 6570 29822 6587
rect 29822 6570 29839 6587
rect 29839 6570 29844 6587
rect 33084 6655 33110 6660
rect 33084 6638 33088 6655
rect 33088 6638 33105 6655
rect 33105 6638 33110 6655
rect 33084 6634 33110 6638
rect 34648 6655 34674 6660
rect 34648 6638 34652 6655
rect 34652 6638 34669 6655
rect 34669 6638 34674 6655
rect 34648 6634 34674 6638
rect 36350 6672 36354 6689
rect 36354 6672 36371 6689
rect 36371 6672 36376 6689
rect 36350 6668 36376 6672
rect 37684 6706 37688 6723
rect 37688 6706 37705 6723
rect 37705 6706 37710 6723
rect 37684 6702 37710 6706
rect 37822 6702 37848 6728
rect 40122 6689 40148 6694
rect 40122 6672 40126 6689
rect 40126 6672 40143 6689
rect 40143 6672 40148 6689
rect 40122 6668 40148 6672
rect 40812 6689 40838 6694
rect 40812 6672 40816 6689
rect 40816 6672 40833 6689
rect 40833 6672 40838 6689
rect 46930 6702 46956 6728
rect 40812 6668 40838 6672
rect 30876 6600 30902 6626
rect 29818 6566 29844 6570
rect 30830 6566 30856 6592
rect 32946 6566 32972 6592
rect 32992 6587 33018 6592
rect 32992 6570 32996 6587
rect 32996 6570 33013 6587
rect 33013 6570 33018 6587
rect 34556 6587 34582 6592
rect 32992 6566 33018 6570
rect 34556 6570 34560 6587
rect 34560 6570 34577 6587
rect 34577 6570 34582 6587
rect 34556 6566 34582 6570
rect 36166 6566 36192 6592
rect 36212 6587 36238 6592
rect 36212 6570 36216 6587
rect 36216 6570 36233 6587
rect 36233 6570 36238 6587
rect 36948 6621 36974 6626
rect 36948 6604 36952 6621
rect 36952 6604 36969 6621
rect 36969 6604 36974 6621
rect 36948 6600 36974 6604
rect 37592 6600 37618 6626
rect 39202 6634 39228 6660
rect 40720 6634 40746 6660
rect 41548 6655 41574 6660
rect 38236 6621 38262 6626
rect 38236 6604 38240 6621
rect 38240 6604 38257 6621
rect 38257 6604 38262 6621
rect 38236 6600 38262 6604
rect 39386 6621 39412 6626
rect 36212 6566 36238 6570
rect 38972 6587 38998 6592
rect 38972 6570 38976 6587
rect 38976 6570 38993 6587
rect 38993 6570 38998 6587
rect 39386 6604 39390 6621
rect 39390 6604 39407 6621
rect 39407 6604 39412 6621
rect 39386 6600 39412 6604
rect 39662 6600 39688 6626
rect 40030 6600 40056 6626
rect 41548 6638 41552 6655
rect 41552 6638 41569 6655
rect 41569 6638 41574 6655
rect 41548 6634 41574 6638
rect 41962 6655 41988 6660
rect 41962 6638 41966 6655
rect 41966 6638 41983 6655
rect 41983 6638 41988 6655
rect 41962 6634 41988 6638
rect 38972 6566 38998 6570
rect 40398 6566 40424 6592
rect 40720 6587 40746 6592
rect 40720 6570 40724 6587
rect 40724 6570 40741 6587
rect 40741 6570 40746 6587
rect 40720 6566 40746 6570
rect 41916 6600 41942 6626
rect 42238 6600 42264 6626
rect 42744 6600 42770 6626
rect 41456 6587 41482 6592
rect 41456 6570 41460 6587
rect 41460 6570 41477 6587
rect 41477 6570 41482 6587
rect 41456 6566 41482 6570
rect 41962 6566 41988 6592
rect 43020 6566 43046 6592
rect 43940 6634 43966 6660
rect 43388 6621 43414 6626
rect 43388 6604 43392 6621
rect 43392 6604 43409 6621
rect 43409 6604 43414 6621
rect 43388 6600 43414 6604
rect 44124 6587 44150 6592
rect 44124 6570 44128 6587
rect 44128 6570 44145 6587
rect 44145 6570 44150 6587
rect 44124 6566 44150 6570
rect 44538 6621 44564 6626
rect 44538 6604 44542 6621
rect 44542 6604 44559 6621
rect 44559 6604 44564 6621
rect 44538 6600 44564 6604
rect 44768 6600 44794 6626
rect 45826 6600 45852 6626
rect 45918 6621 45944 6626
rect 45918 6604 45922 6621
rect 45922 6604 45939 6621
rect 45939 6604 45944 6621
rect 45918 6600 45944 6604
rect 46010 6621 46036 6626
rect 46010 6604 46014 6621
rect 46014 6604 46031 6621
rect 46031 6604 46036 6621
rect 46010 6600 46036 6604
rect 45274 6587 45300 6592
rect 45274 6570 45278 6587
rect 45278 6570 45295 6587
rect 45295 6570 45300 6587
rect 49552 6668 49578 6694
rect 50380 6702 50406 6728
rect 54520 6702 54546 6728
rect 55854 6702 55880 6728
rect 59442 6702 59468 6728
rect 60638 6723 60664 6728
rect 59120 6668 59146 6694
rect 60638 6706 60642 6723
rect 60642 6706 60659 6723
rect 60659 6706 60664 6723
rect 60638 6702 60664 6706
rect 62064 6723 62090 6728
rect 62064 6706 62068 6723
rect 62068 6706 62085 6723
rect 62085 6706 62090 6723
rect 62064 6702 62090 6706
rect 63766 6702 63792 6728
rect 68320 6723 68346 6728
rect 68320 6706 68324 6723
rect 68324 6706 68341 6723
rect 68341 6706 68346 6723
rect 68320 6702 68346 6706
rect 69792 6702 69818 6728
rect 71448 6740 71452 6757
rect 71452 6740 71469 6757
rect 71469 6740 71474 6757
rect 71448 6736 71474 6740
rect 72874 6736 72900 6762
rect 74070 6736 74096 6762
rect 75404 6736 75430 6762
rect 48356 6587 48382 6592
rect 45274 6566 45300 6570
rect 48356 6570 48360 6587
rect 48360 6570 48377 6587
rect 48377 6570 48382 6587
rect 48356 6566 48382 6570
rect 48770 6587 48796 6592
rect 48770 6570 48774 6587
rect 48774 6570 48791 6587
rect 48791 6570 48796 6587
rect 48770 6566 48796 6570
rect 49000 6600 49026 6626
rect 49598 6600 49624 6626
rect 50702 6634 50728 6660
rect 49828 6621 49854 6626
rect 49828 6604 49832 6621
rect 49832 6604 49849 6621
rect 49849 6604 49854 6621
rect 49828 6600 49854 6604
rect 50472 6600 50498 6626
rect 50518 6566 50544 6592
rect 51668 6634 51694 6660
rect 52128 6655 52154 6660
rect 51116 6621 51142 6626
rect 51116 6604 51120 6621
rect 51120 6604 51137 6621
rect 51137 6604 51142 6621
rect 51116 6600 51142 6604
rect 52128 6638 52132 6655
rect 52132 6638 52149 6655
rect 52149 6638 52154 6655
rect 52128 6634 52154 6638
rect 54796 6655 54822 6660
rect 54796 6638 54800 6655
rect 54800 6638 54817 6655
rect 54817 6638 54822 6655
rect 54796 6634 54822 6638
rect 55716 6655 55742 6660
rect 55716 6638 55720 6655
rect 55720 6638 55737 6655
rect 55737 6638 55742 6655
rect 55716 6634 55742 6638
rect 57418 6655 57444 6660
rect 57418 6638 57422 6655
rect 57422 6638 57439 6655
rect 57439 6638 57444 6655
rect 57418 6634 57444 6638
rect 58706 6655 58732 6660
rect 58706 6638 58710 6655
rect 58710 6638 58727 6655
rect 58727 6638 58732 6655
rect 58706 6634 58732 6638
rect 59396 6634 59422 6660
rect 65146 6689 65172 6694
rect 65146 6672 65150 6689
rect 65150 6672 65167 6689
rect 65167 6672 65172 6689
rect 65146 6668 65172 6672
rect 71034 6668 71060 6694
rect 52036 6600 52062 6626
rect 52496 6600 52522 6626
rect 56268 6621 56294 6626
rect 56268 6604 56272 6621
rect 56272 6604 56289 6621
rect 56289 6604 56294 6621
rect 56268 6600 56294 6604
rect 57096 6600 57122 6626
rect 57556 6621 57582 6626
rect 57556 6604 57560 6621
rect 57560 6604 57577 6621
rect 57577 6604 57582 6621
rect 57556 6600 57582 6604
rect 58476 6600 58502 6626
rect 58844 6621 58870 6626
rect 58844 6604 58848 6621
rect 58848 6604 58865 6621
rect 58865 6604 58870 6621
rect 58844 6600 58870 6604
rect 51852 6587 51878 6592
rect 51852 6570 51856 6587
rect 51856 6570 51873 6587
rect 51873 6570 51878 6587
rect 51852 6566 51878 6570
rect 52220 6566 52246 6592
rect 52312 6566 52338 6592
rect 54796 6566 54822 6592
rect 57280 6566 57306 6592
rect 57464 6566 57490 6592
rect 57878 6566 57904 6592
rect 59028 6566 59054 6592
rect 63766 6655 63792 6660
rect 63766 6638 63770 6655
rect 63770 6638 63787 6655
rect 63787 6638 63792 6655
rect 63766 6634 63792 6638
rect 64686 6634 64712 6660
rect 68412 6655 68438 6660
rect 68412 6638 68416 6655
rect 68416 6638 68433 6655
rect 68433 6638 68438 6655
rect 68412 6634 68438 6638
rect 71540 6655 71566 6660
rect 62754 6621 62780 6626
rect 62754 6604 62758 6621
rect 62758 6604 62775 6621
rect 62775 6604 62780 6621
rect 62754 6600 62780 6604
rect 63904 6621 63930 6626
rect 63904 6604 63908 6621
rect 63908 6604 63925 6621
rect 63925 6604 63930 6621
rect 63904 6600 63930 6604
rect 59856 6587 59882 6592
rect 59856 6570 59860 6587
rect 59860 6570 59877 6587
rect 59877 6570 59882 6587
rect 59856 6566 59882 6570
rect 63076 6587 63102 6592
rect 63076 6570 63080 6587
rect 63080 6570 63097 6587
rect 63097 6570 63102 6587
rect 63076 6566 63102 6570
rect 63260 6587 63286 6592
rect 63260 6570 63264 6587
rect 63264 6570 63281 6587
rect 63281 6570 63286 6587
rect 63260 6566 63286 6570
rect 64042 6566 64068 6592
rect 65606 6600 65632 6626
rect 66434 6621 66460 6626
rect 66434 6604 66438 6621
rect 66438 6604 66455 6621
rect 66455 6604 66460 6621
rect 66434 6600 66460 6604
rect 66664 6600 66690 6626
rect 71540 6638 71544 6655
rect 71544 6638 71561 6655
rect 71561 6638 71566 6655
rect 71540 6634 71566 6638
rect 72874 6655 72900 6660
rect 72874 6638 72878 6655
rect 72878 6638 72895 6655
rect 72895 6638 72900 6655
rect 72874 6634 72900 6638
rect 78624 6736 78650 6762
rect 78992 6736 79018 6762
rect 79728 6736 79754 6762
rect 80786 6736 80812 6762
rect 81338 6736 81364 6762
rect 81752 6736 81778 6762
rect 88192 6736 88218 6762
rect 91366 6757 91392 6762
rect 77474 6702 77500 6728
rect 83224 6702 83250 6728
rect 85202 6723 85228 6728
rect 80464 6689 80490 6694
rect 80464 6672 80468 6689
rect 80468 6672 80485 6689
rect 80485 6672 80490 6689
rect 80464 6668 80490 6672
rect 82626 6668 82652 6694
rect 64594 6566 64620 6592
rect 65790 6566 65816 6592
rect 66848 6566 66874 6592
rect 67078 6566 67104 6592
rect 72966 6600 72992 6626
rect 73012 6621 73038 6626
rect 73012 6604 73016 6621
rect 73016 6604 73033 6621
rect 73033 6604 73038 6621
rect 73012 6600 73038 6604
rect 73794 6600 73820 6626
rect 72920 6566 72946 6592
rect 73748 6587 73774 6592
rect 73748 6570 73752 6587
rect 73752 6570 73769 6587
rect 73769 6570 73774 6587
rect 73748 6566 73774 6570
rect 77612 6634 77638 6660
rect 77934 6634 77960 6660
rect 78210 6655 78236 6660
rect 78210 6638 78214 6655
rect 78214 6638 78231 6655
rect 78231 6638 78236 6655
rect 78210 6634 78236 6638
rect 78900 6655 78926 6660
rect 78900 6638 78904 6655
rect 78904 6638 78921 6655
rect 78921 6638 78926 6655
rect 78900 6634 78926 6638
rect 79314 6655 79340 6660
rect 79314 6638 79318 6655
rect 79318 6638 79335 6655
rect 79335 6638 79340 6655
rect 79314 6634 79340 6638
rect 81338 6634 81364 6660
rect 81752 6655 81778 6660
rect 74622 6566 74648 6592
rect 75220 6600 75246 6626
rect 75542 6600 75568 6626
rect 76232 6600 76258 6626
rect 76876 6621 76902 6626
rect 76324 6587 76350 6592
rect 76324 6570 76328 6587
rect 76328 6570 76345 6587
rect 76345 6570 76350 6587
rect 76876 6604 76880 6621
rect 76880 6604 76897 6621
rect 76897 6604 76902 6621
rect 76876 6600 76902 6604
rect 77106 6600 77132 6626
rect 78302 6600 78328 6626
rect 79452 6621 79478 6626
rect 77612 6587 77638 6592
rect 76324 6566 76350 6570
rect 77612 6570 77616 6587
rect 77616 6570 77633 6587
rect 77633 6570 77638 6587
rect 77612 6566 77638 6570
rect 79452 6604 79456 6621
rect 79456 6604 79473 6621
rect 79473 6604 79478 6621
rect 79452 6600 79478 6604
rect 80602 6621 80628 6626
rect 79774 6566 79800 6592
rect 80188 6587 80214 6592
rect 80188 6570 80192 6587
rect 80192 6570 80209 6587
rect 80209 6570 80214 6587
rect 80188 6566 80214 6570
rect 80602 6604 80606 6621
rect 80606 6604 80623 6621
rect 80623 6604 80628 6621
rect 80602 6600 80628 6604
rect 81384 6600 81410 6626
rect 81016 6566 81042 6592
rect 81246 6566 81272 6592
rect 81752 6638 81756 6655
rect 81756 6638 81773 6655
rect 81773 6638 81778 6655
rect 81752 6634 81778 6638
rect 82442 6634 82468 6660
rect 85202 6706 85206 6723
rect 85206 6706 85223 6723
rect 85223 6706 85228 6723
rect 85202 6702 85228 6706
rect 86536 6723 86562 6728
rect 86536 6706 86540 6723
rect 86540 6706 86557 6723
rect 86557 6706 86562 6723
rect 86536 6702 86562 6706
rect 86904 6723 86930 6728
rect 86904 6706 86908 6723
rect 86908 6706 86925 6723
rect 86925 6706 86930 6723
rect 86904 6702 86930 6706
rect 87962 6702 87988 6728
rect 88008 6702 88034 6728
rect 88882 6702 88908 6728
rect 90216 6702 90242 6728
rect 81890 6621 81916 6626
rect 81890 6604 81894 6621
rect 81894 6604 81911 6621
rect 81911 6604 81916 6621
rect 81890 6600 81916 6604
rect 82304 6566 82330 6592
rect 82580 6600 82606 6626
rect 83684 6621 83710 6626
rect 83684 6604 83688 6621
rect 83688 6604 83705 6621
rect 83705 6604 83710 6621
rect 83684 6600 83710 6604
rect 87088 6655 87114 6660
rect 87088 6638 87092 6655
rect 87092 6638 87109 6655
rect 87109 6638 87114 6655
rect 87088 6634 87114 6638
rect 82626 6587 82652 6592
rect 82626 6570 82630 6587
rect 82630 6570 82647 6587
rect 82647 6570 82652 6587
rect 82626 6566 82652 6570
rect 82672 6566 82698 6592
rect 83224 6587 83250 6592
rect 83224 6570 83228 6587
rect 83228 6570 83245 6587
rect 83245 6570 83250 6587
rect 83224 6566 83250 6570
rect 87916 6634 87942 6660
rect 90952 6668 90978 6694
rect 91044 6689 91070 6694
rect 91044 6672 91048 6689
rect 91048 6672 91065 6689
rect 91065 6672 91070 6689
rect 91366 6740 91370 6757
rect 91370 6740 91387 6757
rect 91387 6740 91392 6757
rect 91366 6736 91392 6740
rect 92884 6757 92910 6762
rect 92884 6740 92888 6757
rect 92888 6740 92905 6757
rect 92905 6740 92910 6757
rect 92884 6736 92910 6740
rect 94678 6736 94704 6762
rect 94402 6702 94428 6728
rect 94770 6702 94796 6728
rect 95460 6736 95486 6762
rect 96748 6736 96774 6762
rect 94264 6689 94290 6694
rect 91044 6668 91070 6672
rect 88192 6655 88218 6660
rect 88192 6638 88196 6655
rect 88196 6638 88213 6655
rect 88213 6638 88218 6655
rect 88192 6634 88218 6638
rect 90308 6634 90334 6660
rect 94264 6672 94268 6689
rect 94268 6672 94285 6689
rect 94285 6672 94290 6689
rect 94264 6668 94290 6672
rect 95920 6702 95946 6728
rect 103556 6736 103582 6762
rect 105166 6757 105192 6762
rect 94954 6668 94980 6694
rect 100980 6702 101006 6728
rect 101716 6702 101742 6728
rect 103004 6702 103030 6728
rect 103878 6702 103904 6728
rect 98818 6668 98844 6694
rect 101026 6668 101052 6694
rect 94770 6655 94796 6660
rect 87870 6600 87896 6626
rect 88836 6600 88862 6626
rect 87502 6566 87528 6592
rect 89986 6600 90012 6626
rect 90446 6600 90472 6626
rect 90354 6587 90380 6592
rect 90354 6570 90358 6587
rect 90358 6570 90375 6587
rect 90375 6570 90380 6587
rect 90354 6566 90380 6570
rect 94770 6638 94774 6655
rect 94774 6638 94791 6655
rect 94791 6638 94796 6655
rect 94770 6634 94796 6638
rect 93896 6566 93922 6592
rect 93988 6587 94014 6592
rect 93988 6570 93992 6587
rect 93992 6570 94009 6587
rect 94009 6570 94014 6587
rect 93988 6566 94014 6570
rect 94172 6587 94198 6592
rect 94172 6570 94176 6587
rect 94176 6570 94193 6587
rect 94193 6570 94198 6587
rect 94172 6566 94198 6570
rect 94770 6566 94796 6592
rect 95690 6566 95716 6592
rect 96196 6600 96222 6626
rect 96702 6600 96728 6626
rect 96978 6600 97004 6626
rect 100750 6634 100776 6660
rect 101072 6655 101098 6660
rect 101072 6638 101076 6655
rect 101076 6638 101093 6655
rect 101093 6638 101098 6655
rect 101072 6634 101098 6638
rect 97300 6600 97326 6626
rect 97392 6600 97418 6626
rect 98220 6621 98246 6626
rect 98220 6604 98224 6621
rect 98224 6604 98241 6621
rect 98241 6604 98246 6621
rect 98220 6600 98246 6604
rect 98680 6600 98706 6626
rect 101210 6621 101236 6626
rect 98864 6566 98890 6592
rect 98956 6566 98982 6592
rect 99278 6587 99304 6592
rect 99278 6570 99282 6587
rect 99282 6570 99299 6587
rect 99299 6570 99304 6587
rect 99278 6566 99304 6570
rect 100244 6587 100270 6592
rect 100244 6570 100248 6587
rect 100248 6570 100265 6587
rect 100265 6570 100270 6587
rect 100244 6566 100270 6570
rect 100428 6587 100454 6592
rect 100428 6570 100432 6587
rect 100432 6570 100449 6587
rect 100449 6570 100454 6587
rect 100428 6566 100454 6570
rect 100658 6566 100684 6592
rect 101210 6604 101214 6621
rect 101214 6604 101231 6621
rect 101231 6604 101236 6621
rect 101210 6600 101236 6604
rect 101578 6600 101604 6626
rect 102130 6600 102156 6626
rect 102728 6600 102754 6626
rect 102820 6566 102846 6592
rect 102866 6566 102892 6592
rect 103602 6634 103628 6660
rect 103188 6600 103214 6626
rect 103786 6600 103812 6626
rect 105166 6740 105170 6757
rect 105170 6740 105187 6757
rect 105187 6740 105192 6757
rect 105166 6736 105192 6740
rect 106684 6757 106710 6762
rect 106684 6740 106688 6757
rect 106688 6740 106705 6757
rect 106705 6740 106710 6757
rect 106684 6736 106710 6740
rect 104016 6702 104042 6728
rect 106638 6702 106664 6728
rect 134468 6736 134494 6762
rect 134790 6736 134816 6762
rect 135894 6736 135920 6762
rect 137458 6757 137484 6762
rect 137458 6740 137462 6757
rect 137462 6740 137479 6757
rect 137479 6740 137484 6757
rect 137458 6736 137484 6740
rect 138930 6757 138956 6762
rect 138930 6740 138934 6757
rect 138934 6740 138951 6757
rect 138951 6740 138956 6757
rect 138930 6736 138956 6740
rect 140448 6757 140474 6762
rect 140448 6740 140452 6757
rect 140452 6740 140469 6757
rect 140469 6740 140474 6757
rect 140448 6736 140474 6740
rect 142150 6736 142176 6762
rect 143530 6736 143556 6762
rect 145048 6757 145074 6762
rect 145048 6740 145052 6757
rect 145052 6740 145069 6757
rect 145069 6740 145074 6757
rect 145048 6736 145074 6740
rect 146612 6757 146638 6762
rect 146612 6740 146616 6757
rect 146616 6740 146633 6757
rect 146633 6740 146638 6757
rect 146612 6736 146638 6740
rect 148130 6757 148156 6762
rect 148130 6740 148134 6757
rect 148134 6740 148151 6757
rect 148151 6740 148156 6757
rect 148130 6736 148156 6740
rect 149648 6757 149674 6762
rect 149648 6740 149652 6757
rect 149652 6740 149669 6757
rect 149669 6740 149674 6757
rect 149648 6736 149674 6740
rect 150706 6757 150732 6762
rect 150706 6740 150710 6757
rect 150710 6740 150727 6757
rect 150727 6740 150732 6757
rect 150706 6736 150732 6740
rect 108202 6723 108228 6728
rect 108202 6706 108206 6723
rect 108206 6706 108223 6723
rect 108223 6706 108228 6723
rect 108202 6702 108228 6706
rect 109720 6702 109746 6728
rect 103970 6634 103996 6660
rect 106776 6655 106802 6660
rect 106776 6638 106780 6655
rect 106780 6638 106797 6655
rect 106797 6638 106802 6655
rect 106776 6634 106802 6638
rect 108294 6655 108320 6660
rect 108294 6638 108298 6655
rect 108298 6638 108315 6655
rect 108315 6638 108320 6655
rect 112066 6702 112092 6728
rect 112020 6668 112046 6694
rect 113216 6702 113242 6728
rect 113308 6723 113334 6728
rect 113308 6706 113312 6723
rect 113312 6706 113329 6723
rect 113329 6706 113334 6723
rect 113308 6702 113334 6706
rect 113446 6702 113472 6728
rect 113952 6702 113978 6728
rect 114596 6702 114622 6728
rect 112204 6668 112230 6694
rect 113538 6689 113564 6694
rect 113538 6672 113542 6689
rect 113542 6672 113559 6689
rect 113559 6672 113564 6689
rect 113538 6668 113564 6672
rect 113584 6689 113610 6694
rect 113584 6672 113588 6689
rect 113588 6672 113605 6689
rect 113605 6672 113610 6689
rect 113584 6668 113610 6672
rect 108294 6634 108320 6638
rect 112112 6600 112138 6626
rect 103694 6566 103720 6592
rect 106776 6566 106802 6592
rect 111376 6587 111402 6592
rect 111376 6570 111380 6587
rect 111380 6570 111397 6587
rect 111397 6570 111402 6587
rect 111376 6566 111402 6570
rect 111836 6587 111862 6592
rect 111836 6570 111840 6587
rect 111840 6570 111857 6587
rect 111857 6570 111862 6587
rect 111836 6566 111862 6570
rect 112020 6587 112046 6592
rect 112020 6570 112024 6587
rect 112024 6570 112041 6587
rect 112041 6570 112046 6587
rect 112020 6566 112046 6570
rect 112066 6587 112092 6592
rect 112066 6570 112070 6587
rect 112070 6570 112087 6587
rect 112087 6570 112092 6587
rect 112204 6600 112230 6626
rect 113860 6634 113886 6660
rect 115976 6668 116002 6694
rect 115194 6634 115220 6660
rect 115930 6634 115956 6660
rect 116022 6634 116048 6660
rect 116574 6668 116600 6694
rect 116666 6668 116692 6694
rect 116528 6655 116554 6660
rect 116528 6638 116532 6655
rect 116532 6638 116549 6655
rect 116549 6638 116554 6655
rect 116528 6634 116554 6638
rect 114044 6600 114070 6626
rect 115378 6621 115404 6626
rect 115378 6604 115382 6621
rect 115382 6604 115399 6621
rect 115399 6604 115404 6621
rect 115378 6600 115404 6604
rect 118966 6668 118992 6694
rect 119058 6668 119084 6694
rect 119748 6702 119774 6728
rect 122324 6702 122350 6728
rect 122692 6702 122718 6728
rect 123566 6723 123592 6728
rect 123566 6706 123570 6723
rect 123570 6706 123587 6723
rect 123587 6706 123592 6723
rect 123566 6702 123592 6706
rect 125544 6702 125570 6728
rect 126234 6702 126260 6728
rect 127476 6702 127502 6728
rect 129730 6723 129756 6728
rect 129730 6706 129734 6723
rect 129734 6706 129751 6723
rect 129751 6706 129756 6723
rect 129730 6702 129756 6706
rect 131754 6702 131780 6728
rect 132766 6702 132792 6728
rect 135204 6702 135230 6728
rect 122048 6668 122074 6694
rect 119104 6655 119130 6660
rect 119104 6638 119108 6655
rect 119108 6638 119125 6655
rect 119125 6638 119130 6655
rect 119104 6634 119130 6638
rect 119886 6634 119912 6660
rect 125498 6668 125524 6694
rect 125544 6655 125570 6660
rect 125544 6638 125548 6655
rect 125548 6638 125565 6655
rect 125565 6638 125570 6655
rect 125544 6634 125570 6638
rect 112066 6566 112092 6570
rect 112710 6566 112736 6592
rect 112848 6587 112874 6592
rect 112848 6570 112852 6587
rect 112852 6570 112869 6587
rect 112869 6570 112874 6587
rect 112848 6566 112874 6570
rect 113538 6566 113564 6592
rect 113814 6566 113840 6592
rect 113952 6566 113978 6592
rect 116068 6566 116094 6592
rect 116620 6566 116646 6592
rect 117448 6587 117474 6592
rect 117448 6570 117452 6587
rect 117452 6570 117469 6587
rect 117469 6570 117474 6587
rect 117448 6566 117474 6570
rect 118506 6566 118532 6592
rect 119242 6621 119268 6626
rect 119242 6604 119246 6621
rect 119246 6604 119263 6621
rect 119263 6604 119268 6621
rect 120530 6621 120556 6626
rect 119242 6600 119268 6604
rect 120530 6604 120534 6621
rect 120534 6604 120551 6621
rect 120551 6604 120556 6621
rect 120530 6600 120556 6604
rect 120898 6600 120924 6626
rect 121818 6621 121844 6626
rect 121266 6587 121292 6592
rect 121266 6570 121270 6587
rect 121270 6570 121287 6587
rect 121287 6570 121292 6587
rect 121266 6566 121292 6570
rect 121818 6604 121822 6621
rect 121822 6604 121839 6621
rect 121839 6604 121844 6621
rect 121818 6600 121844 6604
rect 122462 6600 122488 6626
rect 125590 6566 125616 6592
rect 125682 6621 125708 6626
rect 125682 6604 125686 6621
rect 125686 6604 125703 6621
rect 125703 6604 125708 6621
rect 125682 6600 125708 6604
rect 126188 6600 126214 6626
rect 128120 6655 128146 6660
rect 126510 6600 126536 6626
rect 127476 6600 127502 6626
rect 126740 6566 126766 6592
rect 128120 6638 128124 6655
rect 128124 6638 128141 6655
rect 128141 6638 128146 6655
rect 128120 6634 128146 6638
rect 127660 6600 127686 6626
rect 128488 6600 128514 6626
rect 128166 6566 128192 6592
rect 132076 6668 132102 6694
rect 136492 6702 136518 6728
rect 134468 6634 134494 6660
rect 136584 6668 136610 6694
rect 136630 6634 136656 6660
rect 137550 6655 137576 6660
rect 137550 6638 137554 6655
rect 137554 6638 137571 6655
rect 137571 6638 137576 6655
rect 137550 6634 137576 6638
rect 130926 6621 130952 6626
rect 130926 6604 130930 6621
rect 130930 6604 130947 6621
rect 130947 6604 130952 6621
rect 130926 6600 130952 6604
rect 131708 6600 131734 6626
rect 131754 6600 131780 6626
rect 132214 6600 132240 6626
rect 132306 6600 132332 6626
rect 132490 6600 132516 6626
rect 128994 6587 129020 6592
rect 128994 6570 128998 6587
rect 128998 6570 129015 6587
rect 129015 6570 129020 6587
rect 128994 6566 129020 6570
rect 131478 6566 131504 6592
rect 131662 6566 131688 6592
rect 133456 6600 133482 6626
rect 133824 6566 133850 6592
rect 134376 6600 134402 6626
rect 135342 6600 135368 6626
rect 135388 6566 135414 6592
rect 135480 6600 135506 6626
rect 140540 6655 140566 6660
rect 140540 6638 140544 6655
rect 140544 6638 140561 6655
rect 140561 6638 140566 6655
rect 140540 6634 140566 6638
rect 142380 6655 142406 6660
rect 142380 6638 142384 6655
rect 142384 6638 142401 6655
rect 142401 6638 142406 6655
rect 142380 6634 142406 6638
rect 145140 6655 145166 6660
rect 145140 6638 145144 6655
rect 145144 6638 145161 6655
rect 145161 6638 145166 6655
rect 145140 6634 145166 6638
rect 152500 6668 152526 6694
rect 135894 6566 135920 6592
rect 136446 6566 136472 6592
rect 149740 6655 149766 6660
rect 149740 6638 149744 6655
rect 149744 6638 149761 6655
rect 149761 6638 149766 6655
rect 149740 6634 149766 6638
rect 151764 6634 151790 6660
rect 147946 6587 147972 6592
rect 147946 6570 147950 6587
rect 147950 6570 147967 6587
rect 147967 6570 147972 6587
rect 147946 6566 147972 6570
rect 38574 6515 38600 6541
rect 38606 6515 38632 6541
rect 38638 6515 38664 6541
rect 38670 6515 38696 6541
rect 38702 6515 38728 6541
rect 76673 6515 76699 6541
rect 76705 6515 76731 6541
rect 76737 6515 76763 6541
rect 76769 6515 76795 6541
rect 76801 6515 76827 6541
rect 114772 6515 114798 6541
rect 114804 6515 114830 6541
rect 114836 6515 114862 6541
rect 114868 6515 114894 6541
rect 114900 6515 114926 6541
rect 13028 6485 13054 6490
rect 13028 6468 13032 6485
rect 13032 6468 13049 6485
rect 13049 6468 13054 6485
rect 13028 6464 13054 6468
rect 10084 6430 10110 6456
rect 13672 6430 13698 6456
rect 16110 6464 16136 6490
rect 17076 6464 17102 6490
rect 17766 6485 17792 6490
rect 17766 6468 17770 6485
rect 17770 6468 17787 6485
rect 17787 6468 17792 6485
rect 17766 6464 17792 6468
rect 14500 6451 14526 6456
rect 11602 6362 11628 6388
rect 14500 6434 14504 6451
rect 14504 6434 14521 6451
rect 14521 6434 14526 6451
rect 14500 6430 14526 6434
rect 13994 6396 14020 6422
rect 14040 6383 14066 6388
rect 13580 6328 13606 6354
rect 14040 6366 14044 6383
rect 14044 6366 14061 6383
rect 14061 6366 14066 6383
rect 14040 6362 14066 6366
rect 15190 6430 15216 6456
rect 15788 6430 15814 6456
rect 17214 6430 17240 6456
rect 16846 6396 16872 6422
rect 18732 6430 18758 6456
rect 19836 6430 19862 6456
rect 20526 6430 20552 6456
rect 21630 6464 21656 6490
rect 22136 6464 22162 6490
rect 22274 6485 22300 6490
rect 22274 6468 22278 6485
rect 22278 6468 22295 6485
rect 22295 6468 22300 6485
rect 22274 6464 22300 6468
rect 26644 6464 26670 6490
rect 21492 6430 21518 6456
rect 27334 6464 27360 6490
rect 27932 6464 27958 6490
rect 28990 6464 29016 6490
rect 29818 6464 29844 6490
rect 36074 6485 36100 6490
rect 36074 6468 36078 6485
rect 36078 6468 36095 6485
rect 36095 6468 36100 6485
rect 36074 6464 36100 6468
rect 36166 6464 36192 6490
rect 37362 6464 37388 6490
rect 14822 6362 14848 6388
rect 14914 6383 14940 6388
rect 14914 6366 14918 6383
rect 14918 6366 14935 6383
rect 14935 6366 14940 6383
rect 14914 6362 14940 6366
rect 15052 6383 15078 6388
rect 15052 6366 15056 6383
rect 15056 6366 15073 6383
rect 15073 6366 15078 6383
rect 15052 6362 15078 6366
rect 14454 6294 14480 6320
rect 16524 6362 16550 6388
rect 16708 6362 16734 6388
rect 17168 6362 17194 6388
rect 19652 6396 19678 6422
rect 20756 6396 20782 6422
rect 17444 6383 17470 6388
rect 17444 6366 17448 6383
rect 17448 6366 17465 6383
rect 17465 6366 17470 6383
rect 17444 6362 17470 6366
rect 17674 6362 17700 6388
rect 19698 6362 19724 6388
rect 20480 6362 20506 6388
rect 21538 6362 21564 6388
rect 21584 6362 21610 6388
rect 22688 6396 22714 6422
rect 27748 6430 27774 6456
rect 28668 6430 28694 6456
rect 30324 6430 30350 6456
rect 32946 6430 32972 6456
rect 26874 6396 26900 6422
rect 27012 6417 27038 6422
rect 21906 6362 21932 6388
rect 22734 6362 22760 6388
rect 25678 6362 25704 6388
rect 27012 6400 27016 6417
rect 27016 6400 27033 6417
rect 27033 6400 27038 6417
rect 27012 6396 27038 6400
rect 27380 6417 27406 6422
rect 27058 6383 27084 6388
rect 27058 6366 27062 6383
rect 27062 6366 27079 6383
rect 27079 6366 27084 6383
rect 27058 6362 27084 6366
rect 27380 6400 27384 6417
rect 27384 6400 27401 6417
rect 27401 6400 27406 6417
rect 27380 6396 27406 6400
rect 28714 6396 28740 6422
rect 37408 6396 37434 6422
rect 37730 6396 37756 6422
rect 39202 6430 39228 6456
rect 39846 6396 39872 6422
rect 41962 6464 41988 6490
rect 40260 6430 40286 6456
rect 41456 6430 41482 6456
rect 43250 6464 43276 6490
rect 43572 6464 43598 6490
rect 45228 6464 45254 6490
rect 45826 6464 45852 6490
rect 49000 6464 49026 6490
rect 27518 6383 27544 6388
rect 27518 6366 27522 6383
rect 27522 6366 27539 6383
rect 27539 6366 27544 6383
rect 27518 6362 27544 6366
rect 39294 6362 39320 6388
rect 15696 6294 15722 6320
rect 16202 6294 16228 6320
rect 17076 6294 17102 6320
rect 19008 6315 19034 6320
rect 19008 6298 19012 6315
rect 19012 6298 19029 6315
rect 19029 6298 19034 6315
rect 19008 6294 19034 6298
rect 20618 6315 20644 6320
rect 20618 6298 20622 6315
rect 20622 6298 20639 6315
rect 20639 6298 20644 6315
rect 20618 6294 20644 6298
rect 20894 6315 20920 6320
rect 20894 6298 20898 6315
rect 20898 6298 20915 6315
rect 20915 6298 20920 6315
rect 20894 6294 20920 6298
rect 21400 6294 21426 6320
rect 21630 6294 21656 6320
rect 21906 6294 21932 6320
rect 26552 6294 26578 6320
rect 27058 6294 27084 6320
rect 27794 6294 27820 6320
rect 28162 6294 28188 6320
rect 28254 6315 28280 6320
rect 28254 6298 28258 6315
rect 28258 6298 28275 6315
rect 28275 6298 28280 6315
rect 28254 6294 28280 6298
rect 28622 6294 28648 6320
rect 36350 6294 36376 6320
rect 37500 6294 37526 6320
rect 37592 6294 37618 6320
rect 38926 6328 38952 6354
rect 39064 6328 39090 6354
rect 40398 6362 40424 6388
rect 38604 6294 38630 6320
rect 40720 6328 40746 6354
rect 40812 6294 40838 6320
rect 42422 6362 42448 6388
rect 42882 6315 42908 6320
rect 42882 6298 42886 6315
rect 42886 6298 42903 6315
rect 42903 6298 42908 6315
rect 42882 6294 42908 6298
rect 45274 6430 45300 6456
rect 45366 6430 45392 6456
rect 49736 6451 49762 6456
rect 49736 6434 49740 6451
rect 49740 6434 49757 6451
rect 49757 6434 49762 6451
rect 49736 6430 49762 6434
rect 49966 6430 49992 6456
rect 52312 6451 52338 6456
rect 52312 6434 52316 6451
rect 52316 6434 52333 6451
rect 52333 6434 52338 6451
rect 52312 6430 52338 6434
rect 52358 6451 52384 6456
rect 52358 6434 52362 6451
rect 52362 6434 52379 6451
rect 52379 6434 52384 6451
rect 52358 6430 52384 6434
rect 45090 6396 45116 6422
rect 45228 6417 45254 6422
rect 45228 6400 45232 6417
rect 45232 6400 45249 6417
rect 45249 6400 45254 6417
rect 45228 6396 45254 6400
rect 45320 6396 45346 6422
rect 43250 6383 43276 6388
rect 43250 6366 43254 6383
rect 43254 6366 43271 6383
rect 43271 6366 43276 6383
rect 43250 6362 43276 6366
rect 44124 6362 44150 6388
rect 44860 6362 44886 6388
rect 45044 6362 45070 6388
rect 52588 6396 52614 6422
rect 49598 6383 49624 6388
rect 49598 6366 49602 6383
rect 49602 6366 49619 6383
rect 49619 6366 49624 6383
rect 50702 6383 50728 6388
rect 49598 6362 49624 6366
rect 50702 6366 50706 6383
rect 50706 6366 50723 6383
rect 50723 6366 50728 6383
rect 50702 6362 50728 6366
rect 50840 6383 50866 6388
rect 50840 6366 50844 6383
rect 50844 6366 50861 6383
rect 50861 6366 50866 6383
rect 50840 6362 50866 6366
rect 43894 6294 43920 6320
rect 43986 6315 44012 6320
rect 43986 6298 43990 6315
rect 43990 6298 44007 6315
rect 44007 6298 44012 6315
rect 43986 6294 44012 6298
rect 44216 6294 44242 6320
rect 44952 6294 44978 6320
rect 49598 6294 49624 6320
rect 50518 6328 50544 6354
rect 51622 6328 51648 6354
rect 52956 6349 52982 6354
rect 52956 6332 52960 6349
rect 52960 6332 52977 6349
rect 52977 6332 52982 6349
rect 52956 6328 52982 6332
rect 55716 6464 55742 6490
rect 57280 6464 57306 6490
rect 57372 6464 57398 6490
rect 58706 6464 58732 6490
rect 59120 6485 59146 6490
rect 59120 6468 59124 6485
rect 59124 6468 59141 6485
rect 59141 6468 59146 6485
rect 59120 6464 59146 6468
rect 59350 6485 59376 6490
rect 59350 6468 59354 6485
rect 59354 6468 59371 6485
rect 59371 6468 59376 6485
rect 59350 6464 59376 6468
rect 63444 6464 63470 6490
rect 64042 6485 64068 6490
rect 64042 6468 64046 6485
rect 64046 6468 64063 6485
rect 64063 6468 64068 6485
rect 64042 6464 64068 6468
rect 64318 6464 64344 6490
rect 64594 6485 64620 6490
rect 64594 6468 64598 6485
rect 64598 6468 64615 6485
rect 64615 6468 64620 6485
rect 64594 6464 64620 6468
rect 66664 6464 66690 6490
rect 54796 6430 54822 6456
rect 56544 6417 56570 6422
rect 56544 6400 56548 6417
rect 56548 6400 56565 6417
rect 56565 6400 56570 6417
rect 56544 6396 56570 6400
rect 56912 6417 56938 6422
rect 56912 6400 56916 6417
rect 56916 6400 56933 6417
rect 56933 6400 56938 6417
rect 56912 6396 56938 6400
rect 57326 6417 57352 6422
rect 57326 6400 57330 6417
rect 57330 6400 57347 6417
rect 57347 6400 57352 6417
rect 57878 6430 57904 6456
rect 58660 6430 58686 6456
rect 63260 6430 63286 6456
rect 57326 6396 57352 6400
rect 59028 6396 59054 6422
rect 66204 6430 66230 6456
rect 66802 6451 66828 6456
rect 66802 6434 66806 6451
rect 66806 6434 66823 6451
rect 66823 6434 66828 6451
rect 66802 6430 66828 6434
rect 66940 6464 66966 6490
rect 73840 6464 73866 6490
rect 67078 6430 67104 6456
rect 71540 6430 71566 6456
rect 72966 6451 72992 6456
rect 63720 6417 63746 6422
rect 63720 6400 63724 6417
rect 63724 6400 63741 6417
rect 63741 6400 63746 6417
rect 63720 6396 63746 6400
rect 56958 6362 56984 6388
rect 57372 6362 57398 6388
rect 57832 6362 57858 6388
rect 57924 6383 57950 6388
rect 57924 6366 57928 6383
rect 57928 6366 57945 6383
rect 57945 6366 57950 6383
rect 57924 6362 57950 6366
rect 58384 6383 58410 6388
rect 57418 6328 57444 6354
rect 58384 6366 58388 6383
rect 58388 6366 58405 6383
rect 58405 6366 58410 6383
rect 58384 6362 58410 6366
rect 50380 6294 50406 6320
rect 51530 6294 51556 6320
rect 51806 6294 51832 6320
rect 55946 6315 55972 6320
rect 55946 6298 55950 6315
rect 55950 6298 55967 6315
rect 55967 6298 55972 6315
rect 55946 6294 55972 6298
rect 56544 6294 56570 6320
rect 57372 6315 57398 6320
rect 57372 6298 57376 6315
rect 57376 6298 57393 6315
rect 57393 6298 57398 6315
rect 57372 6294 57398 6298
rect 57924 6294 57950 6320
rect 63766 6362 63792 6388
rect 64042 6294 64068 6320
rect 64548 6417 64574 6422
rect 64548 6400 64552 6417
rect 64552 6400 64569 6417
rect 64569 6400 64574 6417
rect 64548 6396 64574 6400
rect 64180 6362 64206 6388
rect 65146 6396 65172 6422
rect 64870 6362 64896 6388
rect 65560 6383 65586 6388
rect 65560 6366 65564 6383
rect 65564 6366 65581 6383
rect 65581 6366 65586 6383
rect 65560 6362 65586 6366
rect 66296 6383 66322 6388
rect 66296 6366 66300 6383
rect 66300 6366 66317 6383
rect 66317 6366 66322 6383
rect 66848 6396 66874 6422
rect 72966 6434 72970 6451
rect 72970 6434 72987 6451
rect 72987 6434 72992 6451
rect 72966 6430 72992 6434
rect 76324 6464 76350 6490
rect 76416 6464 76442 6490
rect 78578 6485 78604 6490
rect 78578 6468 78582 6485
rect 78582 6468 78599 6485
rect 78599 6468 78604 6485
rect 78578 6464 78604 6468
rect 79314 6464 79340 6490
rect 72920 6417 72946 6422
rect 66296 6362 66322 6366
rect 71632 6383 71658 6388
rect 65146 6328 65172 6354
rect 66848 6328 66874 6354
rect 66572 6315 66598 6320
rect 66572 6298 66576 6315
rect 66576 6298 66593 6315
rect 66593 6298 66598 6315
rect 66572 6294 66598 6298
rect 66618 6294 66644 6320
rect 71632 6366 71636 6383
rect 71636 6366 71653 6383
rect 71653 6366 71658 6383
rect 71632 6362 71658 6366
rect 72920 6400 72924 6417
rect 72924 6400 72941 6417
rect 72941 6400 72946 6417
rect 72920 6396 72946 6400
rect 78302 6430 78328 6456
rect 73656 6396 73682 6422
rect 74668 6396 74694 6422
rect 73702 6362 73728 6388
rect 73886 6383 73912 6388
rect 66940 6328 66966 6354
rect 72874 6328 72900 6354
rect 73886 6366 73890 6383
rect 73890 6366 73907 6383
rect 73907 6366 73912 6383
rect 73886 6362 73912 6366
rect 74484 6362 74510 6388
rect 74622 6383 74648 6388
rect 74622 6366 74626 6383
rect 74626 6366 74643 6383
rect 74643 6366 74648 6383
rect 74622 6362 74648 6366
rect 75220 6396 75246 6422
rect 77934 6396 77960 6422
rect 78900 6396 78926 6422
rect 80188 6430 80214 6456
rect 80832 6396 80858 6422
rect 75772 6383 75798 6388
rect 75772 6366 75776 6383
rect 75776 6366 75793 6383
rect 75793 6366 75798 6383
rect 75772 6362 75798 6366
rect 75174 6328 75200 6354
rect 75818 6328 75844 6354
rect 74254 6294 74280 6320
rect 74990 6315 75016 6320
rect 74990 6298 74994 6315
rect 74994 6298 75011 6315
rect 75011 6298 75016 6315
rect 74990 6294 75016 6298
rect 75634 6294 75660 6320
rect 75680 6294 75706 6320
rect 76370 6362 76396 6388
rect 76416 6328 76442 6354
rect 76554 6328 76580 6354
rect 77520 6383 77546 6388
rect 77520 6366 77524 6383
rect 77524 6366 77541 6383
rect 77541 6366 77546 6383
rect 79728 6383 79754 6388
rect 77520 6362 77546 6366
rect 79406 6349 79432 6354
rect 79406 6332 79410 6349
rect 79410 6332 79427 6349
rect 79427 6332 79432 6349
rect 79406 6328 79432 6332
rect 79728 6366 79732 6383
rect 79732 6366 79749 6383
rect 79749 6366 79754 6383
rect 79728 6362 79754 6366
rect 79774 6362 79800 6388
rect 80786 6362 80812 6388
rect 77060 6294 77086 6320
rect 78946 6294 78972 6320
rect 80142 6294 80168 6320
rect 81752 6464 81778 6490
rect 81706 6430 81732 6456
rect 82626 6464 82652 6490
rect 81062 6383 81088 6388
rect 81062 6366 81066 6383
rect 81066 6366 81083 6383
rect 81083 6366 81088 6383
rect 81062 6362 81088 6366
rect 81430 6362 81456 6388
rect 83592 6464 83618 6490
rect 87502 6485 87528 6490
rect 87502 6468 87506 6485
rect 87506 6468 87523 6485
rect 87523 6468 87528 6485
rect 87502 6464 87528 6468
rect 87870 6464 87896 6490
rect 88192 6464 88218 6490
rect 82718 6396 82744 6422
rect 83086 6396 83112 6422
rect 83270 6417 83296 6422
rect 83270 6400 83274 6417
rect 83274 6400 83291 6417
rect 83291 6400 83296 6417
rect 83270 6396 83296 6400
rect 86904 6430 86930 6456
rect 87962 6430 87988 6456
rect 88468 6430 88494 6456
rect 88974 6430 89000 6456
rect 88192 6417 88218 6422
rect 82304 6383 82330 6388
rect 82304 6366 82308 6383
rect 82308 6366 82325 6383
rect 82325 6366 82330 6383
rect 82304 6362 82330 6366
rect 81844 6294 81870 6320
rect 82120 6328 82146 6354
rect 88192 6400 88196 6417
rect 88196 6400 88213 6417
rect 88213 6400 88218 6417
rect 88192 6396 88218 6400
rect 90078 6464 90104 6490
rect 90124 6464 90150 6490
rect 90170 6396 90196 6422
rect 90768 6417 90794 6422
rect 90768 6400 90772 6417
rect 90772 6400 90789 6417
rect 90789 6400 90794 6417
rect 94172 6464 94198 6490
rect 95690 6464 95716 6490
rect 96242 6464 96268 6490
rect 94264 6430 94290 6456
rect 95460 6451 95486 6456
rect 90768 6396 90794 6400
rect 94172 6396 94198 6422
rect 94402 6396 94428 6422
rect 94678 6417 94704 6422
rect 94678 6400 94682 6417
rect 94682 6400 94699 6417
rect 94699 6400 94704 6417
rect 94678 6396 94704 6400
rect 88376 6362 88402 6388
rect 90078 6362 90104 6388
rect 94770 6362 94796 6388
rect 95460 6434 95464 6451
rect 95464 6434 95481 6451
rect 95481 6434 95486 6451
rect 95460 6430 95486 6434
rect 95874 6430 95900 6456
rect 96978 6464 97004 6490
rect 97438 6464 97464 6490
rect 97990 6485 98016 6490
rect 97990 6468 97994 6485
rect 97994 6468 98011 6485
rect 98011 6468 98016 6485
rect 97990 6464 98016 6468
rect 98864 6464 98890 6490
rect 96288 6396 96314 6422
rect 97530 6417 97556 6422
rect 97530 6400 97534 6417
rect 97534 6400 97551 6417
rect 97551 6400 97556 6417
rect 97530 6396 97556 6400
rect 98680 6417 98706 6422
rect 98680 6400 98684 6417
rect 98684 6400 98701 6417
rect 98701 6400 98706 6417
rect 98680 6396 98706 6400
rect 98726 6417 98752 6422
rect 98726 6400 98730 6417
rect 98730 6400 98747 6417
rect 98747 6400 98752 6417
rect 99186 6417 99212 6422
rect 98726 6396 98752 6400
rect 96334 6362 96360 6388
rect 96518 6383 96544 6388
rect 96518 6366 96522 6383
rect 96522 6366 96539 6383
rect 96539 6366 96544 6383
rect 96518 6362 96544 6366
rect 83086 6294 83112 6320
rect 83316 6315 83342 6320
rect 83316 6298 83320 6315
rect 83320 6298 83337 6315
rect 83337 6298 83342 6315
rect 83316 6294 83342 6298
rect 90124 6328 90150 6354
rect 90262 6328 90288 6354
rect 91044 6328 91070 6354
rect 94310 6328 94336 6354
rect 94586 6328 94612 6354
rect 95874 6328 95900 6354
rect 95966 6328 95992 6354
rect 96242 6328 96268 6354
rect 97392 6362 97418 6388
rect 97898 6362 97924 6388
rect 98818 6383 98844 6388
rect 98818 6366 98822 6383
rect 98822 6366 98839 6383
rect 98839 6366 98844 6383
rect 98818 6362 98844 6366
rect 99186 6400 99190 6417
rect 99190 6400 99207 6417
rect 99207 6400 99212 6417
rect 99186 6396 99212 6400
rect 100336 6396 100362 6422
rect 100658 6417 100684 6422
rect 100658 6400 100662 6417
rect 100662 6400 100679 6417
rect 100679 6400 100684 6417
rect 100658 6396 100684 6400
rect 99278 6362 99304 6388
rect 100198 6362 100224 6388
rect 101486 6430 101512 6456
rect 101670 6430 101696 6456
rect 102820 6430 102846 6456
rect 103280 6485 103306 6490
rect 103280 6468 103284 6485
rect 103284 6468 103301 6485
rect 103301 6468 103306 6485
rect 103280 6464 103306 6468
rect 103694 6464 103720 6490
rect 103924 6464 103950 6490
rect 101440 6383 101466 6388
rect 88698 6294 88724 6320
rect 88928 6294 88954 6320
rect 89940 6294 89966 6320
rect 90308 6294 90334 6320
rect 90722 6294 90748 6320
rect 93896 6294 93922 6320
rect 94494 6294 94520 6320
rect 95276 6315 95302 6320
rect 95276 6298 95280 6315
rect 95280 6298 95297 6315
rect 95297 6298 95302 6315
rect 95276 6294 95302 6298
rect 96012 6294 96038 6320
rect 96058 6294 96084 6320
rect 96518 6294 96544 6320
rect 101072 6328 101098 6354
rect 101440 6366 101444 6383
rect 101444 6366 101461 6383
rect 101461 6366 101466 6383
rect 101440 6362 101466 6366
rect 101486 6362 101512 6388
rect 102084 6362 102110 6388
rect 102544 6383 102570 6388
rect 102544 6366 102548 6383
rect 102548 6366 102565 6383
rect 102565 6366 102570 6383
rect 102544 6362 102570 6366
rect 102590 6362 102616 6388
rect 105304 6430 105330 6456
rect 109904 6464 109930 6490
rect 103832 6396 103858 6422
rect 108294 6396 108320 6422
rect 114136 6430 114162 6456
rect 115194 6430 115220 6456
rect 109904 6396 109930 6422
rect 111836 6396 111862 6422
rect 113400 6396 113426 6422
rect 113952 6417 113978 6422
rect 113952 6400 113956 6417
rect 113956 6400 113973 6417
rect 113973 6400 113978 6417
rect 113952 6396 113978 6400
rect 115148 6417 115174 6422
rect 115148 6400 115152 6417
rect 115152 6400 115169 6417
rect 115169 6400 115174 6417
rect 115148 6396 115174 6400
rect 119104 6464 119130 6490
rect 115516 6451 115542 6456
rect 115516 6434 115520 6451
rect 115520 6434 115537 6451
rect 115537 6434 115542 6451
rect 115516 6430 115542 6434
rect 116160 6430 116186 6456
rect 119150 6430 119176 6456
rect 116528 6417 116554 6422
rect 103648 6349 103674 6354
rect 97208 6294 97234 6320
rect 97990 6294 98016 6320
rect 99094 6315 99120 6320
rect 99094 6298 99098 6315
rect 99098 6298 99115 6315
rect 99115 6298 99120 6315
rect 99094 6294 99120 6298
rect 100566 6315 100592 6320
rect 100566 6298 100570 6315
rect 100570 6298 100587 6315
rect 100587 6298 100592 6315
rect 100566 6294 100592 6298
rect 100980 6294 101006 6320
rect 102130 6294 102156 6320
rect 102268 6294 102294 6320
rect 102590 6294 102616 6320
rect 102636 6294 102662 6320
rect 103648 6332 103652 6349
rect 103652 6332 103669 6349
rect 103669 6332 103674 6349
rect 103648 6328 103674 6332
rect 105304 6294 105330 6320
rect 109904 6328 109930 6354
rect 113446 6294 113472 6320
rect 114136 6362 114162 6388
rect 115102 6362 115128 6388
rect 116528 6400 116532 6417
rect 116532 6400 116549 6417
rect 116549 6400 116554 6417
rect 116528 6396 116554 6400
rect 118506 6417 118532 6422
rect 118506 6400 118510 6417
rect 118510 6400 118527 6417
rect 118527 6400 118532 6417
rect 118506 6396 118532 6400
rect 119196 6396 119222 6422
rect 119518 6430 119544 6456
rect 120024 6430 120050 6456
rect 125544 6464 125570 6490
rect 127338 6464 127364 6490
rect 128120 6464 128146 6490
rect 132306 6485 132332 6490
rect 120484 6451 120510 6456
rect 120484 6434 120488 6451
rect 120488 6434 120505 6451
rect 120505 6434 120510 6451
rect 120484 6430 120510 6434
rect 121036 6396 121062 6422
rect 121128 6396 121154 6422
rect 122324 6430 122350 6456
rect 122462 6430 122488 6456
rect 122692 6430 122718 6456
rect 125820 6430 125846 6456
rect 126234 6451 126260 6456
rect 126234 6434 126238 6451
rect 126238 6434 126255 6451
rect 126255 6434 126260 6451
rect 126234 6430 126260 6434
rect 122278 6417 122304 6422
rect 122278 6400 122282 6417
rect 122282 6400 122299 6417
rect 122299 6400 122304 6417
rect 122278 6396 122304 6400
rect 122416 6396 122442 6422
rect 125590 6396 125616 6422
rect 125774 6417 125800 6422
rect 125774 6400 125778 6417
rect 125778 6400 125795 6417
rect 125795 6400 125800 6417
rect 125774 6396 125800 6400
rect 128304 6396 128330 6422
rect 118920 6328 118946 6354
rect 118966 6328 118992 6354
rect 114780 6294 114806 6320
rect 115056 6315 115082 6320
rect 115056 6298 115060 6315
rect 115060 6298 115077 6315
rect 115077 6298 115082 6315
rect 115056 6294 115082 6298
rect 115102 6294 115128 6320
rect 116160 6294 116186 6320
rect 116252 6315 116278 6320
rect 116252 6298 116256 6315
rect 116256 6298 116273 6315
rect 116273 6298 116278 6315
rect 116252 6294 116278 6298
rect 116574 6294 116600 6320
rect 119242 6294 119268 6320
rect 119426 6294 119452 6320
rect 119564 6294 119590 6320
rect 120162 6294 120188 6320
rect 121082 6328 121108 6354
rect 121220 6315 121246 6320
rect 121220 6298 121224 6315
rect 121224 6298 121241 6315
rect 121241 6298 121246 6315
rect 121220 6294 121246 6298
rect 121450 6294 121476 6320
rect 122324 6328 122350 6354
rect 124164 6328 124190 6354
rect 125084 6349 125110 6354
rect 125084 6332 125088 6349
rect 125088 6332 125105 6349
rect 125105 6332 125110 6349
rect 125084 6328 125110 6332
rect 126050 6362 126076 6388
rect 126832 6383 126858 6388
rect 126832 6366 126836 6383
rect 126836 6366 126853 6383
rect 126853 6366 126858 6383
rect 126832 6362 126858 6366
rect 126970 6383 126996 6388
rect 126970 6366 126974 6383
rect 126974 6366 126991 6383
rect 126991 6366 126996 6383
rect 126970 6362 126996 6366
rect 127568 6362 127594 6388
rect 128166 6383 128192 6388
rect 128166 6366 128170 6383
rect 128170 6366 128187 6383
rect 128187 6366 128192 6383
rect 128166 6362 128192 6366
rect 128212 6383 128238 6388
rect 128212 6366 128216 6383
rect 128216 6366 128233 6383
rect 128233 6366 128238 6383
rect 128212 6362 128238 6366
rect 125912 6328 125938 6354
rect 127522 6328 127548 6354
rect 125958 6294 125984 6320
rect 126004 6315 126030 6320
rect 126004 6298 126008 6315
rect 126008 6298 126025 6315
rect 126025 6298 126030 6315
rect 128626 6430 128652 6456
rect 130880 6451 130906 6456
rect 130880 6434 130884 6451
rect 130884 6434 130901 6451
rect 130901 6434 130906 6451
rect 130880 6430 130906 6434
rect 131662 6430 131688 6456
rect 132306 6468 132310 6485
rect 132310 6468 132327 6485
rect 132327 6468 132332 6485
rect 132306 6464 132332 6468
rect 134192 6464 134218 6490
rect 151304 6485 151330 6490
rect 132766 6451 132792 6456
rect 130926 6396 130952 6422
rect 132168 6396 132194 6422
rect 132214 6396 132240 6422
rect 132766 6434 132770 6451
rect 132770 6434 132787 6451
rect 132787 6434 132792 6451
rect 132766 6430 132792 6434
rect 133272 6430 133298 6456
rect 128580 6362 128606 6388
rect 131156 6362 131182 6388
rect 135526 6430 135552 6456
rect 135894 6451 135920 6456
rect 135894 6434 135898 6451
rect 135898 6434 135915 6451
rect 135915 6434 135920 6451
rect 135894 6430 135920 6434
rect 136400 6430 136426 6456
rect 136584 6430 136610 6456
rect 134146 6396 134172 6422
rect 134514 6396 134540 6422
rect 128534 6328 128560 6354
rect 131340 6349 131366 6354
rect 126004 6294 126030 6298
rect 131110 6294 131136 6320
rect 131340 6332 131344 6349
rect 131344 6332 131361 6349
rect 131361 6332 131366 6349
rect 131340 6328 131366 6332
rect 133502 6362 133528 6388
rect 133778 6362 133804 6388
rect 134008 6383 134034 6388
rect 134008 6366 134012 6383
rect 134012 6366 134029 6383
rect 134029 6366 134034 6383
rect 134008 6362 134034 6366
rect 134192 6362 134218 6388
rect 135434 6396 135460 6422
rect 136308 6396 136334 6422
rect 147946 6430 147972 6456
rect 151304 6468 151308 6485
rect 151308 6468 151325 6485
rect 151325 6468 151330 6485
rect 151304 6464 151330 6468
rect 152684 6464 152710 6490
rect 152500 6451 152526 6456
rect 134698 6383 134724 6388
rect 134698 6366 134702 6383
rect 134702 6366 134719 6383
rect 134719 6366 134724 6383
rect 134698 6362 134724 6366
rect 131754 6328 131780 6354
rect 131984 6315 132010 6320
rect 131984 6298 131988 6315
rect 131988 6298 132005 6315
rect 132005 6298 132010 6315
rect 131984 6294 132010 6298
rect 133502 6315 133528 6320
rect 133502 6298 133506 6315
rect 133506 6298 133523 6315
rect 133523 6298 133528 6315
rect 133502 6294 133528 6298
rect 133548 6294 133574 6320
rect 133778 6294 133804 6320
rect 134560 6294 134586 6320
rect 136124 6362 136150 6388
rect 136446 6362 136472 6388
rect 136400 6328 136426 6354
rect 136584 6362 136610 6388
rect 145140 6396 145166 6422
rect 151396 6417 151422 6422
rect 151396 6400 151400 6417
rect 151400 6400 151417 6417
rect 151417 6400 151422 6417
rect 151396 6396 151422 6400
rect 152500 6434 152504 6451
rect 152504 6434 152521 6451
rect 152521 6434 152526 6451
rect 152730 6451 152756 6456
rect 152500 6430 152526 6434
rect 152730 6434 152734 6451
rect 152734 6434 152751 6451
rect 152751 6434 152756 6451
rect 152730 6430 152756 6434
rect 135434 6315 135460 6320
rect 135434 6298 135438 6315
rect 135438 6298 135455 6315
rect 135455 6298 135460 6315
rect 135434 6294 135460 6298
rect 135572 6294 135598 6320
rect 136262 6315 136288 6320
rect 136262 6298 136266 6315
rect 136266 6298 136283 6315
rect 136283 6298 136288 6315
rect 136262 6294 136288 6298
rect 136308 6294 136334 6320
rect 140540 6294 140566 6320
rect 19524 6243 19550 6269
rect 19556 6243 19582 6269
rect 19588 6243 19614 6269
rect 19620 6243 19646 6269
rect 19652 6243 19678 6269
rect 57623 6243 57649 6269
rect 57655 6243 57681 6269
rect 57687 6243 57713 6269
rect 57719 6243 57745 6269
rect 57751 6243 57777 6269
rect 95722 6243 95748 6269
rect 95754 6243 95780 6269
rect 95786 6243 95812 6269
rect 95818 6243 95844 6269
rect 95850 6243 95876 6269
rect 133821 6243 133847 6269
rect 133853 6243 133879 6269
rect 133885 6243 133911 6269
rect 133917 6243 133943 6269
rect 133949 6243 133975 6269
rect 13488 6192 13514 6218
rect 14040 6192 14066 6218
rect 7140 6158 7166 6184
rect 14408 6192 14434 6218
rect 16294 6192 16320 6218
rect 17260 6192 17286 6218
rect 17996 6192 18022 6218
rect 2402 6022 2428 6048
rect 13442 6124 13468 6150
rect 14040 6124 14066 6150
rect 14362 6145 14388 6150
rect 14362 6128 14366 6145
rect 14366 6128 14383 6145
rect 14383 6128 14388 6145
rect 14362 6124 14388 6128
rect 17444 6158 17470 6184
rect 18916 6192 18942 6218
rect 19468 6192 19494 6218
rect 19698 6192 19724 6218
rect 20480 6192 20506 6218
rect 21584 6213 21610 6218
rect 21584 6196 21588 6213
rect 21588 6196 21605 6213
rect 21605 6196 21610 6213
rect 21584 6192 21610 6196
rect 21906 6213 21932 6218
rect 21906 6196 21910 6213
rect 21910 6196 21927 6213
rect 21927 6196 21932 6213
rect 21906 6192 21932 6196
rect 27012 6192 27038 6218
rect 27748 6192 27774 6218
rect 28346 6192 28372 6218
rect 28990 6213 29016 6218
rect 28990 6196 28994 6213
rect 28994 6196 29011 6213
rect 29011 6196 29016 6213
rect 28990 6192 29016 6196
rect 37546 6192 37572 6218
rect 39662 6213 39688 6218
rect 14500 6124 14526 6150
rect 14776 6145 14802 6150
rect 14776 6128 14780 6145
rect 14780 6128 14797 6145
rect 14797 6128 14802 6145
rect 14776 6124 14802 6128
rect 8520 6090 8546 6116
rect 13718 6111 13744 6116
rect 13718 6094 13722 6111
rect 13722 6094 13739 6111
rect 13739 6094 13744 6111
rect 13718 6090 13744 6094
rect 14684 6090 14710 6116
rect 17076 6111 17102 6116
rect 17076 6094 17080 6111
rect 17080 6094 17097 6111
rect 17097 6094 17102 6111
rect 17076 6090 17102 6094
rect 17352 6111 17378 6116
rect 17352 6094 17356 6111
rect 17356 6094 17373 6111
rect 17373 6094 17378 6111
rect 17674 6111 17700 6116
rect 17352 6090 17378 6094
rect 17674 6094 17678 6111
rect 17678 6094 17695 6111
rect 17695 6094 17700 6111
rect 17674 6090 17700 6094
rect 13534 6043 13560 6048
rect 13534 6026 13538 6043
rect 13538 6026 13555 6043
rect 13555 6026 13560 6043
rect 13534 6022 13560 6026
rect 13580 6022 13606 6048
rect 13994 6022 14020 6048
rect 14730 6056 14756 6082
rect 14914 6077 14940 6082
rect 14914 6060 14918 6077
rect 14918 6060 14935 6077
rect 14935 6060 14940 6077
rect 14914 6056 14940 6060
rect 15604 6056 15630 6082
rect 16018 6077 16044 6082
rect 16018 6060 16022 6077
rect 16022 6060 16039 6077
rect 16039 6060 16044 6077
rect 16018 6056 16044 6060
rect 21860 6158 21886 6184
rect 20480 6124 20506 6150
rect 19008 6090 19034 6116
rect 20158 6090 20184 6116
rect 20296 6111 20322 6116
rect 20296 6094 20300 6111
rect 20300 6094 20317 6111
rect 20317 6094 20322 6111
rect 20296 6090 20322 6094
rect 38006 6158 38032 6184
rect 26920 6124 26946 6150
rect 21860 6111 21886 6116
rect 21860 6094 21864 6111
rect 21864 6094 21881 6111
rect 21881 6094 21886 6111
rect 21860 6090 21886 6094
rect 20802 6056 20828 6082
rect 20894 6056 20920 6082
rect 14454 6022 14480 6048
rect 15558 6022 15584 6048
rect 16156 6022 16182 6048
rect 16478 6022 16504 6048
rect 18226 6043 18252 6048
rect 18226 6026 18230 6043
rect 18230 6026 18247 6043
rect 18247 6026 18252 6043
rect 18226 6022 18252 6026
rect 20250 6022 20276 6048
rect 20342 6043 20368 6048
rect 20342 6026 20346 6043
rect 20346 6026 20363 6043
rect 20363 6026 20368 6043
rect 20342 6022 20368 6026
rect 28208 6124 28234 6150
rect 37408 6124 37434 6150
rect 38604 6158 38630 6184
rect 39202 6158 39228 6184
rect 27656 6090 27682 6116
rect 28254 6090 28280 6116
rect 38466 6145 38492 6150
rect 38466 6128 38470 6145
rect 38470 6128 38487 6145
rect 38487 6128 38492 6145
rect 39064 6145 39090 6150
rect 38466 6124 38492 6128
rect 39064 6128 39068 6145
rect 39068 6128 39085 6145
rect 39085 6128 39090 6145
rect 39064 6124 39090 6128
rect 26322 6077 26348 6082
rect 26322 6060 26326 6077
rect 26326 6060 26343 6077
rect 26343 6060 26348 6077
rect 26322 6056 26348 6060
rect 26552 6056 26578 6082
rect 38972 6111 38998 6116
rect 38972 6094 38976 6111
rect 38976 6094 38993 6111
rect 38993 6094 38998 6111
rect 38972 6090 38998 6094
rect 39662 6196 39666 6213
rect 39666 6196 39683 6213
rect 39683 6196 39688 6213
rect 39662 6192 39688 6196
rect 40260 6192 40286 6218
rect 42744 6192 42770 6218
rect 43204 6213 43230 6218
rect 43204 6196 43208 6213
rect 43208 6196 43225 6213
rect 43225 6196 43230 6213
rect 43204 6192 43230 6196
rect 43940 6192 43966 6218
rect 45090 6213 45116 6218
rect 45090 6196 45094 6213
rect 45094 6196 45111 6213
rect 45111 6196 45116 6213
rect 45090 6192 45116 6196
rect 49736 6192 49762 6218
rect 49966 6192 49992 6218
rect 52496 6192 52522 6218
rect 52588 6213 52614 6218
rect 52588 6196 52592 6213
rect 52592 6196 52609 6213
rect 52609 6196 52614 6213
rect 52588 6192 52614 6196
rect 56268 6192 56294 6218
rect 57510 6192 57536 6218
rect 58476 6192 58502 6218
rect 63904 6192 63930 6218
rect 64548 6192 64574 6218
rect 65468 6192 65494 6218
rect 66204 6192 66230 6218
rect 73886 6192 73912 6218
rect 76232 6192 76258 6218
rect 39294 6090 39320 6116
rect 43066 6158 43092 6184
rect 43710 6158 43736 6184
rect 40720 6124 40746 6150
rect 42330 6145 42356 6150
rect 42330 6128 42334 6145
rect 42334 6128 42351 6145
rect 42351 6128 42356 6145
rect 42330 6124 42356 6128
rect 41916 6090 41942 6116
rect 42882 6124 42908 6150
rect 43158 6124 43184 6150
rect 44078 6145 44104 6150
rect 44078 6128 44082 6145
rect 44082 6128 44099 6145
rect 44099 6128 44104 6145
rect 44078 6124 44104 6128
rect 42744 6111 42770 6116
rect 42744 6094 42748 6111
rect 42748 6094 42765 6111
rect 42765 6094 42770 6111
rect 42744 6090 42770 6094
rect 43020 6090 43046 6116
rect 44124 6090 44150 6116
rect 44584 6124 44610 6150
rect 44492 6090 44518 6116
rect 46010 6090 46036 6116
rect 49552 6124 49578 6150
rect 51024 6124 51050 6150
rect 51622 6124 51648 6150
rect 51668 6124 51694 6150
rect 57878 6158 57904 6184
rect 48770 6090 48796 6116
rect 51852 6090 51878 6116
rect 50380 6077 50406 6082
rect 27932 6022 27958 6048
rect 28024 6043 28050 6048
rect 28024 6026 28028 6043
rect 28028 6026 28045 6043
rect 28045 6026 28050 6043
rect 28024 6022 28050 6026
rect 28668 6022 28694 6048
rect 38144 6043 38170 6048
rect 38144 6026 38148 6043
rect 38148 6026 38165 6043
rect 38165 6026 38170 6043
rect 38144 6022 38170 6026
rect 40122 6022 40148 6048
rect 42008 6043 42034 6048
rect 42008 6026 42012 6043
rect 42012 6026 42029 6043
rect 42029 6026 42034 6043
rect 42008 6022 42034 6026
rect 42330 6022 42356 6048
rect 43158 6022 43184 6048
rect 43756 6022 43782 6048
rect 43894 6022 43920 6048
rect 43986 6022 44012 6048
rect 44354 6022 44380 6048
rect 50380 6060 50384 6077
rect 50384 6060 50401 6077
rect 50401 6060 50406 6077
rect 50380 6056 50406 6060
rect 50518 6056 50544 6082
rect 50978 6077 51004 6082
rect 50978 6060 50982 6077
rect 50982 6060 50999 6077
rect 50999 6060 51004 6077
rect 50978 6056 51004 6060
rect 51070 6077 51096 6082
rect 51070 6060 51074 6077
rect 51074 6060 51091 6077
rect 51091 6060 51096 6077
rect 55946 6090 55972 6116
rect 57142 6090 57168 6116
rect 59442 6124 59468 6150
rect 70988 6158 71014 6184
rect 73794 6158 73820 6184
rect 75818 6158 75844 6184
rect 51070 6056 51096 6060
rect 56912 6056 56938 6082
rect 50196 6043 50222 6048
rect 50196 6026 50200 6043
rect 50200 6026 50217 6043
rect 50217 6026 50222 6043
rect 50196 6022 50222 6026
rect 51162 6022 51188 6048
rect 51300 6043 51326 6048
rect 51300 6026 51304 6043
rect 51304 6026 51321 6043
rect 51321 6026 51326 6043
rect 51300 6022 51326 6026
rect 51530 6043 51556 6048
rect 51530 6026 51534 6043
rect 51534 6026 51551 6043
rect 51551 6026 51556 6043
rect 51530 6022 51556 6026
rect 56958 6022 56984 6048
rect 57832 6022 57858 6048
rect 58200 6022 58226 6048
rect 59028 6090 59054 6116
rect 59166 6111 59192 6116
rect 59166 6094 59170 6111
rect 59170 6094 59187 6111
rect 59187 6094 59192 6111
rect 59166 6090 59192 6094
rect 63076 6090 63102 6116
rect 64318 6111 64344 6116
rect 64318 6094 64322 6111
rect 64322 6094 64339 6111
rect 64339 6094 64344 6111
rect 64318 6090 64344 6094
rect 65514 6124 65540 6150
rect 66618 6124 66644 6150
rect 74530 6124 74556 6150
rect 59120 6056 59146 6082
rect 65238 6090 65264 6116
rect 66204 6090 66230 6116
rect 66296 6111 66322 6116
rect 66296 6094 66300 6111
rect 66300 6094 66317 6111
rect 66317 6094 66322 6111
rect 66296 6090 66322 6094
rect 68872 6111 68898 6116
rect 68872 6094 68876 6111
rect 68876 6094 68893 6111
rect 68893 6094 68898 6111
rect 68872 6090 68898 6094
rect 74024 6090 74050 6116
rect 74668 6090 74694 6116
rect 74714 6111 74740 6116
rect 74714 6094 74718 6111
rect 74718 6094 74735 6111
rect 74735 6094 74740 6111
rect 74714 6090 74740 6094
rect 75680 6090 75706 6116
rect 76370 6158 76396 6184
rect 66250 6056 66276 6082
rect 69010 6077 69036 6082
rect 69010 6060 69014 6077
rect 69014 6060 69031 6077
rect 69031 6060 69036 6077
rect 69010 6056 69036 6060
rect 76876 6192 76902 6218
rect 78624 6192 78650 6218
rect 80464 6192 80490 6218
rect 80786 6192 80812 6218
rect 77520 6158 77546 6184
rect 79452 6158 79478 6184
rect 83224 6192 83250 6218
rect 88238 6192 88264 6218
rect 89756 6192 89782 6218
rect 94586 6192 94612 6218
rect 94816 6192 94842 6218
rect 95414 6192 95440 6218
rect 97024 6192 97050 6218
rect 82718 6158 82744 6184
rect 83040 6179 83066 6184
rect 83040 6162 83044 6179
rect 83044 6162 83061 6179
rect 83061 6162 83066 6179
rect 83040 6158 83066 6162
rect 77060 6124 77086 6150
rect 80188 6124 80214 6150
rect 80740 6145 80766 6150
rect 80740 6128 80744 6145
rect 80744 6128 80761 6145
rect 80761 6128 80766 6145
rect 81246 6145 81272 6150
rect 80740 6124 80766 6128
rect 81246 6128 81250 6145
rect 81250 6128 81267 6145
rect 81267 6128 81272 6145
rect 81246 6124 81272 6128
rect 81338 6145 81364 6150
rect 81338 6128 81342 6145
rect 81342 6128 81359 6145
rect 81359 6128 81364 6145
rect 81338 6124 81364 6128
rect 81798 6145 81824 6150
rect 81798 6128 81802 6145
rect 81802 6128 81819 6145
rect 81819 6128 81824 6145
rect 81798 6124 81824 6128
rect 88882 6158 88908 6184
rect 90446 6179 90472 6184
rect 90446 6162 90450 6179
rect 90450 6162 90467 6179
rect 90467 6162 90472 6179
rect 90446 6158 90472 6162
rect 96288 6179 96314 6184
rect 88560 6145 88586 6150
rect 88560 6128 88564 6145
rect 88564 6128 88581 6145
rect 88581 6128 88586 6145
rect 88560 6124 88586 6128
rect 79406 6090 79432 6116
rect 80878 6090 80904 6116
rect 93988 6124 94014 6150
rect 88928 6090 88954 6116
rect 89572 6111 89598 6116
rect 89572 6094 89576 6111
rect 89576 6094 89593 6111
rect 89593 6094 89598 6111
rect 89572 6090 89598 6094
rect 90354 6090 90380 6116
rect 94770 6111 94796 6116
rect 65790 6022 65816 6048
rect 77934 6056 77960 6082
rect 78210 6056 78236 6082
rect 81292 6056 81318 6082
rect 81338 6056 81364 6082
rect 82166 6056 82192 6082
rect 82948 6077 82974 6082
rect 82948 6060 82952 6077
rect 82952 6060 82969 6077
rect 82969 6060 82974 6077
rect 82948 6056 82974 6060
rect 83270 6056 83296 6082
rect 89710 6077 89736 6082
rect 74760 6022 74786 6048
rect 75818 6043 75844 6048
rect 75818 6026 75822 6043
rect 75822 6026 75839 6043
rect 75839 6026 75844 6043
rect 75818 6022 75844 6026
rect 75864 6022 75890 6048
rect 76094 6022 76120 6048
rect 76278 6022 76304 6048
rect 80556 6022 80582 6048
rect 81108 6022 81134 6048
rect 81430 6022 81456 6048
rect 88330 6022 88356 6048
rect 89020 6043 89046 6048
rect 89020 6026 89024 6043
rect 89024 6026 89041 6043
rect 89041 6026 89046 6043
rect 89020 6022 89046 6026
rect 89710 6060 89714 6077
rect 89714 6060 89731 6077
rect 89731 6060 89736 6077
rect 89710 6056 89736 6060
rect 90722 6056 90748 6082
rect 94770 6094 94774 6111
rect 94774 6094 94791 6111
rect 94791 6094 94796 6111
rect 94770 6090 94796 6094
rect 96288 6162 96292 6179
rect 96292 6162 96309 6179
rect 96309 6162 96314 6179
rect 96288 6158 96314 6162
rect 95920 6124 95946 6150
rect 96334 6124 96360 6150
rect 97208 6111 97234 6116
rect 95414 6056 95440 6082
rect 95552 6077 95578 6082
rect 95552 6060 95556 6077
rect 95556 6060 95573 6077
rect 95573 6060 95578 6077
rect 95552 6056 95578 6060
rect 95598 6056 95624 6082
rect 90078 6022 90104 6048
rect 96702 6077 96728 6082
rect 96702 6060 96706 6077
rect 96706 6060 96723 6077
rect 96723 6060 96728 6077
rect 96702 6056 96728 6060
rect 96518 6043 96544 6048
rect 96518 6026 96522 6043
rect 96522 6026 96539 6043
rect 96539 6026 96544 6043
rect 96518 6022 96544 6026
rect 96840 6022 96866 6048
rect 97208 6094 97212 6111
rect 97212 6094 97229 6111
rect 97229 6094 97234 6111
rect 97208 6090 97234 6094
rect 97346 6077 97372 6082
rect 97346 6060 97350 6077
rect 97350 6060 97367 6077
rect 97367 6060 97372 6077
rect 97346 6056 97372 6060
rect 98726 6158 98752 6184
rect 101210 6192 101236 6218
rect 102820 6192 102846 6218
rect 103832 6192 103858 6218
rect 115056 6192 115082 6218
rect 115930 6192 115956 6218
rect 119518 6192 119544 6218
rect 120070 6192 120096 6218
rect 114412 6158 114438 6184
rect 115562 6158 115588 6184
rect 116252 6158 116278 6184
rect 97484 6022 97510 6048
rect 100244 6124 100270 6150
rect 98726 6111 98752 6116
rect 98726 6094 98730 6111
rect 98730 6094 98747 6111
rect 98747 6094 98752 6111
rect 98726 6090 98752 6094
rect 99186 6090 99212 6116
rect 100290 6090 100316 6116
rect 100520 6111 100546 6116
rect 100520 6094 100524 6111
rect 100524 6094 100541 6111
rect 100541 6094 100546 6111
rect 100520 6090 100546 6094
rect 101026 6124 101052 6150
rect 101762 6145 101788 6150
rect 101762 6128 101766 6145
rect 101766 6128 101783 6145
rect 101783 6128 101788 6145
rect 101762 6124 101788 6128
rect 102268 6090 102294 6116
rect 114964 6111 114990 6116
rect 114964 6094 114968 6111
rect 114968 6094 114985 6111
rect 114985 6094 114990 6111
rect 114964 6090 114990 6094
rect 115654 6090 115680 6116
rect 102498 6077 102524 6082
rect 102498 6060 102502 6077
rect 102502 6060 102519 6077
rect 102519 6060 102524 6077
rect 102498 6056 102524 6060
rect 98404 6043 98430 6048
rect 98404 6026 98408 6043
rect 98408 6026 98425 6043
rect 98425 6026 98430 6043
rect 98404 6022 98430 6026
rect 98496 6043 98522 6048
rect 98496 6026 98500 6043
rect 98500 6026 98517 6043
rect 98517 6026 98522 6043
rect 98496 6022 98522 6026
rect 98680 6043 98706 6048
rect 98680 6026 98684 6043
rect 98684 6026 98701 6043
rect 98701 6026 98706 6043
rect 98680 6022 98706 6026
rect 101532 6022 101558 6048
rect 101716 6022 101742 6048
rect 102130 6022 102156 6048
rect 115424 6056 115450 6082
rect 115562 6056 115588 6082
rect 115838 6124 115864 6150
rect 119426 6124 119452 6150
rect 119656 6145 119682 6150
rect 119656 6128 119660 6145
rect 119660 6128 119677 6145
rect 119677 6128 119682 6145
rect 119656 6124 119682 6128
rect 116068 6111 116094 6116
rect 116068 6094 116072 6111
rect 116072 6094 116089 6111
rect 116089 6094 116094 6111
rect 116068 6090 116094 6094
rect 116528 6090 116554 6116
rect 119012 6111 119038 6116
rect 119012 6094 119016 6111
rect 119016 6094 119033 6111
rect 119033 6094 119038 6111
rect 119012 6090 119038 6094
rect 119196 6090 119222 6116
rect 119564 6111 119590 6116
rect 119564 6094 119568 6111
rect 119568 6094 119585 6111
rect 119585 6094 119590 6111
rect 119564 6090 119590 6094
rect 119748 6090 119774 6116
rect 119978 6124 120004 6150
rect 121128 6158 121154 6184
rect 121220 6124 121246 6150
rect 121496 6158 121522 6184
rect 121450 6145 121476 6150
rect 121450 6128 121454 6145
rect 121454 6128 121471 6145
rect 121471 6128 121476 6145
rect 121450 6124 121476 6128
rect 121082 6090 121108 6116
rect 121818 6192 121844 6218
rect 122094 6213 122120 6218
rect 122094 6196 122098 6213
rect 122098 6196 122115 6213
rect 122115 6196 122120 6213
rect 122094 6192 122120 6196
rect 125682 6192 125708 6218
rect 125958 6192 125984 6218
rect 125728 6158 125754 6184
rect 126050 6179 126076 6184
rect 126050 6162 126054 6179
rect 126054 6162 126071 6179
rect 126071 6162 126076 6179
rect 126050 6158 126076 6162
rect 127154 6179 127180 6184
rect 127154 6162 127158 6179
rect 127158 6162 127175 6179
rect 127175 6162 127180 6179
rect 127154 6158 127180 6162
rect 127614 6158 127640 6184
rect 121588 6124 121614 6150
rect 124164 6124 124190 6150
rect 124624 6124 124650 6150
rect 125636 6111 125662 6116
rect 125636 6094 125640 6111
rect 125640 6094 125657 6111
rect 125657 6094 125662 6111
rect 125958 6111 125984 6116
rect 125636 6090 125662 6094
rect 125958 6094 125962 6111
rect 125962 6094 125979 6111
rect 125979 6094 125984 6111
rect 125958 6090 125984 6094
rect 127568 6111 127594 6116
rect 127568 6094 127572 6111
rect 127572 6094 127589 6111
rect 127589 6094 127594 6111
rect 127568 6090 127594 6094
rect 124532 6077 124558 6082
rect 114412 6022 114438 6048
rect 115608 6022 115634 6048
rect 124532 6060 124536 6077
rect 124536 6060 124553 6077
rect 124553 6060 124558 6077
rect 124532 6056 124558 6060
rect 124624 6077 124650 6082
rect 124624 6060 124628 6077
rect 124628 6060 124645 6077
rect 124645 6060 124650 6077
rect 124624 6056 124650 6060
rect 126556 6056 126582 6082
rect 127798 6124 127824 6150
rect 128258 6192 128284 6218
rect 131248 6213 131274 6218
rect 131248 6196 131252 6213
rect 131252 6196 131269 6213
rect 131269 6196 131274 6213
rect 131248 6192 131274 6196
rect 132766 6192 132792 6218
rect 128488 6158 128514 6184
rect 132490 6158 132516 6184
rect 134008 6192 134034 6218
rect 134192 6192 134218 6218
rect 135526 6213 135552 6218
rect 135526 6196 135530 6213
rect 135530 6196 135547 6213
rect 135547 6196 135552 6213
rect 135526 6192 135552 6196
rect 152730 6213 152756 6218
rect 152730 6196 152734 6213
rect 152734 6196 152751 6213
rect 152751 6196 152756 6213
rect 152730 6192 152756 6196
rect 130926 6124 130952 6150
rect 131202 6124 131228 6150
rect 128120 6111 128146 6116
rect 128120 6094 128124 6111
rect 128124 6094 128141 6111
rect 128141 6094 128146 6111
rect 128120 6090 128146 6094
rect 128166 6090 128192 6116
rect 131524 6090 131550 6116
rect 132076 6124 132102 6150
rect 132582 6124 132608 6150
rect 132168 6090 132194 6116
rect 132812 6124 132838 6150
rect 134560 6124 134586 6150
rect 134836 6124 134862 6150
rect 135572 6124 135598 6150
rect 136124 6145 136150 6150
rect 136124 6128 136128 6145
rect 136128 6128 136145 6145
rect 136145 6128 136150 6145
rect 136124 6124 136150 6128
rect 136400 6124 136426 6150
rect 115700 6043 115726 6048
rect 115700 6026 115704 6043
rect 115704 6026 115721 6043
rect 115721 6026 115726 6043
rect 115700 6022 115726 6026
rect 115884 6022 115910 6048
rect 116528 6022 116554 6048
rect 120438 6043 120464 6048
rect 120438 6026 120442 6043
rect 120442 6026 120459 6043
rect 120459 6026 120464 6043
rect 120438 6022 120464 6026
rect 120760 6022 120786 6048
rect 121266 6022 121292 6048
rect 122048 6022 122074 6048
rect 127200 6022 127226 6048
rect 127522 6022 127548 6048
rect 127614 6043 127640 6048
rect 127614 6026 127618 6043
rect 127618 6026 127635 6043
rect 127635 6026 127640 6043
rect 127614 6022 127640 6026
rect 128166 6022 128192 6048
rect 132582 6056 132608 6082
rect 134054 6090 134080 6116
rect 134330 6090 134356 6116
rect 133410 6077 133436 6082
rect 133410 6060 133414 6077
rect 133414 6060 133431 6077
rect 133431 6060 133436 6077
rect 133410 6056 133436 6060
rect 133640 6056 133666 6082
rect 134100 6056 134126 6082
rect 134744 6056 134770 6082
rect 133502 6022 133528 6048
rect 134238 6022 134264 6048
rect 134330 6022 134356 6048
rect 135664 6090 135690 6116
rect 136446 6090 136472 6116
rect 135204 6022 135230 6048
rect 142380 6022 142406 6048
rect 38574 5971 38600 5997
rect 38606 5971 38632 5997
rect 38638 5971 38664 5997
rect 38670 5971 38696 5997
rect 38702 5971 38728 5997
rect 76673 5971 76699 5997
rect 76705 5971 76731 5997
rect 76737 5971 76763 5997
rect 76769 5971 76795 5997
rect 76801 5971 76827 5997
rect 114772 5971 114798 5997
rect 114804 5971 114830 5997
rect 114836 5971 114862 5997
rect 114868 5971 114894 5997
rect 114900 5971 114926 5997
rect 14546 5920 14572 5946
rect 14730 5920 14756 5946
rect 15466 5920 15492 5946
rect 16110 5920 16136 5946
rect 16892 5941 16918 5946
rect 16892 5924 16896 5941
rect 16896 5924 16913 5941
rect 16913 5924 16918 5941
rect 16892 5920 16918 5924
rect 17214 5941 17240 5946
rect 17214 5924 17218 5941
rect 17218 5924 17235 5941
rect 17235 5924 17240 5941
rect 17214 5920 17240 5924
rect 19192 5941 19218 5946
rect 13856 5886 13882 5912
rect 14362 5886 14388 5912
rect 14500 5886 14526 5912
rect 14454 5839 14480 5844
rect 14454 5822 14458 5839
rect 14458 5822 14475 5839
rect 14475 5822 14480 5839
rect 14454 5818 14480 5822
rect 15006 5886 15032 5912
rect 16018 5886 16044 5912
rect 19192 5924 19196 5941
rect 19196 5924 19213 5941
rect 19213 5924 19218 5941
rect 19192 5920 19218 5924
rect 19790 5920 19816 5946
rect 14776 5852 14802 5878
rect 16202 5852 16228 5878
rect 14960 5839 14986 5844
rect 14960 5822 14964 5839
rect 14964 5822 14981 5839
rect 14981 5822 14986 5839
rect 14960 5818 14986 5822
rect 14224 5771 14250 5776
rect 14224 5754 14228 5771
rect 14228 5754 14245 5771
rect 14245 5754 14250 5771
rect 14224 5750 14250 5754
rect 16294 5818 16320 5844
rect 17352 5852 17378 5878
rect 19974 5920 20000 5946
rect 20710 5920 20736 5946
rect 21446 5920 21472 5946
rect 26322 5920 26348 5946
rect 26828 5941 26854 5946
rect 26828 5924 26832 5941
rect 26832 5924 26849 5941
rect 26849 5924 26854 5941
rect 26828 5920 26854 5924
rect 27196 5941 27222 5946
rect 27196 5924 27200 5941
rect 27200 5924 27217 5941
rect 27217 5924 27222 5941
rect 27196 5920 27222 5924
rect 27656 5941 27682 5946
rect 27656 5924 27660 5941
rect 27660 5924 27677 5941
rect 27677 5924 27682 5941
rect 27656 5920 27682 5924
rect 28300 5920 28326 5946
rect 29312 5920 29338 5946
rect 37730 5920 37756 5946
rect 37822 5920 37848 5946
rect 38236 5920 38262 5946
rect 38926 5941 38952 5946
rect 38926 5924 38930 5941
rect 38930 5924 38947 5941
rect 38947 5924 38952 5941
rect 38926 5920 38952 5924
rect 39248 5941 39274 5946
rect 39248 5924 39252 5941
rect 39252 5924 39269 5941
rect 39269 5924 39274 5941
rect 39248 5920 39274 5924
rect 42146 5920 42172 5946
rect 43020 5941 43046 5946
rect 17030 5818 17056 5844
rect 15558 5784 15584 5810
rect 20342 5886 20368 5912
rect 20618 5886 20644 5912
rect 26874 5886 26900 5912
rect 20158 5852 20184 5878
rect 21400 5852 21426 5878
rect 21492 5852 21518 5878
rect 26506 5873 26532 5878
rect 20480 5818 20506 5844
rect 20710 5818 20736 5844
rect 26506 5856 26510 5873
rect 26510 5856 26527 5873
rect 26527 5856 26532 5873
rect 26506 5852 26532 5856
rect 28714 5886 28740 5912
rect 42468 5886 42494 5912
rect 27334 5818 27360 5844
rect 27794 5839 27820 5844
rect 27794 5822 27798 5839
rect 27798 5822 27815 5839
rect 27815 5822 27820 5839
rect 27794 5818 27820 5822
rect 27932 5818 27958 5844
rect 38006 5852 38032 5878
rect 38144 5852 38170 5878
rect 39294 5852 39320 5878
rect 40720 5852 40746 5878
rect 43020 5924 43024 5941
rect 43024 5924 43041 5941
rect 43041 5924 43046 5941
rect 43020 5920 43046 5924
rect 43066 5920 43092 5946
rect 43940 5941 43966 5946
rect 43940 5924 43944 5941
rect 43944 5924 43961 5941
rect 43961 5924 43966 5941
rect 43940 5920 43966 5924
rect 44768 5920 44794 5946
rect 49828 5920 49854 5946
rect 50472 5941 50498 5946
rect 50472 5924 50476 5941
rect 50476 5924 50493 5941
rect 50493 5924 50498 5941
rect 50472 5920 50498 5924
rect 51530 5920 51556 5946
rect 51760 5920 51786 5946
rect 56912 5941 56938 5946
rect 42652 5886 42678 5912
rect 56912 5924 56916 5941
rect 56916 5924 56933 5941
rect 56933 5924 56938 5941
rect 56912 5920 56938 5924
rect 57142 5920 57168 5946
rect 57832 5920 57858 5946
rect 58384 5920 58410 5946
rect 58660 5920 58686 5946
rect 59396 5920 59422 5946
rect 64686 5941 64712 5946
rect 64686 5924 64690 5941
rect 64690 5924 64707 5941
rect 64707 5924 64712 5941
rect 64686 5920 64712 5924
rect 65146 5920 65172 5946
rect 65468 5941 65494 5946
rect 65468 5924 65472 5941
rect 65472 5924 65489 5941
rect 65489 5924 65494 5941
rect 65468 5920 65494 5924
rect 65560 5920 65586 5946
rect 68872 5920 68898 5946
rect 75542 5941 75568 5946
rect 37500 5818 37526 5844
rect 38466 5818 38492 5844
rect 42008 5818 42034 5844
rect 42882 5852 42908 5878
rect 43480 5873 43506 5878
rect 43480 5856 43484 5873
rect 43484 5856 43501 5873
rect 43501 5856 43506 5873
rect 43480 5852 43506 5856
rect 43158 5839 43184 5844
rect 43158 5822 43162 5839
rect 43162 5822 43179 5839
rect 43179 5822 43184 5839
rect 43158 5818 43184 5822
rect 44584 5852 44610 5878
rect 50196 5873 50222 5878
rect 50196 5856 50200 5873
rect 50200 5856 50217 5873
rect 50217 5856 50222 5873
rect 50196 5852 50222 5856
rect 51070 5852 51096 5878
rect 51806 5852 51832 5878
rect 28024 5784 28050 5810
rect 45228 5818 45254 5844
rect 50380 5818 50406 5844
rect 51024 5839 51050 5844
rect 51024 5822 51028 5839
rect 51028 5822 51045 5839
rect 51045 5822 51050 5839
rect 51024 5818 51050 5822
rect 51162 5818 51188 5844
rect 51760 5818 51786 5844
rect 57280 5886 57306 5912
rect 57004 5873 57030 5878
rect 57004 5856 57008 5873
rect 57008 5856 57025 5873
rect 57025 5856 57030 5873
rect 57004 5852 57030 5856
rect 69010 5886 69036 5912
rect 74990 5886 75016 5912
rect 75542 5924 75546 5941
rect 75546 5924 75563 5941
rect 75563 5924 75568 5941
rect 75542 5920 75568 5924
rect 76002 5941 76028 5946
rect 76002 5924 76006 5941
rect 76006 5924 76023 5941
rect 76023 5924 76028 5941
rect 76002 5920 76028 5924
rect 77106 5920 77132 5946
rect 57510 5852 57536 5878
rect 58200 5873 58226 5878
rect 58200 5856 58204 5873
rect 58204 5856 58221 5873
rect 58221 5856 58226 5873
rect 58200 5852 58226 5856
rect 57832 5818 57858 5844
rect 57878 5818 57904 5844
rect 59166 5852 59192 5878
rect 64180 5852 64206 5878
rect 65146 5852 65172 5878
rect 65790 5852 65816 5878
rect 64870 5818 64896 5844
rect 65514 5839 65540 5844
rect 65514 5822 65518 5839
rect 65518 5822 65535 5839
rect 65535 5822 65540 5839
rect 65514 5818 65540 5822
rect 66250 5852 66276 5878
rect 73840 5852 73866 5878
rect 75634 5873 75660 5878
rect 75634 5856 75638 5873
rect 75638 5856 75655 5873
rect 75655 5856 75660 5873
rect 75634 5852 75660 5856
rect 76094 5873 76120 5878
rect 76094 5856 76098 5873
rect 76098 5856 76115 5873
rect 76115 5856 76120 5873
rect 76094 5852 76120 5856
rect 76370 5852 76396 5878
rect 80556 5873 80582 5878
rect 80556 5856 80560 5873
rect 80560 5856 80577 5873
rect 80577 5856 80582 5873
rect 80556 5852 80582 5856
rect 80878 5873 80904 5878
rect 80878 5856 80882 5873
rect 80882 5856 80899 5873
rect 80899 5856 80904 5873
rect 80878 5852 80904 5856
rect 68872 5818 68898 5844
rect 74162 5839 74188 5844
rect 74162 5822 74166 5839
rect 74166 5822 74183 5839
rect 74183 5822 74188 5839
rect 74162 5818 74188 5822
rect 74300 5839 74326 5844
rect 74300 5822 74304 5839
rect 74304 5822 74321 5839
rect 74321 5822 74326 5839
rect 74300 5818 74326 5822
rect 71632 5784 71658 5810
rect 73012 5784 73038 5810
rect 80602 5784 80628 5810
rect 80648 5784 80674 5810
rect 81016 5920 81042 5946
rect 81384 5920 81410 5946
rect 81890 5920 81916 5946
rect 82166 5920 82192 5946
rect 82442 5941 82468 5946
rect 82442 5924 82446 5941
rect 82446 5924 82463 5941
rect 82463 5924 82468 5941
rect 82442 5920 82468 5924
rect 88376 5920 88402 5946
rect 88698 5920 88724 5946
rect 88928 5920 88954 5946
rect 89940 5920 89966 5946
rect 89986 5920 90012 5946
rect 90078 5920 90104 5946
rect 94172 5920 94198 5946
rect 95874 5920 95900 5946
rect 95920 5920 95946 5946
rect 81292 5886 81318 5912
rect 94770 5886 94796 5912
rect 96932 5886 96958 5912
rect 81844 5873 81870 5878
rect 81844 5856 81848 5873
rect 81848 5856 81865 5873
rect 81865 5856 81870 5873
rect 81844 5852 81870 5856
rect 81752 5818 81778 5844
rect 83316 5852 83342 5878
rect 88330 5873 88356 5878
rect 88330 5856 88334 5873
rect 88334 5856 88351 5873
rect 88351 5856 88356 5873
rect 88330 5852 88356 5856
rect 89940 5852 89966 5878
rect 88560 5818 88586 5844
rect 82948 5784 82974 5810
rect 15696 5771 15722 5776
rect 15696 5754 15700 5771
rect 15700 5754 15717 5771
rect 15717 5754 15722 5771
rect 15696 5750 15722 5754
rect 16478 5750 16504 5776
rect 27748 5750 27774 5776
rect 42422 5750 42448 5776
rect 43204 5750 43230 5776
rect 50932 5750 50958 5776
rect 52036 5750 52062 5776
rect 57004 5750 57030 5776
rect 65928 5771 65954 5776
rect 65928 5754 65932 5771
rect 65932 5754 65949 5771
rect 65949 5754 65954 5771
rect 65928 5750 65954 5754
rect 73656 5750 73682 5776
rect 75864 5750 75890 5776
rect 90032 5852 90058 5878
rect 90308 5852 90334 5878
rect 90400 5818 90426 5844
rect 90768 5818 90794 5844
rect 94816 5873 94842 5878
rect 94816 5856 94820 5873
rect 94820 5856 94837 5873
rect 94837 5856 94842 5873
rect 94816 5852 94842 5856
rect 95414 5852 95440 5878
rect 95920 5873 95946 5878
rect 95920 5856 95924 5873
rect 95924 5856 95941 5873
rect 95941 5856 95946 5873
rect 95920 5852 95946 5856
rect 97208 5920 97234 5946
rect 97346 5920 97372 5946
rect 101440 5941 101466 5946
rect 101440 5924 101444 5941
rect 101444 5924 101461 5941
rect 101461 5924 101466 5941
rect 101440 5920 101466 5924
rect 102268 5920 102294 5946
rect 103280 5920 103306 5946
rect 113906 5920 113932 5946
rect 114412 5920 114438 5946
rect 98404 5886 98430 5912
rect 101578 5886 101604 5912
rect 102774 5886 102800 5912
rect 113860 5886 113886 5912
rect 114964 5920 114990 5946
rect 115194 5941 115220 5946
rect 115194 5924 115198 5941
rect 115198 5924 115215 5941
rect 115215 5924 115220 5941
rect 115194 5920 115220 5924
rect 115516 5920 115542 5946
rect 115838 5920 115864 5946
rect 120162 5941 120188 5946
rect 120162 5924 120166 5941
rect 120166 5924 120183 5941
rect 120183 5924 120188 5941
rect 120162 5920 120188 5924
rect 120530 5941 120556 5946
rect 120530 5924 120534 5941
rect 120534 5924 120551 5941
rect 120551 5924 120556 5941
rect 120530 5920 120556 5924
rect 120898 5941 120924 5946
rect 120898 5924 120902 5941
rect 120902 5924 120919 5941
rect 120919 5924 120924 5941
rect 120898 5920 120924 5924
rect 126464 5920 126490 5946
rect 127338 5920 127364 5946
rect 127384 5920 127410 5946
rect 127522 5920 127548 5946
rect 133410 5920 133436 5946
rect 98956 5852 98982 5878
rect 100520 5852 100546 5878
rect 101532 5873 101558 5878
rect 101532 5856 101536 5873
rect 101536 5856 101553 5873
rect 101553 5856 101558 5873
rect 101532 5852 101558 5856
rect 96058 5839 96084 5844
rect 96058 5822 96062 5839
rect 96062 5822 96079 5839
rect 96079 5822 96084 5839
rect 96058 5818 96084 5822
rect 97162 5839 97188 5844
rect 97162 5822 97166 5839
rect 97166 5822 97183 5839
rect 97183 5822 97188 5839
rect 97162 5818 97188 5822
rect 97208 5818 97234 5844
rect 90170 5784 90196 5810
rect 98680 5818 98706 5844
rect 100658 5818 100684 5844
rect 101440 5818 101466 5844
rect 103188 5852 103214 5878
rect 115424 5886 115450 5912
rect 114688 5852 114714 5878
rect 120070 5886 120096 5912
rect 101762 5818 101788 5844
rect 103924 5818 103950 5844
rect 113630 5818 113656 5844
rect 90262 5750 90288 5776
rect 94724 5771 94750 5776
rect 94724 5754 94728 5771
rect 94728 5754 94745 5771
rect 94745 5754 94750 5771
rect 94724 5750 94750 5754
rect 98726 5784 98752 5810
rect 101716 5784 101742 5810
rect 102452 5784 102478 5810
rect 115148 5784 115174 5810
rect 96656 5750 96682 5776
rect 96748 5750 96774 5776
rect 97898 5750 97924 5776
rect 97944 5750 97970 5776
rect 98496 5750 98522 5776
rect 100750 5750 100776 5776
rect 102406 5771 102432 5776
rect 102406 5754 102410 5771
rect 102410 5754 102427 5771
rect 102427 5754 102432 5771
rect 102406 5750 102432 5754
rect 114688 5750 114714 5776
rect 115608 5852 115634 5878
rect 120760 5886 120786 5912
rect 119656 5818 119682 5844
rect 119978 5818 120004 5844
rect 116068 5784 116094 5810
rect 121266 5873 121292 5878
rect 121266 5856 121270 5873
rect 121270 5856 121287 5873
rect 121287 5856 121292 5873
rect 121266 5852 121292 5856
rect 120990 5818 121016 5844
rect 122416 5886 122442 5912
rect 127154 5886 127180 5912
rect 135342 5920 135368 5946
rect 135388 5920 135414 5946
rect 134146 5886 134172 5912
rect 134928 5886 134954 5912
rect 126004 5873 126030 5878
rect 126004 5856 126008 5873
rect 126008 5856 126025 5873
rect 126025 5856 126030 5873
rect 126004 5852 126030 5856
rect 126372 5873 126398 5878
rect 126372 5856 126376 5873
rect 126376 5856 126393 5873
rect 126393 5856 126398 5873
rect 126372 5852 126398 5856
rect 126510 5852 126536 5878
rect 128120 5852 128146 5878
rect 128626 5852 128652 5878
rect 132168 5873 132194 5878
rect 132168 5856 132172 5873
rect 132172 5856 132189 5873
rect 132189 5856 132194 5873
rect 132168 5852 132194 5856
rect 132582 5873 132608 5878
rect 132582 5856 132586 5873
rect 132586 5856 132603 5873
rect 132603 5856 132608 5873
rect 132582 5852 132608 5856
rect 132628 5852 132654 5878
rect 121358 5818 121384 5844
rect 122278 5818 122304 5844
rect 126050 5818 126076 5844
rect 127798 5818 127824 5844
rect 128212 5818 128238 5844
rect 131984 5818 132010 5844
rect 134238 5852 134264 5878
rect 134560 5873 134586 5878
rect 134560 5856 134564 5873
rect 134564 5856 134581 5873
rect 134581 5856 134586 5873
rect 134560 5852 134586 5856
rect 135664 5873 135690 5878
rect 135664 5856 135668 5873
rect 135668 5856 135685 5873
rect 135685 5856 135690 5873
rect 135664 5852 135690 5856
rect 115838 5750 115864 5776
rect 119702 5750 119728 5776
rect 120622 5750 120648 5776
rect 125820 5784 125846 5810
rect 124532 5750 124558 5776
rect 126648 5750 126674 5776
rect 134008 5784 134034 5810
rect 130880 5750 130906 5776
rect 131340 5750 131366 5776
rect 133134 5750 133160 5776
rect 133180 5750 133206 5776
rect 134698 5839 134724 5844
rect 134698 5822 134702 5839
rect 134702 5822 134719 5839
rect 134719 5822 134724 5839
rect 134698 5818 134724 5822
rect 134974 5818 135000 5844
rect 136584 5818 136610 5844
rect 137550 5750 137576 5776
rect 19524 5699 19550 5725
rect 19556 5699 19582 5725
rect 19588 5699 19614 5725
rect 19620 5699 19646 5725
rect 19652 5699 19678 5725
rect 57623 5699 57649 5725
rect 57655 5699 57681 5725
rect 57687 5699 57713 5725
rect 57719 5699 57745 5725
rect 57751 5699 57777 5725
rect 95722 5699 95748 5725
rect 95754 5699 95780 5725
rect 95786 5699 95812 5725
rect 95818 5699 95844 5725
rect 95850 5699 95876 5725
rect 133821 5699 133847 5725
rect 133853 5699 133879 5725
rect 133885 5699 133911 5725
rect 133917 5699 133943 5725
rect 133949 5699 133975 5725
rect 14960 5648 14986 5674
rect 15006 5648 15032 5674
rect 14454 5614 14480 5640
rect 16202 5648 16228 5674
rect 16662 5648 16688 5674
rect 16800 5669 16826 5674
rect 16800 5652 16804 5669
rect 16804 5652 16821 5669
rect 16821 5652 16826 5669
rect 16800 5648 16826 5652
rect 20204 5648 20230 5674
rect 20526 5669 20552 5674
rect 20526 5652 20530 5669
rect 20530 5652 20547 5669
rect 20547 5652 20552 5669
rect 20526 5648 20552 5652
rect 20802 5669 20828 5674
rect 20802 5652 20806 5669
rect 20806 5652 20823 5669
rect 20823 5652 20828 5669
rect 20802 5648 20828 5652
rect 27518 5648 27544 5674
rect 28852 5648 28878 5674
rect 38190 5648 38216 5674
rect 39386 5648 39412 5674
rect 42238 5648 42264 5674
rect 43572 5648 43598 5674
rect 44538 5648 44564 5674
rect 51438 5669 51464 5674
rect 51438 5652 51442 5669
rect 51442 5652 51459 5669
rect 51459 5652 51464 5669
rect 51438 5648 51464 5652
rect 57556 5648 57582 5674
rect 58844 5648 58870 5674
rect 65192 5648 65218 5674
rect 65606 5669 65632 5674
rect 65606 5652 65610 5669
rect 65610 5652 65627 5669
rect 65627 5652 65632 5669
rect 65606 5648 65632 5652
rect 66434 5648 66460 5674
rect 74024 5669 74050 5674
rect 74024 5652 74028 5669
rect 74028 5652 74045 5669
rect 74045 5652 74050 5669
rect 74024 5648 74050 5652
rect 75404 5669 75430 5674
rect 75404 5652 75408 5669
rect 75408 5652 75425 5669
rect 75425 5652 75430 5669
rect 75404 5648 75430 5652
rect 78624 5648 78650 5674
rect 81062 5648 81088 5674
rect 81338 5669 81364 5674
rect 81338 5652 81342 5669
rect 81342 5652 81359 5669
rect 81359 5652 81364 5669
rect 81338 5648 81364 5652
rect 81706 5648 81732 5674
rect 82948 5648 82974 5674
rect 119702 5648 119728 5674
rect 119886 5648 119912 5674
rect 120024 5648 120050 5674
rect 120484 5648 120510 5674
rect 121036 5648 121062 5674
rect 126234 5648 126260 5674
rect 126556 5669 126582 5674
rect 126556 5652 126560 5669
rect 126560 5652 126577 5669
rect 126577 5652 126582 5669
rect 126556 5648 126582 5652
rect 127016 5648 127042 5674
rect 132720 5648 132746 5674
rect 133134 5648 133160 5674
rect 13534 5580 13560 5606
rect 14730 5580 14756 5606
rect 14776 5580 14802 5606
rect 18226 5614 18252 5640
rect 20664 5614 20690 5640
rect 43388 5614 43414 5640
rect 51116 5614 51142 5640
rect 57096 5614 57122 5640
rect 73702 5614 73728 5640
rect 15696 5580 15722 5606
rect 16156 5601 16182 5606
rect 16156 5584 16160 5601
rect 16160 5584 16177 5601
rect 16177 5584 16182 5601
rect 16156 5580 16182 5584
rect 13810 5546 13836 5572
rect 16110 5567 16136 5572
rect 16110 5550 16114 5567
rect 16114 5550 16131 5567
rect 16131 5550 16136 5567
rect 16110 5546 16136 5550
rect 13994 5512 14020 5538
rect 14960 5533 14986 5538
rect 14960 5516 14964 5533
rect 14964 5516 14981 5533
rect 14981 5516 14986 5533
rect 14960 5512 14986 5516
rect 15834 5512 15860 5538
rect 15880 5512 15906 5538
rect 16294 5580 16320 5606
rect 17352 5546 17378 5572
rect 20250 5567 20276 5572
rect 20250 5550 20254 5567
rect 20254 5550 20271 5567
rect 20271 5550 20276 5567
rect 20250 5546 20276 5550
rect 20710 5546 20736 5572
rect 22504 5580 22530 5606
rect 42744 5580 42770 5606
rect 21216 5567 21242 5572
rect 21216 5550 21220 5567
rect 21220 5550 21237 5567
rect 21237 5550 21242 5567
rect 21216 5546 21242 5550
rect 27748 5567 27774 5572
rect 27748 5550 27752 5567
rect 27752 5550 27769 5567
rect 27769 5550 27774 5567
rect 27748 5546 27774 5550
rect 28622 5546 28648 5572
rect 37362 5546 37388 5572
rect 39202 5567 39228 5572
rect 39202 5550 39206 5567
rect 39206 5550 39223 5567
rect 39223 5550 39228 5567
rect 39202 5546 39228 5550
rect 43204 5567 43230 5572
rect 43204 5550 43208 5567
rect 43208 5550 43225 5567
rect 43225 5550 43230 5567
rect 43204 5546 43230 5550
rect 44584 5580 44610 5606
rect 51024 5580 51050 5606
rect 51300 5580 51326 5606
rect 43894 5567 43920 5572
rect 43894 5550 43898 5567
rect 43898 5550 43915 5567
rect 43915 5550 43920 5567
rect 43894 5546 43920 5550
rect 44216 5567 44242 5572
rect 44216 5550 44220 5567
rect 44220 5550 44237 5567
rect 44237 5550 44242 5567
rect 44216 5546 44242 5550
rect 51208 5546 51234 5572
rect 51530 5567 51556 5572
rect 51530 5550 51534 5567
rect 51534 5550 51551 5567
rect 51551 5550 51556 5567
rect 51530 5546 51556 5550
rect 65146 5580 65172 5606
rect 57372 5546 57398 5572
rect 57878 5546 57904 5572
rect 57924 5546 57950 5572
rect 59856 5546 59882 5572
rect 65468 5546 65494 5572
rect 66296 5580 66322 5606
rect 71632 5580 71658 5606
rect 66572 5546 66598 5572
rect 71034 5567 71060 5572
rect 71034 5550 71038 5567
rect 71038 5550 71055 5567
rect 71055 5550 71060 5567
rect 71034 5546 71060 5550
rect 72874 5546 72900 5572
rect 73748 5580 73774 5606
rect 78210 5614 78236 5640
rect 82718 5614 82744 5640
rect 75680 5580 75706 5606
rect 40812 5512 40838 5538
rect 43940 5512 43966 5538
rect 56866 5512 56892 5538
rect 70344 5512 70370 5538
rect 76554 5546 76580 5572
rect 81108 5567 81134 5572
rect 81108 5550 81112 5567
rect 81112 5550 81129 5567
rect 81129 5550 81134 5567
rect 81108 5546 81134 5550
rect 82672 5580 82698 5606
rect 88836 5580 88862 5606
rect 88974 5580 89000 5606
rect 81752 5567 81778 5572
rect 81752 5550 81756 5567
rect 81756 5550 81773 5567
rect 81773 5550 81778 5567
rect 81752 5546 81778 5550
rect 89020 5546 89046 5572
rect 90400 5580 90426 5606
rect 95598 5580 95624 5606
rect 95920 5580 95946 5606
rect 126372 5614 126398 5640
rect 126602 5614 126628 5640
rect 132582 5614 132608 5640
rect 134652 5648 134678 5674
rect 96748 5580 96774 5606
rect 97208 5580 97234 5606
rect 97300 5580 97326 5606
rect 90216 5546 90242 5572
rect 94494 5546 94520 5572
rect 95322 5546 95348 5572
rect 95414 5567 95440 5572
rect 95414 5550 95418 5567
rect 95418 5550 95435 5567
rect 95435 5550 95440 5567
rect 95414 5546 95440 5550
rect 95966 5546 95992 5572
rect 97438 5546 97464 5572
rect 98220 5580 98246 5606
rect 100520 5580 100546 5606
rect 97898 5567 97924 5572
rect 15926 5499 15952 5504
rect 15926 5482 15930 5499
rect 15930 5482 15947 5499
rect 15947 5482 15952 5499
rect 15926 5478 15952 5482
rect 74530 5478 74556 5504
rect 74760 5478 74786 5504
rect 78072 5512 78098 5538
rect 89710 5512 89736 5538
rect 94724 5512 94750 5538
rect 96656 5512 96682 5538
rect 97898 5550 97902 5567
rect 97902 5550 97919 5567
rect 97919 5550 97924 5567
rect 97898 5546 97924 5550
rect 101348 5546 101374 5572
rect 101670 5580 101696 5606
rect 97208 5499 97234 5504
rect 97208 5482 97212 5499
rect 97212 5482 97229 5499
rect 97229 5482 97234 5499
rect 97208 5478 97234 5482
rect 97622 5512 97648 5538
rect 102498 5580 102524 5606
rect 119012 5580 119038 5606
rect 121358 5580 121384 5606
rect 133640 5580 133666 5606
rect 134008 5580 134034 5606
rect 102038 5512 102064 5538
rect 102452 5567 102478 5572
rect 102452 5550 102456 5567
rect 102456 5550 102473 5567
rect 102473 5550 102478 5567
rect 114688 5567 114714 5572
rect 102452 5546 102478 5550
rect 114688 5550 114692 5567
rect 114692 5550 114709 5567
rect 114709 5550 114714 5567
rect 114688 5546 114714 5550
rect 102728 5512 102754 5538
rect 115378 5512 115404 5538
rect 120438 5546 120464 5572
rect 120990 5546 121016 5572
rect 125774 5546 125800 5572
rect 126510 5546 126536 5572
rect 126648 5567 126674 5572
rect 126648 5550 126652 5567
rect 126652 5550 126669 5567
rect 126669 5550 126674 5567
rect 126648 5546 126674 5550
rect 127200 5546 127226 5572
rect 127338 5546 127364 5572
rect 132168 5546 132194 5572
rect 132444 5567 132470 5572
rect 132444 5550 132448 5567
rect 132448 5550 132465 5567
rect 132465 5550 132470 5567
rect 132444 5546 132470 5550
rect 132812 5546 132838 5572
rect 134238 5580 134264 5606
rect 134468 5580 134494 5606
rect 136124 5580 136150 5606
rect 134836 5546 134862 5572
rect 135204 5567 135230 5572
rect 135204 5550 135208 5567
rect 135208 5550 135225 5567
rect 135225 5550 135230 5567
rect 135204 5546 135230 5550
rect 135434 5546 135460 5572
rect 134146 5512 134172 5538
rect 134468 5512 134494 5538
rect 134974 5512 135000 5538
rect 134422 5499 134448 5504
rect 134422 5482 134426 5499
rect 134426 5482 134443 5499
rect 134443 5482 134448 5499
rect 134422 5478 134448 5482
rect 135020 5499 135046 5504
rect 135020 5482 135024 5499
rect 135024 5482 135041 5499
rect 135041 5482 135046 5499
rect 135020 5478 135046 5482
rect 38574 5427 38600 5453
rect 38606 5427 38632 5453
rect 38638 5427 38664 5453
rect 38670 5427 38696 5453
rect 38702 5427 38728 5453
rect 76673 5427 76699 5453
rect 76705 5427 76731 5453
rect 76737 5427 76763 5453
rect 76769 5427 76795 5453
rect 76801 5427 76827 5453
rect 114772 5427 114798 5453
rect 114804 5427 114830 5453
rect 114836 5427 114862 5453
rect 114868 5427 114894 5453
rect 114900 5427 114926 5453
rect 14914 5376 14940 5402
rect 15236 5376 15262 5402
rect 15374 5397 15400 5402
rect 15374 5380 15378 5397
rect 15378 5380 15395 5397
rect 15395 5380 15400 5397
rect 15374 5376 15400 5380
rect 14868 5342 14894 5368
rect 14224 5308 14250 5334
rect 15098 5342 15124 5368
rect 16340 5376 16366 5402
rect 16524 5376 16550 5402
rect 50840 5397 50866 5402
rect 50840 5380 50844 5397
rect 50844 5380 50861 5397
rect 50861 5380 50866 5397
rect 50840 5376 50866 5380
rect 65238 5397 65264 5402
rect 65238 5380 65242 5397
rect 65242 5380 65259 5397
rect 65259 5380 65264 5397
rect 65238 5376 65264 5380
rect 70988 5397 71014 5402
rect 70988 5380 70992 5397
rect 70992 5380 71009 5397
rect 71009 5380 71014 5397
rect 70988 5376 71014 5380
rect 74300 5376 74326 5402
rect 74484 5376 74510 5402
rect 95552 5376 95578 5402
rect 15880 5342 15906 5368
rect 15926 5342 15952 5368
rect 70344 5363 70370 5368
rect 16478 5329 16504 5334
rect 16478 5312 16482 5329
rect 16482 5312 16499 5329
rect 16499 5312 16504 5329
rect 16478 5308 16504 5312
rect 70344 5346 70348 5363
rect 70348 5346 70365 5363
rect 70365 5346 70370 5363
rect 70344 5342 70370 5346
rect 50932 5329 50958 5334
rect 50932 5312 50936 5329
rect 50936 5312 50953 5329
rect 50953 5312 50958 5329
rect 50932 5308 50958 5312
rect 65146 5308 65172 5334
rect 75818 5342 75844 5368
rect 78072 5363 78098 5368
rect 78072 5346 78076 5363
rect 78076 5346 78093 5363
rect 78093 5346 78098 5363
rect 78072 5342 78098 5346
rect 75174 5308 75200 5334
rect 96104 5342 96130 5368
rect 95276 5308 95302 5334
rect 96150 5308 96176 5334
rect 96610 5342 96636 5368
rect 96932 5376 96958 5402
rect 102544 5376 102570 5402
rect 127614 5376 127640 5402
rect 133272 5397 133298 5402
rect 133272 5380 133276 5397
rect 133276 5380 133293 5397
rect 133293 5380 133298 5397
rect 133272 5376 133298 5380
rect 134100 5376 134126 5402
rect 134698 5376 134724 5402
rect 97530 5342 97556 5368
rect 132444 5342 132470 5368
rect 97070 5329 97096 5334
rect 97070 5312 97074 5329
rect 97074 5312 97091 5329
rect 97091 5312 97096 5329
rect 97070 5308 97096 5312
rect 97484 5308 97510 5334
rect 102406 5308 102432 5334
rect 127476 5308 127502 5334
rect 133180 5308 133206 5334
rect 135020 5342 135046 5368
rect 93758 5295 93784 5300
rect 93758 5278 93762 5295
rect 93762 5278 93779 5295
rect 93779 5278 93784 5295
rect 93758 5274 93784 5278
rect 96058 5240 96084 5266
rect 100520 5274 100546 5300
rect 134514 5308 134540 5334
rect 135158 5308 135184 5334
rect 136262 5274 136288 5300
rect 89572 5206 89598 5232
rect 134376 5240 134402 5266
rect 101762 5206 101788 5232
rect 134790 5206 134816 5232
rect 19524 5155 19550 5181
rect 19556 5155 19582 5181
rect 19588 5155 19614 5181
rect 19620 5155 19646 5181
rect 19652 5155 19678 5181
rect 57623 5155 57649 5181
rect 57655 5155 57681 5181
rect 57687 5155 57713 5181
rect 57719 5155 57745 5181
rect 57751 5155 57777 5181
rect 95722 5155 95748 5181
rect 95754 5155 95780 5181
rect 95786 5155 95812 5181
rect 95818 5155 95844 5181
rect 95850 5155 95876 5181
rect 133821 5155 133847 5181
rect 133853 5155 133879 5181
rect 133885 5155 133911 5181
rect 133917 5155 133943 5181
rect 133949 5155 133975 5181
rect 15052 5104 15078 5130
rect 15834 5125 15860 5130
rect 15834 5108 15838 5125
rect 15838 5108 15855 5125
rect 15855 5108 15860 5125
rect 15834 5104 15860 5108
rect 16064 5104 16090 5130
rect 16662 5104 16688 5130
rect 95644 5104 95670 5130
rect 96242 5104 96268 5130
rect 133456 5104 133482 5130
rect 134284 5104 134310 5130
rect 13764 5070 13790 5096
rect 15788 5070 15814 5096
rect 81798 5036 81824 5062
rect 14730 5002 14756 5028
rect 15466 5002 15492 5028
rect 16708 5002 16734 5028
rect 16846 5002 16872 5028
rect 70344 5002 70370 5028
rect 78072 5002 78098 5028
rect 96288 5002 96314 5028
rect 97944 5036 97970 5062
rect 133870 5036 133896 5062
rect 97208 5002 97234 5028
rect 134192 5070 134218 5096
rect 134744 5070 134770 5096
rect 134422 5036 134448 5062
rect 134054 5002 134080 5028
rect 134514 5002 134540 5028
rect 134606 5023 134632 5028
rect 134606 5006 134610 5023
rect 134610 5006 134627 5023
rect 134627 5006 134632 5023
rect 134606 5002 134632 5006
rect 152224 5023 152250 5028
rect 152224 5006 152228 5023
rect 152228 5006 152245 5023
rect 152245 5006 152250 5023
rect 152224 5002 152250 5006
rect 126372 4968 126398 4994
rect 58706 4934 58732 4960
rect 97162 4934 97188 4960
rect 133870 4934 133896 4960
rect 135480 4934 135506 4960
rect 38574 4883 38600 4909
rect 38606 4883 38632 4909
rect 38638 4883 38664 4909
rect 38670 4883 38696 4909
rect 38702 4883 38728 4909
rect 76673 4883 76699 4909
rect 76705 4883 76731 4909
rect 76737 4883 76763 4909
rect 76769 4883 76795 4909
rect 76801 4883 76827 4909
rect 114772 4883 114798 4909
rect 114804 4883 114830 4909
rect 114836 4883 114862 4909
rect 114868 4883 114894 4909
rect 114900 4883 114926 4909
rect 15604 4798 15630 4824
rect 70344 4819 70370 4824
rect 70344 4802 70348 4819
rect 70348 4802 70365 4819
rect 70365 4802 70370 4819
rect 70344 4798 70370 4802
rect 78072 4819 78098 4824
rect 78072 4802 78076 4819
rect 78076 4802 78093 4819
rect 78093 4802 78098 4819
rect 78072 4798 78098 4802
rect 79314 4798 79340 4824
rect 95322 4798 95348 4824
rect 13672 4764 13698 4790
rect 16846 4764 16872 4790
rect 96656 4798 96682 4824
rect 134928 4798 134954 4824
rect 15282 4730 15308 4756
rect 97070 4764 97096 4790
rect 134054 4764 134080 4790
rect 97990 4730 98016 4756
rect 14960 4696 14986 4722
rect 97254 4696 97280 4722
rect 52128 4662 52154 4688
rect 74162 4662 74188 4688
rect 19524 4611 19550 4637
rect 19556 4611 19582 4637
rect 19588 4611 19614 4637
rect 19620 4611 19646 4637
rect 19652 4611 19678 4637
rect 57623 4611 57649 4637
rect 57655 4611 57681 4637
rect 57687 4611 57713 4637
rect 57719 4611 57745 4637
rect 57751 4611 57777 4637
rect 95722 4611 95748 4637
rect 95754 4611 95780 4637
rect 95786 4611 95812 4637
rect 95818 4611 95844 4637
rect 95850 4611 95876 4637
rect 133821 4611 133847 4637
rect 133853 4611 133879 4637
rect 133885 4611 133911 4637
rect 133917 4611 133943 4637
rect 133949 4611 133975 4637
rect 38574 4339 38600 4365
rect 38606 4339 38632 4365
rect 38638 4339 38664 4365
rect 38670 4339 38696 4365
rect 38702 4339 38728 4365
rect 76673 4339 76699 4365
rect 76705 4339 76731 4365
rect 76737 4339 76763 4365
rect 76769 4339 76795 4365
rect 76801 4339 76827 4365
rect 114772 4339 114798 4365
rect 114804 4339 114830 4365
rect 114836 4339 114862 4365
rect 114868 4339 114894 4365
rect 114900 4339 114926 4365
rect 700 4173 726 4178
rect 700 4156 704 4173
rect 704 4156 721 4173
rect 721 4156 726 4173
rect 700 4152 726 4156
rect 93758 4152 93784 4178
rect 19524 4067 19550 4093
rect 19556 4067 19582 4093
rect 19588 4067 19614 4093
rect 19620 4067 19646 4093
rect 19652 4067 19678 4093
rect 57623 4067 57649 4093
rect 57655 4067 57681 4093
rect 57687 4067 57713 4093
rect 57719 4067 57745 4093
rect 57751 4067 57777 4093
rect 95722 4067 95748 4093
rect 95754 4067 95780 4093
rect 95786 4067 95812 4093
rect 95818 4067 95844 4093
rect 95850 4067 95876 4093
rect 133821 4067 133847 4093
rect 133853 4067 133879 4093
rect 133885 4067 133911 4093
rect 133917 4067 133943 4093
rect 133949 4067 133975 4093
rect 38574 3795 38600 3821
rect 38606 3795 38632 3821
rect 38638 3795 38664 3821
rect 38670 3795 38696 3821
rect 38702 3795 38728 3821
rect 76673 3795 76699 3821
rect 76705 3795 76731 3821
rect 76737 3795 76763 3821
rect 76769 3795 76795 3821
rect 76801 3795 76827 3821
rect 114772 3795 114798 3821
rect 114804 3795 114830 3821
rect 114836 3795 114862 3821
rect 114868 3795 114894 3821
rect 114900 3795 114926 3821
rect 19524 3523 19550 3549
rect 19556 3523 19582 3549
rect 19588 3523 19614 3549
rect 19620 3523 19646 3549
rect 19652 3523 19678 3549
rect 57623 3523 57649 3549
rect 57655 3523 57681 3549
rect 57687 3523 57713 3549
rect 57719 3523 57745 3549
rect 57751 3523 57777 3549
rect 95722 3523 95748 3549
rect 95754 3523 95780 3549
rect 95786 3523 95812 3549
rect 95818 3523 95844 3549
rect 95850 3523 95876 3549
rect 133821 3523 133847 3549
rect 133853 3523 133879 3549
rect 133885 3523 133911 3549
rect 133917 3523 133943 3549
rect 133949 3523 133975 3549
rect 38574 3251 38600 3277
rect 38606 3251 38632 3277
rect 38638 3251 38664 3277
rect 38670 3251 38696 3277
rect 38702 3251 38728 3277
rect 76673 3251 76699 3277
rect 76705 3251 76731 3277
rect 76737 3251 76763 3277
rect 76769 3251 76795 3277
rect 76801 3251 76827 3277
rect 114772 3251 114798 3277
rect 114804 3251 114830 3277
rect 114836 3251 114862 3277
rect 114868 3251 114894 3277
rect 114900 3251 114926 3277
rect 151994 3153 152020 3158
rect 151994 3136 151998 3153
rect 151998 3136 152015 3153
rect 152015 3136 152020 3153
rect 151994 3132 152020 3136
rect 124532 3098 124558 3124
rect 19524 2979 19550 3005
rect 19556 2979 19582 3005
rect 19588 2979 19614 3005
rect 19620 2979 19646 3005
rect 19652 2979 19678 3005
rect 57623 2979 57649 3005
rect 57655 2979 57681 3005
rect 57687 2979 57713 3005
rect 57719 2979 57745 3005
rect 57751 2979 57777 3005
rect 95722 2979 95748 3005
rect 95754 2979 95780 3005
rect 95786 2979 95812 3005
rect 95818 2979 95844 3005
rect 95850 2979 95876 3005
rect 133821 2979 133847 3005
rect 133853 2979 133879 3005
rect 133885 2979 133911 3005
rect 133917 2979 133943 3005
rect 133949 2979 133975 3005
rect 38574 2707 38600 2733
rect 38606 2707 38632 2733
rect 38638 2707 38664 2733
rect 38670 2707 38696 2733
rect 38702 2707 38728 2733
rect 76673 2707 76699 2733
rect 76705 2707 76731 2733
rect 76737 2707 76763 2733
rect 76769 2707 76795 2733
rect 76801 2707 76827 2733
rect 114772 2707 114798 2733
rect 114804 2707 114830 2733
rect 114836 2707 114862 2733
rect 114868 2707 114894 2733
rect 114900 2707 114926 2733
rect 19524 2435 19550 2461
rect 19556 2435 19582 2461
rect 19588 2435 19614 2461
rect 19620 2435 19646 2461
rect 19652 2435 19678 2461
rect 57623 2435 57649 2461
rect 57655 2435 57681 2461
rect 57687 2435 57713 2461
rect 57719 2435 57745 2461
rect 57751 2435 57777 2461
rect 95722 2435 95748 2461
rect 95754 2435 95780 2461
rect 95786 2435 95812 2461
rect 95818 2435 95844 2461
rect 95850 2435 95876 2461
rect 133821 2435 133847 2461
rect 133853 2435 133879 2461
rect 133885 2435 133911 2461
rect 133917 2435 133943 2461
rect 133949 2435 133975 2461
rect 38574 2163 38600 2189
rect 38606 2163 38632 2189
rect 38638 2163 38664 2189
rect 38670 2163 38696 2189
rect 38702 2163 38728 2189
rect 76673 2163 76699 2189
rect 76705 2163 76731 2189
rect 76737 2163 76763 2189
rect 76769 2163 76795 2189
rect 76801 2163 76827 2189
rect 114772 2163 114798 2189
rect 114804 2163 114830 2189
rect 114836 2163 114862 2189
rect 114868 2163 114894 2189
rect 114900 2163 114926 2189
rect 19524 1891 19550 1917
rect 19556 1891 19582 1917
rect 19588 1891 19614 1917
rect 19620 1891 19646 1917
rect 19652 1891 19678 1917
rect 57623 1891 57649 1917
rect 57655 1891 57681 1917
rect 57687 1891 57713 1917
rect 57719 1891 57745 1917
rect 57751 1891 57777 1917
rect 95722 1891 95748 1917
rect 95754 1891 95780 1917
rect 95786 1891 95812 1917
rect 95818 1891 95844 1917
rect 95850 1891 95876 1917
rect 133821 1891 133847 1917
rect 133853 1891 133879 1917
rect 133885 1891 133911 1917
rect 133917 1891 133943 1917
rect 133949 1891 133975 1917
rect 38574 1619 38600 1645
rect 38606 1619 38632 1645
rect 38638 1619 38664 1645
rect 38670 1619 38696 1645
rect 38702 1619 38728 1645
rect 76673 1619 76699 1645
rect 76705 1619 76731 1645
rect 76737 1619 76763 1645
rect 76769 1619 76795 1645
rect 76801 1619 76827 1645
rect 114772 1619 114798 1645
rect 114804 1619 114830 1645
rect 114836 1619 114862 1645
rect 114868 1619 114894 1645
rect 114900 1619 114926 1645
rect 19524 1347 19550 1373
rect 19556 1347 19582 1373
rect 19588 1347 19614 1373
rect 19620 1347 19646 1373
rect 19652 1347 19678 1373
rect 57623 1347 57649 1373
rect 57655 1347 57681 1373
rect 57687 1347 57713 1373
rect 57719 1347 57745 1373
rect 57751 1347 57777 1373
rect 95722 1347 95748 1373
rect 95754 1347 95780 1373
rect 95786 1347 95812 1373
rect 95818 1347 95844 1373
rect 95850 1347 95876 1373
rect 133821 1347 133847 1373
rect 133853 1347 133879 1373
rect 133885 1347 133911 1373
rect 133917 1347 133943 1373
rect 133949 1347 133975 1373
rect 74714 1296 74740 1322
rect 151120 1296 151146 1322
rect 38574 1075 38600 1101
rect 38606 1075 38632 1101
rect 38638 1075 38664 1101
rect 38670 1075 38696 1101
rect 38702 1075 38728 1101
rect 76673 1075 76699 1101
rect 76705 1075 76731 1101
rect 76737 1075 76763 1101
rect 76769 1075 76795 1101
rect 76801 1075 76827 1101
rect 114772 1075 114798 1101
rect 114804 1075 114830 1101
rect 114836 1075 114862 1101
rect 114868 1075 114894 1101
rect 114900 1075 114926 1101
<< metal2 >>
rect 745 7657 773 8000
rect 2263 7657 2291 8000
rect 3781 7657 3809 8000
rect 5345 7657 5373 8000
rect 745 7643 812 7657
rect 745 7600 773 7643
rect 798 6765 812 7643
rect 2263 7643 2330 7657
rect 2263 7600 2291 7643
rect 2316 6765 2330 7643
rect 3781 7643 3848 7657
rect 3781 7600 3809 7643
rect 3834 6765 3848 7643
rect 5345 7643 5412 7657
rect 5345 7600 5373 7643
rect 5398 6765 5412 7643
rect 6863 7600 6891 8000
rect 8381 7657 8409 8000
rect 9945 7657 9973 8000
rect 11463 7657 11491 8000
rect 12981 7657 13009 8000
rect 8381 7643 8448 7657
rect 8381 7600 8409 7643
rect 792 6762 818 6765
rect 792 6733 818 6736
rect 2310 6762 2336 6765
rect 2310 6733 2336 6736
rect 3828 6762 3854 6765
rect 3828 6733 3854 6736
rect 5392 6762 5418 6765
rect 6870 6756 6884 7600
rect 8434 6765 8448 7643
rect 9945 7643 10012 7657
rect 9945 7600 9973 7643
rect 9998 6765 10012 7643
rect 11463 7643 11530 7657
rect 11463 7600 11491 7643
rect 11516 6765 11530 7643
rect 12981 7643 13048 7657
rect 12981 7600 13009 7643
rect 6910 6762 6936 6765
rect 6870 6742 6910 6756
rect 5392 6733 5418 6736
rect 6910 6733 6936 6736
rect 8428 6762 8454 6765
rect 8428 6733 8454 6736
rect 9992 6762 10018 6765
rect 9992 6733 10018 6736
rect 11510 6762 11536 6765
rect 11510 6733 11536 6736
rect 2402 6660 2428 6663
rect 2402 6631 2428 6634
rect 7140 6660 7166 6663
rect 7140 6631 7166 6634
rect 8520 6660 8546 6663
rect 8520 6631 8546 6634
rect 10084 6660 10110 6663
rect 10084 6631 10110 6634
rect 11602 6660 11628 6663
rect 11602 6631 11628 6634
rect 2408 6051 2422 6631
rect 7146 6187 7160 6631
rect 7140 6184 7166 6187
rect 7140 6155 7166 6158
rect 8526 6119 8540 6631
rect 10090 6459 10104 6631
rect 10084 6456 10110 6459
rect 10084 6427 10110 6430
rect 11608 6391 11622 6631
rect 13034 6493 13048 7643
rect 14545 7600 14573 8000
rect 16063 7600 16091 8000
rect 17627 7657 17655 8000
rect 19145 7657 19173 8000
rect 17627 7643 17786 7657
rect 17627 7600 17655 7643
rect 14500 6898 14526 6901
rect 14500 6869 14526 6872
rect 13580 6864 13606 6867
rect 13580 6835 13606 6838
rect 13586 6731 13600 6835
rect 13724 6827 13876 6841
rect 13580 6728 13606 6731
rect 13580 6699 13606 6702
rect 13488 6694 13514 6697
rect 13488 6665 13514 6668
rect 13028 6490 13054 6493
rect 13028 6461 13054 6464
rect 11602 6388 11628 6391
rect 11602 6359 11628 6362
rect 13494 6221 13508 6665
rect 13586 6357 13600 6699
rect 13626 6592 13652 6595
rect 13626 6563 13652 6566
rect 13632 6501 13646 6563
rect 13724 6501 13738 6827
rect 13862 6765 13876 6827
rect 13810 6762 13836 6765
rect 13810 6733 13836 6736
rect 13856 6762 13882 6765
rect 13856 6733 13882 6736
rect 13764 6626 13790 6629
rect 13764 6597 13790 6600
rect 13632 6487 13738 6501
rect 13672 6456 13698 6459
rect 13672 6427 13698 6430
rect 13580 6354 13606 6357
rect 13580 6325 13606 6328
rect 13488 6218 13514 6221
rect 13488 6189 13514 6192
rect 13442 6150 13468 6153
rect 13442 6121 13468 6124
rect 8520 6116 8546 6119
rect 8520 6087 8546 6090
rect 13448 6093 13462 6121
rect 13448 6079 13600 6093
rect 13586 6051 13600 6079
rect 2402 6048 2428 6051
rect 2402 6019 2428 6022
rect 13534 6048 13560 6051
rect 13534 6019 13560 6022
rect 13580 6048 13606 6051
rect 13580 6019 13606 6022
rect 13540 5609 13554 6019
rect 13534 5606 13560 5609
rect 13534 5577 13560 5580
rect 13678 4793 13692 6427
rect 13724 6119 13738 6487
rect 13718 6116 13744 6119
rect 13718 6087 13744 6090
rect 13770 5099 13784 6597
rect 13816 5575 13830 6733
rect 13856 6592 13882 6595
rect 13856 6563 13882 6566
rect 13862 5915 13876 6563
rect 14506 6459 14520 6869
rect 14500 6456 14526 6459
rect 14500 6427 14526 6430
rect 13994 6422 14020 6425
rect 13994 6393 14020 6396
rect 14000 6051 14014 6393
rect 14040 6388 14066 6391
rect 14040 6359 14066 6362
rect 14046 6221 14060 6359
rect 14454 6320 14480 6323
rect 14454 6291 14480 6294
rect 14040 6218 14066 6221
rect 14040 6189 14066 6192
rect 14408 6218 14434 6221
rect 14408 6189 14434 6192
rect 14046 6153 14060 6189
rect 14414 6161 14428 6189
rect 14368 6153 14428 6161
rect 14040 6150 14066 6153
rect 14040 6121 14066 6124
rect 14362 6150 14428 6153
rect 14388 6147 14428 6150
rect 14362 6121 14388 6124
rect 13994 6048 14020 6051
rect 13994 6019 14020 6022
rect 13856 5912 13882 5915
rect 13856 5883 13882 5886
rect 13810 5572 13836 5575
rect 13810 5543 13836 5546
rect 14000 5541 14014 6019
rect 14368 5915 14382 6121
rect 14460 6051 14474 6291
rect 14500 6150 14526 6153
rect 14500 6121 14526 6124
rect 14454 6048 14480 6051
rect 14454 6019 14480 6022
rect 14506 5915 14520 6121
rect 14552 5949 14566 7600
rect 15236 6762 15262 6765
rect 15236 6733 15262 6736
rect 15242 6705 15256 6733
rect 15196 6691 15256 6705
rect 14914 6660 14940 6663
rect 14914 6631 14940 6634
rect 14920 6391 14934 6631
rect 15098 6626 15124 6629
rect 15098 6597 15124 6600
rect 14822 6388 14848 6391
rect 14822 6359 14848 6362
rect 14914 6388 14940 6391
rect 14914 6359 14940 6362
rect 15052 6388 15078 6391
rect 15052 6359 15078 6362
rect 14828 6217 14842 6359
rect 14828 6203 14888 6217
rect 14776 6150 14802 6153
rect 14776 6121 14802 6124
rect 14684 6116 14710 6119
rect 14683 6100 14684 6104
rect 14710 6100 14711 6104
rect 14683 6067 14711 6072
rect 14730 6082 14756 6085
rect 14730 6053 14756 6056
rect 14736 5949 14750 6053
rect 14546 5946 14572 5949
rect 14546 5917 14572 5920
rect 14730 5946 14756 5949
rect 14730 5917 14756 5920
rect 14362 5912 14388 5915
rect 14362 5883 14388 5886
rect 14500 5912 14526 5915
rect 14500 5883 14526 5886
rect 14782 5881 14796 6121
rect 14776 5878 14802 5881
rect 14776 5849 14802 5852
rect 14454 5844 14480 5847
rect 14454 5815 14480 5818
rect 14224 5776 14250 5779
rect 14224 5747 14250 5750
rect 13994 5538 14020 5541
rect 13994 5509 14020 5512
rect 14230 5337 14244 5747
rect 14460 5643 14474 5815
rect 14454 5640 14480 5643
rect 14454 5611 14480 5614
rect 14782 5609 14796 5849
rect 14730 5606 14756 5609
rect 14730 5577 14756 5580
rect 14776 5606 14802 5609
rect 14776 5577 14802 5580
rect 14224 5334 14250 5337
rect 14224 5305 14250 5308
rect 13764 5096 13790 5099
rect 13764 5067 13790 5070
rect 14736 5031 14750 5577
rect 14874 5371 14888 6203
rect 14914 6082 14940 6085
rect 14914 6053 14940 6056
rect 14920 5405 14934 6053
rect 15006 5912 15032 5915
rect 15006 5883 15032 5886
rect 14960 5844 14986 5847
rect 14960 5815 14986 5818
rect 14966 5677 14980 5815
rect 15012 5677 15026 5883
rect 14960 5674 14986 5677
rect 14960 5645 14986 5648
rect 15006 5674 15032 5677
rect 15006 5645 15032 5648
rect 14960 5538 14986 5541
rect 14960 5509 14986 5512
rect 14914 5402 14940 5405
rect 14914 5373 14940 5376
rect 14868 5368 14894 5371
rect 14868 5339 14894 5342
rect 14730 5028 14756 5031
rect 14730 4999 14756 5002
rect 13672 4790 13698 4793
rect 13672 4761 13698 4764
rect 14966 4725 14980 5509
rect 15058 5133 15072 6359
rect 15104 5371 15118 6597
rect 15196 6459 15210 6691
rect 15236 6592 15262 6595
rect 15236 6563 15262 6566
rect 15190 6456 15216 6459
rect 15190 6427 15216 6430
rect 15196 5685 15210 6427
rect 15242 6217 15256 6563
rect 15788 6456 15814 6459
rect 15788 6427 15814 6430
rect 15696 6320 15722 6323
rect 15696 6291 15722 6294
rect 15242 6203 15302 6217
rect 15196 5671 15256 5685
rect 15242 5405 15256 5671
rect 15236 5402 15262 5405
rect 15236 5373 15262 5376
rect 15098 5368 15124 5371
rect 15098 5339 15124 5342
rect 15052 5130 15078 5133
rect 15052 5101 15078 5104
rect 15288 4759 15302 6203
rect 15702 6104 15716 6291
rect 15373 6100 15401 6104
rect 15695 6100 15723 6104
rect 15373 6067 15401 6072
rect 15604 6082 15630 6085
rect 15380 5405 15394 6067
rect 15695 6067 15723 6072
rect 15604 6053 15630 6056
rect 15558 6048 15584 6051
rect 15558 6019 15584 6022
rect 15466 5946 15492 5949
rect 15466 5917 15492 5920
rect 15374 5402 15400 5405
rect 15374 5373 15400 5376
rect 15472 5031 15486 5917
rect 15564 5813 15578 6019
rect 15558 5810 15584 5813
rect 15558 5781 15584 5784
rect 15466 5028 15492 5031
rect 15466 4999 15492 5002
rect 15610 4827 15624 6053
rect 15696 5776 15722 5779
rect 15696 5747 15722 5750
rect 15702 5609 15716 5747
rect 15696 5606 15722 5609
rect 15696 5577 15722 5580
rect 15794 5099 15808 6427
rect 16018 6082 16044 6085
rect 16018 6053 16044 6056
rect 16024 5915 16038 6053
rect 16018 5912 16044 5915
rect 16018 5883 16044 5886
rect 15834 5538 15860 5541
rect 15834 5509 15860 5512
rect 15880 5538 15906 5541
rect 15880 5509 15906 5512
rect 15840 5133 15854 5509
rect 15886 5371 15900 5509
rect 15926 5504 15952 5507
rect 15926 5475 15952 5478
rect 15932 5371 15946 5475
rect 15880 5368 15906 5371
rect 15880 5339 15906 5342
rect 15926 5368 15952 5371
rect 15926 5339 15952 5342
rect 16070 5133 16084 7600
rect 16478 6898 16504 6901
rect 16478 6869 16504 6872
rect 16202 6660 16228 6663
rect 16202 6631 16228 6634
rect 16110 6490 16136 6493
rect 16110 6461 16136 6464
rect 16116 5949 16130 6461
rect 16208 6323 16222 6631
rect 16340 6626 16366 6629
rect 16340 6597 16366 6600
rect 16202 6320 16228 6323
rect 16202 6291 16228 6294
rect 16294 6218 16320 6221
rect 16294 6189 16320 6192
rect 16156 6048 16182 6051
rect 16156 6019 16182 6022
rect 16110 5946 16136 5949
rect 16110 5917 16136 5920
rect 16116 5575 16130 5917
rect 16162 5609 16176 6019
rect 16202 5878 16228 5881
rect 16202 5849 16228 5852
rect 16208 5677 16222 5849
rect 16300 5847 16314 6189
rect 16294 5844 16320 5847
rect 16294 5815 16320 5818
rect 16202 5674 16228 5677
rect 16202 5645 16228 5648
rect 16300 5609 16314 5815
rect 16156 5606 16182 5609
rect 16156 5577 16182 5580
rect 16294 5606 16320 5609
rect 16294 5577 16320 5580
rect 16110 5572 16136 5575
rect 16110 5543 16136 5546
rect 16346 5405 16360 6597
rect 16484 6051 16498 6869
rect 16892 6660 16918 6663
rect 16892 6631 16918 6634
rect 16800 6592 16826 6595
rect 16800 6563 16826 6566
rect 16524 6388 16550 6391
rect 16524 6359 16550 6362
rect 16708 6388 16734 6391
rect 16708 6359 16734 6362
rect 16478 6048 16504 6051
rect 16478 6019 16504 6022
rect 16478 5776 16504 5779
rect 16478 5747 16504 5750
rect 16340 5402 16366 5405
rect 16340 5373 16366 5376
rect 16484 5337 16498 5747
rect 16530 5405 16544 6359
rect 16662 5674 16688 5677
rect 16662 5645 16688 5648
rect 16524 5402 16550 5405
rect 16524 5373 16550 5376
rect 16478 5334 16504 5337
rect 16478 5305 16504 5308
rect 16668 5133 16682 5645
rect 15834 5130 15860 5133
rect 15834 5101 15860 5104
rect 16064 5130 16090 5133
rect 16064 5101 16090 5104
rect 16662 5130 16688 5133
rect 16662 5101 16688 5104
rect 15788 5096 15814 5099
rect 15788 5067 15814 5070
rect 16714 5031 16728 6359
rect 16806 5677 16820 6563
rect 16846 6422 16872 6425
rect 16846 6393 16872 6396
rect 16800 5674 16826 5677
rect 16800 5645 16826 5648
rect 16852 5031 16866 6393
rect 16898 5949 16912 6631
rect 17260 6626 17286 6629
rect 17260 6597 17286 6600
rect 17076 6592 17102 6595
rect 17076 6563 17102 6566
rect 17168 6592 17194 6595
rect 17168 6563 17194 6566
rect 17082 6493 17096 6563
rect 17076 6490 17102 6493
rect 17076 6461 17102 6464
rect 17082 6416 17096 6461
rect 17036 6402 17096 6416
rect 16892 5946 16918 5949
rect 16892 5917 16918 5920
rect 17036 5847 17050 6402
rect 17174 6391 17188 6563
rect 17214 6456 17240 6459
rect 17214 6427 17240 6430
rect 17168 6388 17194 6391
rect 17168 6359 17194 6362
rect 17076 6320 17102 6323
rect 17076 6291 17102 6294
rect 17082 6119 17096 6291
rect 17076 6116 17102 6119
rect 17076 6087 17102 6090
rect 17220 5949 17234 6427
rect 17266 6221 17280 6597
rect 17772 6493 17786 7643
rect 19145 7643 19212 7657
rect 19145 7600 19173 7643
rect 18272 6864 18298 6867
rect 18272 6835 18298 6838
rect 18278 6765 18292 6835
rect 18272 6762 18298 6765
rect 18272 6733 18298 6736
rect 17996 6626 18022 6629
rect 17996 6597 18022 6600
rect 18916 6626 18942 6629
rect 18916 6597 18942 6600
rect 17766 6490 17792 6493
rect 17766 6461 17792 6464
rect 17444 6388 17470 6391
rect 17444 6359 17470 6362
rect 17674 6388 17700 6391
rect 17674 6359 17700 6362
rect 17260 6218 17286 6221
rect 17260 6189 17286 6192
rect 17450 6187 17464 6359
rect 17444 6184 17470 6187
rect 17444 6155 17470 6158
rect 17680 6119 17694 6359
rect 18002 6221 18016 6597
rect 18732 6592 18758 6595
rect 18732 6563 18758 6566
rect 18738 6459 18752 6563
rect 18732 6456 18758 6459
rect 18732 6427 18758 6430
rect 18922 6221 18936 6597
rect 19008 6320 19034 6323
rect 19008 6291 19034 6294
rect 17996 6218 18022 6221
rect 17996 6189 18022 6192
rect 18916 6218 18942 6221
rect 18916 6189 18942 6192
rect 19014 6119 19028 6291
rect 17352 6116 17378 6119
rect 17352 6087 17378 6090
rect 17674 6116 17700 6119
rect 17674 6087 17700 6090
rect 19008 6116 19034 6119
rect 19008 6087 19034 6090
rect 17214 5946 17240 5949
rect 17214 5917 17240 5920
rect 17358 5881 17372 6087
rect 18226 6048 18252 6051
rect 18226 6019 18252 6022
rect 17352 5878 17378 5881
rect 17352 5849 17378 5852
rect 17030 5844 17056 5847
rect 17030 5815 17056 5818
rect 17358 5575 17372 5849
rect 18232 5643 18246 6019
rect 19198 5949 19212 7643
rect 20663 7600 20691 8000
rect 22227 7657 22255 8000
rect 23745 7657 23773 8000
rect 22227 7643 22294 7657
rect 22227 7600 22255 7643
rect 19524 6814 19678 6818
rect 19524 6813 19527 6814
rect 19555 6813 19567 6814
rect 19595 6813 19607 6814
rect 19635 6813 19647 6814
rect 19675 6813 19678 6814
rect 19555 6787 19556 6813
rect 19646 6787 19647 6813
rect 19524 6786 19527 6787
rect 19555 6786 19567 6787
rect 19595 6786 19607 6787
rect 19635 6786 19647 6787
rect 19675 6786 19678 6787
rect 19524 6781 19678 6786
rect 19468 6660 19494 6663
rect 19468 6631 19494 6634
rect 19474 6221 19488 6631
rect 20204 6626 20230 6629
rect 20204 6597 20230 6600
rect 19652 6592 19678 6595
rect 19652 6563 19678 6566
rect 19974 6592 20000 6595
rect 19974 6563 20000 6566
rect 19658 6425 19672 6563
rect 19836 6456 19862 6459
rect 19836 6427 19862 6430
rect 19652 6422 19678 6425
rect 19652 6393 19678 6396
rect 19698 6388 19724 6391
rect 19698 6359 19724 6362
rect 19524 6270 19678 6274
rect 19524 6269 19527 6270
rect 19555 6269 19567 6270
rect 19595 6269 19607 6270
rect 19635 6269 19647 6270
rect 19675 6269 19678 6270
rect 19555 6243 19556 6269
rect 19646 6243 19647 6269
rect 19524 6242 19527 6243
rect 19555 6242 19567 6243
rect 19595 6242 19607 6243
rect 19635 6242 19647 6243
rect 19675 6242 19678 6243
rect 19524 6237 19678 6242
rect 19704 6221 19718 6359
rect 19468 6218 19494 6221
rect 19468 6189 19494 6192
rect 19698 6218 19724 6221
rect 19698 6189 19724 6192
rect 19192 5946 19218 5949
rect 19192 5917 19218 5920
rect 19790 5946 19816 5949
rect 19842 5940 19856 6427
rect 19980 5949 19994 6563
rect 20158 6116 20184 6119
rect 20158 6087 20184 6090
rect 19816 5926 19856 5940
rect 19974 5946 20000 5949
rect 19790 5917 19816 5920
rect 19974 5917 20000 5920
rect 20164 5881 20178 6087
rect 20158 5878 20184 5881
rect 20158 5849 20184 5852
rect 19524 5726 19678 5730
rect 19524 5725 19527 5726
rect 19555 5725 19567 5726
rect 19595 5725 19607 5726
rect 19635 5725 19647 5726
rect 19675 5725 19678 5726
rect 19555 5699 19556 5725
rect 19646 5699 19647 5725
rect 19524 5698 19527 5699
rect 19555 5698 19567 5699
rect 19595 5698 19607 5699
rect 19635 5698 19647 5699
rect 19675 5698 19678 5699
rect 19524 5693 19678 5698
rect 20210 5677 20224 6597
rect 20526 6456 20552 6459
rect 20526 6427 20552 6430
rect 20480 6388 20506 6391
rect 20480 6359 20506 6362
rect 20486 6221 20500 6359
rect 20480 6218 20506 6221
rect 20480 6189 20506 6192
rect 20486 6153 20500 6189
rect 20480 6150 20506 6153
rect 20480 6121 20506 6124
rect 20296 6116 20322 6119
rect 20295 6100 20296 6104
rect 20322 6100 20323 6104
rect 20295 6067 20323 6072
rect 20250 6048 20276 6051
rect 20250 6019 20276 6022
rect 20342 6048 20368 6051
rect 20342 6019 20368 6022
rect 20204 5674 20230 5677
rect 20204 5645 20230 5648
rect 18226 5640 18252 5643
rect 18226 5611 18252 5614
rect 20256 5575 20270 6019
rect 20348 5915 20362 6019
rect 20342 5912 20368 5915
rect 20342 5883 20368 5886
rect 20486 5847 20500 6121
rect 20480 5844 20506 5847
rect 20480 5815 20506 5818
rect 20532 5677 20546 6427
rect 20618 6320 20644 6323
rect 20618 6291 20644 6294
rect 20624 5915 20638 6291
rect 20618 5912 20644 5915
rect 20618 5883 20644 5886
rect 20526 5674 20552 5677
rect 20526 5645 20552 5648
rect 20670 5643 20684 7600
rect 21262 6864 21288 6867
rect 21262 6835 21288 6838
rect 21268 6663 21282 6835
rect 22090 6728 22116 6731
rect 22182 6728 22208 6731
rect 22116 6708 22182 6722
rect 22090 6699 22116 6702
rect 22182 6699 22208 6702
rect 21262 6660 21288 6663
rect 21262 6631 21288 6634
rect 22136 6660 22162 6663
rect 22136 6631 22162 6634
rect 20710 6626 20736 6629
rect 20710 6597 20736 6600
rect 21446 6626 21472 6629
rect 21446 6597 21472 6600
rect 21630 6626 21656 6629
rect 21630 6597 21656 6600
rect 20716 5949 20730 6597
rect 21216 6592 21242 6595
rect 21216 6563 21242 6566
rect 20756 6422 20782 6425
rect 20756 6393 20782 6396
rect 20710 5946 20736 5949
rect 20710 5917 20736 5920
rect 20710 5844 20736 5847
rect 20762 5838 20776 6393
rect 20894 6320 20920 6323
rect 20894 6291 20920 6294
rect 20900 6085 20914 6291
rect 21222 6104 21236 6563
rect 21400 6320 21426 6323
rect 21400 6291 21426 6294
rect 21215 6100 21243 6104
rect 20802 6082 20828 6085
rect 20802 6053 20828 6056
rect 20894 6082 20920 6085
rect 21215 6067 21243 6072
rect 20894 6053 20920 6056
rect 20736 5824 20776 5838
rect 20710 5815 20736 5818
rect 20664 5640 20690 5643
rect 20664 5611 20690 5614
rect 20716 5575 20730 5815
rect 20808 5677 20822 6053
rect 20802 5674 20828 5677
rect 20802 5645 20828 5648
rect 21222 5575 21236 6067
rect 21406 5881 21420 6291
rect 21452 5949 21466 6597
rect 21636 6493 21650 6597
rect 22142 6493 22156 6631
rect 22280 6493 22294 7643
rect 23745 7643 23812 7657
rect 23745 7600 23773 7643
rect 23102 6898 23128 6901
rect 23102 6869 23128 6872
rect 23108 6765 23122 6869
rect 23798 6765 23812 7643
rect 25263 7600 25291 8000
rect 26827 7600 26855 8000
rect 28345 7600 28373 8000
rect 29909 7600 29937 8000
rect 31427 7657 31455 8000
rect 32945 7657 32973 8000
rect 34509 7657 34537 8000
rect 36027 7657 36055 8000
rect 31427 7643 31540 7657
rect 31427 7600 31455 7643
rect 23930 6864 23956 6867
rect 23930 6835 23956 6838
rect 23102 6762 23128 6765
rect 23102 6733 23128 6736
rect 23792 6762 23818 6765
rect 23792 6733 23818 6736
rect 22780 6694 22806 6697
rect 22780 6665 22806 6668
rect 22504 6592 22530 6595
rect 22504 6563 22530 6566
rect 22688 6592 22714 6595
rect 22688 6563 22714 6566
rect 21630 6490 21656 6493
rect 21630 6461 21656 6464
rect 22136 6490 22162 6493
rect 22136 6461 22162 6464
rect 22274 6490 22300 6493
rect 22274 6461 22300 6464
rect 21492 6456 21518 6459
rect 21492 6427 21518 6430
rect 21446 5946 21472 5949
rect 21446 5917 21472 5920
rect 21498 5881 21512 6427
rect 21544 6419 21650 6433
rect 21544 6391 21558 6419
rect 21538 6388 21564 6391
rect 21538 6359 21564 6362
rect 21584 6388 21610 6391
rect 21584 6359 21610 6362
rect 21590 6221 21604 6359
rect 21636 6323 21650 6419
rect 21906 6388 21932 6391
rect 21906 6359 21932 6362
rect 21912 6323 21926 6359
rect 21630 6320 21656 6323
rect 21630 6291 21656 6294
rect 21906 6320 21932 6323
rect 21906 6291 21932 6294
rect 21912 6221 21926 6291
rect 21584 6218 21610 6221
rect 21584 6189 21610 6192
rect 21906 6218 21932 6221
rect 21906 6189 21932 6192
rect 21860 6184 21886 6187
rect 21860 6155 21886 6158
rect 21866 6119 21880 6155
rect 21860 6116 21886 6119
rect 21860 6087 21886 6090
rect 21400 5878 21426 5881
rect 21400 5849 21426 5852
rect 21492 5878 21518 5881
rect 21492 5849 21518 5852
rect 22510 5609 22524 6563
rect 22694 6425 22708 6563
rect 22688 6422 22714 6425
rect 22688 6393 22714 6396
rect 22734 6388 22760 6391
rect 22786 6382 22800 6665
rect 23936 6629 23950 6835
rect 25270 6765 25284 7600
rect 25816 6864 25842 6867
rect 25816 6835 25842 6838
rect 25264 6762 25290 6765
rect 25264 6733 25290 6736
rect 25822 6697 25836 6835
rect 26506 6762 26532 6765
rect 26506 6733 26532 6736
rect 25816 6694 25842 6697
rect 25816 6665 25842 6668
rect 25678 6660 25704 6663
rect 25678 6631 25704 6634
rect 23930 6626 23956 6629
rect 23930 6597 23956 6600
rect 25684 6391 25698 6631
rect 22760 6368 22800 6382
rect 25678 6388 25704 6391
rect 22734 6359 22760 6362
rect 25678 6359 25704 6362
rect 26322 6082 26348 6085
rect 26322 6053 26348 6056
rect 26328 5949 26342 6053
rect 26322 5946 26348 5949
rect 26322 5917 26348 5920
rect 26512 5881 26526 6733
rect 26644 6626 26670 6629
rect 26644 6597 26670 6600
rect 26650 6493 26664 6597
rect 26644 6490 26670 6493
rect 26644 6461 26670 6464
rect 26552 6320 26578 6323
rect 26552 6291 26578 6294
rect 26558 6085 26572 6291
rect 26552 6082 26578 6085
rect 26552 6053 26578 6056
rect 26834 5949 26848 7600
rect 27058 6864 27084 6867
rect 27058 6835 27084 6838
rect 26874 6422 26900 6425
rect 26874 6393 26900 6396
rect 27012 6422 27038 6425
rect 27012 6393 27038 6396
rect 26880 6161 26894 6393
rect 27018 6221 27032 6393
rect 27064 6391 27078 6835
rect 27794 6762 27820 6765
rect 27794 6733 27820 6736
rect 27800 6663 27814 6733
rect 27196 6660 27222 6663
rect 27196 6631 27222 6634
rect 27380 6660 27406 6663
rect 27380 6631 27406 6634
rect 27794 6660 27820 6663
rect 27794 6631 27820 6634
rect 27058 6388 27084 6391
rect 27058 6359 27084 6362
rect 27064 6323 27078 6359
rect 27058 6320 27084 6323
rect 27058 6291 27084 6294
rect 27012 6218 27038 6221
rect 27012 6189 27038 6192
rect 26880 6153 26940 6161
rect 26880 6150 26946 6153
rect 26880 6147 26920 6150
rect 26828 5946 26854 5949
rect 26828 5917 26854 5920
rect 26880 5915 26894 6147
rect 26920 6121 26946 6124
rect 27202 5949 27216 6631
rect 27334 6592 27360 6595
rect 27334 6563 27360 6566
rect 27340 6493 27354 6563
rect 27334 6490 27360 6493
rect 27334 6461 27360 6464
rect 27196 5946 27222 5949
rect 27196 5917 27222 5920
rect 26874 5912 26900 5915
rect 26874 5883 26900 5886
rect 26506 5878 26532 5881
rect 26506 5849 26532 5852
rect 27340 5847 27354 6461
rect 27386 6425 27400 6631
rect 27932 6626 27958 6629
rect 27932 6597 27958 6600
rect 28300 6626 28326 6629
rect 28300 6597 28326 6600
rect 27938 6493 27952 6597
rect 27932 6490 27958 6493
rect 27932 6461 27958 6464
rect 27748 6456 27774 6459
rect 27748 6427 27774 6430
rect 27380 6422 27406 6425
rect 27380 6393 27406 6396
rect 27518 6388 27544 6391
rect 27518 6359 27544 6362
rect 27334 5844 27360 5847
rect 27334 5815 27360 5818
rect 27524 5677 27538 6359
rect 27754 6221 27768 6427
rect 27794 6320 27820 6323
rect 27794 6291 27820 6294
rect 28162 6320 28188 6323
rect 28162 6291 28188 6294
rect 28254 6320 28280 6323
rect 28254 6291 28280 6294
rect 27748 6218 27774 6221
rect 27748 6189 27774 6192
rect 27656 6116 27682 6119
rect 27656 6087 27682 6090
rect 27662 5949 27676 6087
rect 27656 5946 27682 5949
rect 27656 5917 27682 5920
rect 27800 5847 27814 6291
rect 28168 6217 28182 6291
rect 28168 6203 28228 6217
rect 28214 6153 28228 6203
rect 28208 6150 28234 6153
rect 28208 6121 28234 6124
rect 28260 6119 28274 6291
rect 28254 6116 28280 6119
rect 28254 6087 28280 6090
rect 27932 6048 27958 6051
rect 27932 6019 27958 6022
rect 28024 6048 28050 6051
rect 28024 6019 28050 6022
rect 27938 5847 27952 6019
rect 27794 5844 27820 5847
rect 27794 5815 27820 5818
rect 27932 5844 27958 5847
rect 27932 5815 27958 5818
rect 28030 5813 28044 6019
rect 28306 5949 28320 6597
rect 28352 6221 28366 7600
rect 28944 6762 28970 6765
rect 28944 6733 28970 6736
rect 28950 6663 28964 6733
rect 29916 6731 29930 7600
rect 30876 6762 30902 6765
rect 30876 6733 30902 6736
rect 29910 6728 29936 6731
rect 29910 6699 29936 6702
rect 28944 6660 28970 6663
rect 28944 6631 28970 6634
rect 30324 6660 30350 6663
rect 30324 6631 30350 6634
rect 28852 6626 28878 6629
rect 28852 6597 28878 6600
rect 29312 6626 29338 6629
rect 29312 6597 29338 6600
rect 28668 6592 28694 6595
rect 28668 6563 28694 6566
rect 28674 6459 28688 6563
rect 28668 6456 28694 6459
rect 28668 6427 28694 6430
rect 28622 6320 28648 6323
rect 28622 6291 28648 6294
rect 28346 6218 28372 6221
rect 28346 6189 28372 6192
rect 28300 5946 28326 5949
rect 28300 5917 28326 5920
rect 28024 5810 28050 5813
rect 28024 5781 28050 5784
rect 27748 5776 27774 5779
rect 27748 5747 27774 5750
rect 27518 5674 27544 5677
rect 27518 5645 27544 5648
rect 22504 5606 22530 5609
rect 22504 5577 22530 5580
rect 27754 5575 27768 5747
rect 28628 5575 28642 6291
rect 28674 6051 28688 6427
rect 28714 6422 28740 6425
rect 28714 6393 28740 6396
rect 28668 6048 28694 6051
rect 28668 6019 28694 6022
rect 28720 5915 28734 6393
rect 28714 5912 28740 5915
rect 28714 5883 28740 5886
rect 28858 5677 28872 6597
rect 28990 6490 29016 6493
rect 28990 6461 29016 6464
rect 28996 6221 29010 6461
rect 28990 6218 29016 6221
rect 28990 6189 29016 6192
rect 29318 5949 29332 6597
rect 29818 6592 29844 6595
rect 29818 6563 29844 6566
rect 29824 6493 29838 6563
rect 29818 6490 29844 6493
rect 29818 6461 29844 6464
rect 30330 6459 30344 6631
rect 30744 6629 30850 6637
rect 30882 6629 30896 6733
rect 31526 6731 31540 7643
rect 32945 7643 33012 7657
rect 32945 7600 32973 7643
rect 31704 6898 31730 6901
rect 31704 6869 31730 6872
rect 31710 6765 31724 6869
rect 31704 6762 31730 6765
rect 31704 6733 31730 6736
rect 31520 6728 31546 6731
rect 31520 6699 31546 6702
rect 30738 6626 30850 6629
rect 30764 6623 30850 6626
rect 30738 6597 30764 6600
rect 30836 6595 30850 6623
rect 30876 6626 30902 6629
rect 30876 6597 30902 6600
rect 32998 6595 33012 7643
rect 34509 7643 34576 7657
rect 34509 7600 34537 7643
rect 33084 6864 33110 6867
rect 33084 6835 33110 6838
rect 33090 6663 33104 6835
rect 33084 6660 33110 6663
rect 33084 6631 33110 6634
rect 34562 6595 34576 7643
rect 36027 7643 36094 7657
rect 36027 7600 36055 7643
rect 34648 6898 34674 6901
rect 34648 6869 34674 6872
rect 34654 6663 34668 6869
rect 34648 6660 34674 6663
rect 34648 6631 34674 6634
rect 30830 6592 30856 6595
rect 30830 6563 30856 6566
rect 32946 6592 32972 6595
rect 32946 6563 32972 6566
rect 32992 6592 33018 6595
rect 32992 6563 33018 6566
rect 34556 6592 34582 6595
rect 34556 6563 34582 6566
rect 32952 6459 32966 6563
rect 36080 6493 36094 7643
rect 37545 7600 37573 8000
rect 39109 7657 39137 8000
rect 40627 7657 40655 8000
rect 39109 7643 39268 7657
rect 39109 7600 39137 7643
rect 36212 6864 36238 6867
rect 36212 6835 36238 6838
rect 36948 6864 36974 6867
rect 36948 6835 36974 6838
rect 36218 6595 36232 6835
rect 36350 6694 36376 6697
rect 36350 6665 36376 6668
rect 36166 6592 36192 6595
rect 36166 6563 36192 6566
rect 36212 6592 36238 6595
rect 36212 6563 36238 6566
rect 36172 6493 36186 6563
rect 36074 6490 36100 6493
rect 36074 6461 36100 6464
rect 36166 6490 36192 6493
rect 36166 6461 36192 6464
rect 30324 6456 30350 6459
rect 30324 6427 30350 6430
rect 32946 6456 32972 6459
rect 32946 6427 32972 6430
rect 36356 6323 36370 6665
rect 36954 6629 36968 6835
rect 36948 6626 36974 6629
rect 36948 6597 36974 6600
rect 37362 6490 37388 6493
rect 37362 6461 37388 6464
rect 36350 6320 36376 6323
rect 36350 6291 36376 6294
rect 29312 5946 29338 5949
rect 29312 5917 29338 5920
rect 28852 5674 28878 5677
rect 28852 5645 28878 5648
rect 37368 5575 37382 6461
rect 37408 6422 37434 6425
rect 37408 6393 37434 6396
rect 37414 6153 37428 6393
rect 37500 6320 37526 6323
rect 37500 6291 37526 6294
rect 37408 6150 37434 6153
rect 37408 6121 37434 6124
rect 37506 5847 37520 6291
rect 37552 6221 37566 7600
rect 37684 6898 37710 6901
rect 37684 6869 37710 6872
rect 38006 6898 38032 6901
rect 38006 6869 38032 6872
rect 37690 6731 37704 6869
rect 37684 6728 37710 6731
rect 37684 6699 37710 6702
rect 37822 6728 37848 6731
rect 37822 6699 37848 6702
rect 37592 6626 37618 6629
rect 37592 6597 37618 6600
rect 37598 6323 37612 6597
rect 37730 6422 37756 6425
rect 37730 6393 37756 6396
rect 37592 6320 37618 6323
rect 37592 6291 37618 6294
rect 37546 6218 37572 6221
rect 37546 6189 37572 6192
rect 37736 5949 37750 6393
rect 37828 5949 37842 6699
rect 38012 6187 38026 6869
rect 38190 6864 38216 6867
rect 38190 6835 38216 6838
rect 38006 6184 38032 6187
rect 38006 6155 38032 6158
rect 37730 5946 37756 5949
rect 37730 5917 37756 5920
rect 37822 5946 37848 5949
rect 37822 5917 37848 5920
rect 38012 5881 38026 6155
rect 38144 6048 38170 6051
rect 38144 6019 38170 6022
rect 38150 5881 38164 6019
rect 38006 5878 38032 5881
rect 38006 5849 38032 5852
rect 38144 5878 38170 5881
rect 38144 5849 38170 5852
rect 37500 5844 37526 5847
rect 37500 5815 37526 5818
rect 38196 5677 38210 6835
rect 39202 6660 39228 6663
rect 39202 6631 39228 6634
rect 38236 6626 38262 6629
rect 38236 6597 38262 6600
rect 38242 5949 38256 6597
rect 38972 6592 38998 6595
rect 38972 6563 38998 6566
rect 38574 6542 38728 6546
rect 38574 6541 38577 6542
rect 38605 6541 38617 6542
rect 38645 6541 38657 6542
rect 38685 6541 38697 6542
rect 38725 6541 38728 6542
rect 38605 6515 38606 6541
rect 38696 6515 38697 6541
rect 38574 6514 38577 6515
rect 38605 6514 38617 6515
rect 38645 6514 38657 6515
rect 38685 6514 38697 6515
rect 38725 6514 38728 6515
rect 38574 6509 38728 6514
rect 38926 6354 38952 6357
rect 38926 6325 38952 6328
rect 38604 6320 38630 6323
rect 38604 6291 38630 6294
rect 38610 6187 38624 6291
rect 38604 6184 38630 6187
rect 38604 6155 38630 6158
rect 38466 6150 38492 6153
rect 38466 6121 38492 6124
rect 38236 5946 38262 5949
rect 38236 5917 38262 5920
rect 38472 5847 38486 6121
rect 38574 5998 38728 6002
rect 38574 5997 38577 5998
rect 38605 5997 38617 5998
rect 38645 5997 38657 5998
rect 38685 5997 38697 5998
rect 38725 5997 38728 5998
rect 38605 5971 38606 5997
rect 38696 5971 38697 5997
rect 38574 5970 38577 5971
rect 38605 5970 38617 5971
rect 38645 5970 38657 5971
rect 38685 5970 38697 5971
rect 38725 5970 38728 5971
rect 38574 5965 38728 5970
rect 38932 5949 38946 6325
rect 38978 6119 38992 6563
rect 39208 6459 39222 6631
rect 39202 6456 39228 6459
rect 39202 6427 39228 6430
rect 39064 6354 39090 6357
rect 39064 6325 39090 6328
rect 39070 6153 39084 6325
rect 39202 6184 39228 6187
rect 39202 6155 39228 6158
rect 39064 6150 39090 6153
rect 39064 6121 39090 6124
rect 38972 6116 38998 6119
rect 38972 6087 38998 6090
rect 38926 5946 38952 5949
rect 38926 5917 38952 5920
rect 38466 5844 38492 5847
rect 38466 5815 38492 5818
rect 38190 5674 38216 5677
rect 38190 5645 38216 5648
rect 39208 5575 39222 6155
rect 39254 5949 39268 7643
rect 40627 7643 40694 7657
rect 40627 7600 40655 7643
rect 40680 6705 40694 7643
rect 42145 7600 42173 8000
rect 43709 7600 43737 8000
rect 45227 7600 45255 8000
rect 46791 7657 46819 8000
rect 48309 7657 48337 8000
rect 46791 7643 46904 7657
rect 46791 7600 46819 7643
rect 41548 6864 41574 6867
rect 41548 6835 41574 6838
rect 40122 6694 40148 6697
rect 40680 6691 40740 6705
rect 40122 6665 40148 6668
rect 39990 6629 40050 6637
rect 39386 6626 39412 6629
rect 39386 6597 39412 6600
rect 39662 6626 39688 6629
rect 39662 6597 39688 6600
rect 39990 6626 40056 6629
rect 39990 6623 40030 6626
rect 39294 6388 39320 6391
rect 39294 6359 39320 6362
rect 39300 6119 39314 6359
rect 39294 6116 39320 6119
rect 39294 6087 39320 6090
rect 39248 5946 39274 5949
rect 39248 5917 39274 5920
rect 39300 5881 39314 6087
rect 39294 5878 39320 5881
rect 39294 5849 39320 5852
rect 39392 5677 39406 6597
rect 39668 6221 39682 6597
rect 39990 6433 40004 6623
rect 40030 6597 40056 6600
rect 39852 6425 40004 6433
rect 39846 6422 40004 6425
rect 39872 6419 40004 6422
rect 39846 6393 39872 6396
rect 39662 6218 39688 6221
rect 39662 6189 39688 6192
rect 40128 6051 40142 6665
rect 40726 6663 40740 6691
rect 40812 6694 40838 6697
rect 40812 6665 40838 6668
rect 40720 6660 40746 6663
rect 40720 6631 40746 6634
rect 40398 6592 40424 6595
rect 40398 6563 40424 6566
rect 40720 6592 40746 6595
rect 40720 6563 40746 6566
rect 40260 6456 40286 6459
rect 40260 6427 40286 6430
rect 40266 6221 40280 6427
rect 40404 6391 40418 6563
rect 40398 6388 40424 6391
rect 40398 6359 40424 6362
rect 40726 6357 40740 6563
rect 40720 6354 40746 6357
rect 40720 6325 40746 6328
rect 40260 6218 40286 6221
rect 40260 6189 40286 6192
rect 40726 6153 40740 6325
rect 40818 6323 40832 6665
rect 41554 6663 41568 6835
rect 41548 6660 41574 6663
rect 41548 6631 41574 6634
rect 41962 6660 41988 6663
rect 41962 6631 41988 6634
rect 41916 6626 41942 6629
rect 41916 6597 41942 6600
rect 41456 6592 41482 6595
rect 41456 6563 41482 6566
rect 41462 6459 41476 6563
rect 41456 6456 41482 6459
rect 41456 6427 41482 6430
rect 40812 6320 40838 6323
rect 40812 6291 40838 6294
rect 40720 6150 40746 6153
rect 40720 6121 40746 6124
rect 40122 6048 40148 6051
rect 40122 6019 40148 6022
rect 40726 5881 40740 6121
rect 40720 5878 40746 5881
rect 40720 5849 40746 5852
rect 39386 5674 39412 5677
rect 39386 5645 39412 5648
rect 17352 5572 17378 5575
rect 17352 5543 17378 5546
rect 20250 5572 20276 5575
rect 20250 5543 20276 5546
rect 20710 5572 20736 5575
rect 20710 5543 20736 5546
rect 21216 5572 21242 5575
rect 21216 5543 21242 5546
rect 27748 5572 27774 5575
rect 27748 5543 27774 5546
rect 28622 5572 28648 5575
rect 28622 5543 28648 5546
rect 37362 5572 37388 5575
rect 37362 5543 37388 5546
rect 39202 5572 39228 5575
rect 39202 5543 39228 5546
rect 40818 5541 40832 6291
rect 41922 6119 41936 6597
rect 41968 6595 41982 6631
rect 41962 6592 41988 6595
rect 41962 6563 41988 6566
rect 41968 6493 41982 6563
rect 41962 6490 41988 6493
rect 41962 6461 41988 6464
rect 41916 6116 41942 6119
rect 41916 6087 41942 6090
rect 42008 6048 42034 6051
rect 42008 6019 42034 6022
rect 42014 5847 42028 6019
rect 42152 5949 42166 7600
rect 43204 6864 43230 6867
rect 43204 6835 43230 6838
rect 42238 6626 42264 6629
rect 42238 6597 42264 6600
rect 42744 6626 42770 6629
rect 42744 6597 42770 6600
rect 42146 5946 42172 5949
rect 42146 5917 42172 5920
rect 42008 5844 42034 5847
rect 42008 5815 42034 5818
rect 42244 5677 42258 6597
rect 42422 6388 42448 6391
rect 42422 6359 42448 6362
rect 42330 6150 42356 6153
rect 42330 6121 42356 6124
rect 42336 6051 42350 6121
rect 42330 6048 42356 6051
rect 42330 6019 42356 6022
rect 42428 5779 42442 6359
rect 42750 6221 42764 6597
rect 43020 6592 43046 6595
rect 43020 6563 43046 6566
rect 42882 6320 42908 6323
rect 42882 6291 42908 6294
rect 42744 6218 42770 6221
rect 42744 6189 42770 6192
rect 42888 6153 42902 6291
rect 42882 6150 42908 6153
rect 42882 6121 42908 6124
rect 42744 6116 42770 6119
rect 42744 6087 42770 6090
rect 42468 5912 42494 5915
rect 42652 5912 42678 5915
rect 42494 5886 42652 5889
rect 42468 5883 42678 5886
rect 42474 5875 42672 5883
rect 42422 5776 42448 5779
rect 42422 5747 42448 5750
rect 42238 5674 42264 5677
rect 42238 5645 42264 5648
rect 42750 5609 42764 6087
rect 42888 5881 42902 6121
rect 43026 6119 43040 6563
rect 43210 6221 43224 6835
rect 43388 6626 43414 6629
rect 43388 6597 43414 6600
rect 43250 6490 43276 6493
rect 43250 6461 43276 6464
rect 43256 6391 43270 6461
rect 43250 6388 43276 6391
rect 43250 6359 43276 6362
rect 43204 6218 43230 6221
rect 43204 6189 43230 6192
rect 43066 6184 43092 6187
rect 43066 6155 43092 6158
rect 43020 6116 43046 6119
rect 43020 6087 43046 6090
rect 43026 5949 43040 6087
rect 43072 5949 43086 6155
rect 43158 6150 43184 6153
rect 43158 6121 43184 6124
rect 43164 6051 43178 6121
rect 43158 6048 43184 6051
rect 43158 6019 43184 6022
rect 43020 5946 43046 5949
rect 43020 5917 43046 5920
rect 43066 5946 43092 5949
rect 43066 5917 43092 5920
rect 42882 5878 42908 5881
rect 42882 5849 42908 5852
rect 43164 5847 43178 6019
rect 43158 5844 43184 5847
rect 43158 5815 43184 5818
rect 43204 5776 43230 5779
rect 43204 5747 43230 5750
rect 42744 5606 42770 5609
rect 42744 5577 42770 5580
rect 43210 5575 43224 5747
rect 43394 5643 43408 6597
rect 43479 6576 43507 6580
rect 43479 6543 43507 6548
rect 43486 5881 43500 6543
rect 43572 6490 43598 6493
rect 43572 6461 43598 6464
rect 43480 5878 43506 5881
rect 43480 5849 43506 5852
rect 43578 5677 43592 6461
rect 43716 6187 43730 7600
rect 43940 6660 43966 6663
rect 43940 6631 43966 6634
rect 43893 6372 43921 6376
rect 43893 6339 43921 6344
rect 43900 6323 43914 6339
rect 43894 6320 43920 6323
rect 43894 6291 43920 6294
rect 43946 6221 43960 6631
rect 44538 6626 44564 6629
rect 44538 6597 44564 6600
rect 44768 6626 44794 6629
rect 44768 6597 44794 6600
rect 44124 6592 44150 6595
rect 44124 6563 44150 6566
rect 44130 6391 44144 6563
rect 44124 6388 44150 6391
rect 44124 6359 44150 6362
rect 43986 6320 44012 6323
rect 43986 6291 44012 6294
rect 43940 6218 43966 6221
rect 43940 6189 43966 6192
rect 43710 6184 43736 6187
rect 43710 6155 43736 6158
rect 43992 6093 44006 6291
rect 44077 6168 44105 6172
rect 44077 6135 44078 6140
rect 44104 6135 44105 6140
rect 44078 6121 44104 6124
rect 44130 6119 44144 6359
rect 44216 6320 44242 6323
rect 44216 6291 44242 6294
rect 43762 6079 44006 6093
rect 44124 6116 44150 6119
rect 44124 6087 44150 6090
rect 43762 6051 43776 6079
rect 43992 6051 44006 6079
rect 43756 6048 43782 6051
rect 43756 6019 43782 6022
rect 43894 6048 43920 6051
rect 43894 6019 43920 6022
rect 43986 6048 44012 6051
rect 43986 6019 44012 6022
rect 43572 5674 43598 5677
rect 43572 5645 43598 5648
rect 43388 5640 43414 5643
rect 43388 5611 43414 5614
rect 43900 5575 43914 6019
rect 43940 5946 43966 5949
rect 43940 5917 43966 5920
rect 43204 5572 43230 5575
rect 43204 5543 43230 5546
rect 43894 5572 43920 5575
rect 43894 5543 43920 5546
rect 43946 5541 43960 5917
rect 44222 5575 44236 6291
rect 44492 6116 44518 6119
rect 44360 6090 44492 6093
rect 44360 6087 44518 6090
rect 44360 6079 44512 6087
rect 44360 6051 44374 6079
rect 44354 6048 44380 6051
rect 44354 6019 44380 6022
rect 44544 5677 44558 6597
rect 44584 6150 44610 6153
rect 44584 6121 44610 6124
rect 44590 5881 44604 6121
rect 44774 5949 44788 6597
rect 45234 6493 45248 7600
rect 45320 6898 45346 6901
rect 45320 6869 45346 6872
rect 45274 6592 45300 6595
rect 45274 6563 45300 6566
rect 45228 6490 45254 6493
rect 45228 6461 45254 6464
rect 45280 6459 45294 6563
rect 45274 6456 45300 6459
rect 45274 6427 45300 6430
rect 45326 6425 45340 6869
rect 45918 6864 45944 6867
rect 45918 6835 45944 6838
rect 45924 6629 45938 6835
rect 46890 6773 46904 7643
rect 48309 7643 48376 7657
rect 48309 7600 48337 7643
rect 46890 6759 46950 6773
rect 46936 6731 46950 6759
rect 46930 6728 46956 6731
rect 46930 6699 46956 6702
rect 45826 6626 45852 6629
rect 45826 6597 45852 6600
rect 45918 6626 45944 6629
rect 45918 6597 45944 6600
rect 46010 6626 46036 6629
rect 46010 6597 46036 6600
rect 45832 6493 45846 6597
rect 45924 6580 45938 6597
rect 45917 6576 45945 6580
rect 45917 6543 45945 6548
rect 45826 6490 45852 6493
rect 45826 6461 45852 6464
rect 45366 6456 45392 6459
rect 45366 6427 45392 6430
rect 45090 6422 45116 6425
rect 45090 6393 45116 6396
rect 45228 6422 45254 6425
rect 45228 6393 45254 6396
rect 45320 6422 45346 6425
rect 45320 6393 45346 6396
rect 44860 6388 44886 6391
rect 45044 6388 45070 6391
rect 44886 6368 45044 6382
rect 44860 6359 44886 6362
rect 45044 6359 45070 6362
rect 44952 6320 44978 6323
rect 44952 6291 44978 6294
rect 44958 6172 44972 6291
rect 45096 6221 45110 6393
rect 45090 6218 45116 6221
rect 45090 6189 45116 6192
rect 44951 6168 44979 6172
rect 44951 6135 44979 6140
rect 44768 5946 44794 5949
rect 44768 5917 44794 5920
rect 44584 5878 44610 5881
rect 44584 5849 44610 5852
rect 44538 5674 44564 5677
rect 44538 5645 44564 5648
rect 44590 5609 44604 5849
rect 45234 5847 45248 6393
rect 45372 6376 45386 6427
rect 45365 6372 45393 6376
rect 45365 6339 45393 6344
rect 46016 6119 46030 6597
rect 48362 6595 48376 7643
rect 49827 7600 49855 8000
rect 51391 7657 51419 8000
rect 52909 7657 52937 8000
rect 54427 7657 54455 8000
rect 55991 7657 56019 8000
rect 51391 7643 51458 7657
rect 51391 7600 51419 7643
rect 49834 6705 49848 7600
rect 51208 6898 51234 6901
rect 51208 6869 51234 6872
rect 50978 6864 51004 6867
rect 50978 6835 51004 6838
rect 49552 6694 49578 6697
rect 49552 6665 49578 6668
rect 49696 6691 49848 6705
rect 50380 6728 50406 6731
rect 50380 6699 50406 6702
rect 49000 6626 49026 6629
rect 49000 6597 49026 6600
rect 48356 6592 48382 6595
rect 48356 6563 48382 6566
rect 48770 6592 48796 6595
rect 48770 6563 48796 6566
rect 48776 6119 48790 6563
rect 49006 6493 49020 6597
rect 49000 6490 49026 6493
rect 49000 6461 49026 6464
rect 49558 6153 49572 6665
rect 49598 6626 49624 6629
rect 49598 6597 49624 6600
rect 49604 6391 49618 6597
rect 49598 6388 49624 6391
rect 49598 6359 49624 6362
rect 49598 6320 49624 6323
rect 49696 6314 49710 6691
rect 49828 6626 49854 6629
rect 49828 6597 49854 6600
rect 49736 6456 49762 6459
rect 49736 6427 49762 6430
rect 49624 6300 49710 6314
rect 49598 6291 49624 6294
rect 49742 6221 49756 6427
rect 49736 6218 49762 6221
rect 49736 6189 49762 6192
rect 49552 6150 49578 6153
rect 49552 6121 49578 6124
rect 46010 6116 46036 6119
rect 46010 6087 46036 6090
rect 48770 6116 48796 6119
rect 48770 6087 48796 6090
rect 49834 5949 49848 6597
rect 49966 6456 49992 6459
rect 49966 6427 49992 6430
rect 49972 6221 49986 6427
rect 50386 6323 50400 6699
rect 50702 6660 50728 6663
rect 50702 6631 50728 6634
rect 50472 6626 50498 6629
rect 50472 6597 50498 6600
rect 50380 6320 50406 6323
rect 50380 6291 50406 6294
rect 49966 6218 49992 6221
rect 49966 6189 49992 6192
rect 50386 6085 50400 6291
rect 50380 6082 50406 6085
rect 50380 6053 50406 6056
rect 50196 6048 50222 6051
rect 50196 6019 50222 6022
rect 49828 5946 49854 5949
rect 49828 5917 49854 5920
rect 50202 5881 50216 6019
rect 50196 5878 50222 5881
rect 50196 5849 50222 5852
rect 50386 5847 50400 6053
rect 50478 5949 50492 6597
rect 50518 6592 50544 6595
rect 50518 6563 50544 6566
rect 50524 6357 50538 6563
rect 50708 6391 50722 6631
rect 50702 6388 50728 6391
rect 50702 6359 50728 6362
rect 50840 6388 50866 6391
rect 50840 6359 50866 6362
rect 50518 6354 50544 6357
rect 50518 6325 50544 6328
rect 50524 6085 50538 6325
rect 50518 6082 50544 6085
rect 50518 6053 50544 6056
rect 50472 5946 50498 5949
rect 50472 5917 50498 5920
rect 45228 5844 45254 5847
rect 45228 5815 45254 5818
rect 50380 5844 50406 5847
rect 50380 5815 50406 5818
rect 44584 5606 44610 5609
rect 44584 5577 44610 5580
rect 44216 5572 44242 5575
rect 44216 5543 44242 5546
rect 40812 5538 40838 5541
rect 40812 5509 40838 5512
rect 43940 5538 43966 5541
rect 43940 5509 43966 5512
rect 38574 5454 38728 5458
rect 38574 5453 38577 5454
rect 38605 5453 38617 5454
rect 38645 5453 38657 5454
rect 38685 5453 38697 5454
rect 38725 5453 38728 5454
rect 38605 5427 38606 5453
rect 38696 5427 38697 5453
rect 38574 5426 38577 5427
rect 38605 5426 38617 5427
rect 38645 5426 38657 5427
rect 38685 5426 38697 5427
rect 38725 5426 38728 5427
rect 38574 5421 38728 5426
rect 50846 5405 50860 6359
rect 50984 6085 50998 6835
rect 51116 6626 51142 6629
rect 51116 6597 51142 6600
rect 51024 6150 51050 6153
rect 51024 6121 51050 6124
rect 50978 6082 51004 6085
rect 50978 6053 51004 6056
rect 51030 5847 51044 6121
rect 51070 6082 51096 6085
rect 51070 6053 51096 6056
rect 51076 5881 51090 6053
rect 51070 5878 51096 5881
rect 51070 5849 51096 5852
rect 51024 5844 51050 5847
rect 51024 5815 51050 5818
rect 50932 5776 50958 5779
rect 50932 5747 50958 5750
rect 50840 5402 50866 5405
rect 50840 5373 50866 5376
rect 50938 5337 50952 5747
rect 51030 5609 51044 5815
rect 51122 5643 51136 6597
rect 51162 6048 51188 6051
rect 51162 6019 51188 6022
rect 51168 5847 51182 6019
rect 51162 5844 51188 5847
rect 51162 5815 51188 5818
rect 51116 5640 51142 5643
rect 51116 5611 51142 5614
rect 51024 5606 51050 5609
rect 51024 5577 51050 5580
rect 51214 5575 51228 6869
rect 51300 6048 51326 6051
rect 51300 6019 51326 6022
rect 51306 5609 51320 6019
rect 51444 5677 51458 7643
rect 52909 7643 52976 7657
rect 52909 7600 52937 7643
rect 51668 6660 51694 6663
rect 51668 6631 51694 6634
rect 52128 6660 52154 6663
rect 52128 6631 52154 6634
rect 51622 6354 51648 6357
rect 51622 6325 51648 6328
rect 51530 6320 51556 6323
rect 51530 6291 51556 6294
rect 51536 6051 51550 6291
rect 51628 6153 51642 6325
rect 51674 6153 51688 6631
rect 52036 6626 52062 6629
rect 52036 6597 52062 6600
rect 51852 6592 51878 6595
rect 51852 6563 51878 6566
rect 51806 6320 51832 6323
rect 51806 6291 51832 6294
rect 51622 6150 51648 6153
rect 51622 6121 51648 6124
rect 51668 6150 51694 6153
rect 51668 6121 51694 6124
rect 51530 6048 51556 6051
rect 51530 6019 51556 6022
rect 51536 5949 51550 6019
rect 51530 5946 51556 5949
rect 51530 5917 51556 5920
rect 51760 5946 51786 5949
rect 51760 5917 51786 5920
rect 51438 5674 51464 5677
rect 51438 5645 51464 5648
rect 51300 5606 51326 5609
rect 51300 5577 51326 5580
rect 51536 5575 51550 5917
rect 51766 5847 51780 5917
rect 51812 5881 51826 6291
rect 51858 6119 51872 6563
rect 51852 6116 51878 6119
rect 51852 6087 51878 6090
rect 51806 5878 51832 5881
rect 51806 5849 51832 5852
rect 51760 5844 51786 5847
rect 51760 5815 51786 5818
rect 52042 5779 52056 6597
rect 52036 5776 52062 5779
rect 52036 5747 52062 5750
rect 51208 5572 51234 5575
rect 51208 5543 51234 5546
rect 51530 5572 51556 5575
rect 51530 5543 51556 5546
rect 50932 5334 50958 5337
rect 50932 5305 50958 5308
rect 19524 5182 19678 5186
rect 19524 5181 19527 5182
rect 19555 5181 19567 5182
rect 19595 5181 19607 5182
rect 19635 5181 19647 5182
rect 19675 5181 19678 5182
rect 19555 5155 19556 5181
rect 19646 5155 19647 5181
rect 19524 5154 19527 5155
rect 19555 5154 19567 5155
rect 19595 5154 19607 5155
rect 19635 5154 19647 5155
rect 19675 5154 19678 5155
rect 19524 5149 19678 5154
rect 16708 5028 16734 5031
rect 16708 4999 16734 5002
rect 16846 5028 16872 5031
rect 16846 4999 16872 5002
rect 15604 4824 15630 4827
rect 15604 4795 15630 4798
rect 16852 4793 16866 4999
rect 38574 4910 38728 4914
rect 38574 4909 38577 4910
rect 38605 4909 38617 4910
rect 38645 4909 38657 4910
rect 38685 4909 38697 4910
rect 38725 4909 38728 4910
rect 38605 4883 38606 4909
rect 38696 4883 38697 4909
rect 38574 4882 38577 4883
rect 38605 4882 38617 4883
rect 38645 4882 38657 4883
rect 38685 4882 38697 4883
rect 38725 4882 38728 4883
rect 38574 4877 38728 4882
rect 16846 4790 16872 4793
rect 16846 4761 16872 4764
rect 15282 4756 15308 4759
rect 15282 4727 15308 4730
rect 14960 4722 14986 4725
rect 14960 4693 14986 4696
rect 52134 4691 52148 6631
rect 52226 6623 52378 6637
rect 52226 6595 52240 6623
rect 52220 6592 52246 6595
rect 52220 6563 52246 6566
rect 52312 6592 52338 6595
rect 52312 6563 52338 6566
rect 52318 6459 52332 6563
rect 52364 6459 52378 6623
rect 52496 6626 52522 6629
rect 52496 6597 52522 6600
rect 52312 6456 52338 6459
rect 52312 6427 52338 6430
rect 52358 6456 52384 6459
rect 52358 6427 52384 6430
rect 52502 6221 52516 6597
rect 52588 6422 52614 6425
rect 52588 6393 52614 6396
rect 52594 6221 52608 6393
rect 52962 6357 52976 7643
rect 54427 7643 54494 7657
rect 54427 7600 54455 7643
rect 54480 6773 54494 7643
rect 55906 7643 56019 7657
rect 55906 6773 55920 7643
rect 55991 7600 56019 7643
rect 57509 7600 57537 8000
rect 59073 7657 59101 8000
rect 60591 7657 60619 8000
rect 59073 7643 59324 7657
rect 59073 7600 59101 7643
rect 56912 6898 56938 6901
rect 56912 6869 56938 6872
rect 54480 6759 54540 6773
rect 54526 6731 54540 6759
rect 55860 6759 55920 6773
rect 55860 6731 55874 6759
rect 54520 6728 54546 6731
rect 54520 6699 54546 6702
rect 55854 6728 55880 6731
rect 55854 6699 55880 6702
rect 54796 6660 54822 6663
rect 54796 6631 54822 6634
rect 55716 6660 55742 6663
rect 55716 6631 55742 6634
rect 54802 6595 54816 6631
rect 54796 6592 54822 6595
rect 54796 6563 54822 6566
rect 54802 6459 54816 6563
rect 55722 6493 55736 6631
rect 56268 6626 56294 6629
rect 56268 6597 56294 6600
rect 55716 6490 55742 6493
rect 55716 6461 55742 6464
rect 54796 6456 54822 6459
rect 54796 6427 54822 6430
rect 52956 6354 52982 6357
rect 52956 6325 52982 6328
rect 55946 6320 55972 6323
rect 55946 6291 55972 6294
rect 52496 6218 52522 6221
rect 52496 6189 52522 6192
rect 52588 6218 52614 6221
rect 52588 6189 52614 6192
rect 55952 6119 55966 6291
rect 56274 6221 56288 6597
rect 56918 6425 56932 6869
rect 57326 6864 57352 6867
rect 57326 6835 57352 6838
rect 57096 6626 57122 6629
rect 57096 6597 57122 6600
rect 56544 6422 56570 6425
rect 56544 6393 56570 6396
rect 56912 6422 56938 6425
rect 56912 6393 56938 6396
rect 56550 6323 56564 6393
rect 56544 6320 56570 6323
rect 56544 6291 56570 6294
rect 56268 6218 56294 6221
rect 56268 6189 56294 6192
rect 56918 6161 56932 6393
rect 56958 6388 56984 6391
rect 56958 6359 56984 6362
rect 56872 6147 56932 6161
rect 55946 6116 55972 6119
rect 55946 6087 55972 6090
rect 56872 5541 56886 6147
rect 56912 6082 56938 6085
rect 56912 6053 56938 6056
rect 56918 5949 56932 6053
rect 56964 6051 56978 6359
rect 56958 6048 56984 6051
rect 56958 6019 56984 6022
rect 56912 5946 56938 5949
rect 56912 5917 56938 5920
rect 57004 5878 57030 5881
rect 57004 5849 57030 5852
rect 57010 5779 57024 5849
rect 57004 5776 57030 5779
rect 57004 5747 57030 5750
rect 57102 5643 57116 6597
rect 57280 6592 57306 6595
rect 57280 6563 57306 6566
rect 57286 6493 57300 6563
rect 57280 6490 57306 6493
rect 57280 6461 57306 6464
rect 57332 6425 57346 6835
rect 57418 6660 57444 6663
rect 57418 6631 57444 6634
rect 57372 6490 57398 6493
rect 57372 6461 57398 6464
rect 57326 6422 57352 6425
rect 57326 6393 57352 6396
rect 57332 6161 57346 6393
rect 57378 6391 57392 6461
rect 57372 6388 57398 6391
rect 57372 6359 57398 6362
rect 57424 6357 57438 6631
rect 57464 6592 57490 6595
rect 57464 6563 57490 6566
rect 57418 6354 57444 6357
rect 57418 6325 57444 6328
rect 57372 6320 57398 6323
rect 57372 6291 57398 6294
rect 57286 6147 57346 6161
rect 57142 6116 57168 6119
rect 57142 6087 57168 6090
rect 57148 5949 57162 6087
rect 57142 5946 57168 5949
rect 57142 5917 57168 5920
rect 57286 5915 57300 6147
rect 57280 5912 57306 5915
rect 57280 5883 57306 5886
rect 57096 5640 57122 5643
rect 57096 5611 57122 5614
rect 57378 5575 57392 6291
rect 57470 6161 57484 6563
rect 57516 6221 57530 7600
rect 59310 6841 59324 7643
rect 60591 7643 60658 7657
rect 60591 7600 60619 7643
rect 59310 6827 59370 6841
rect 57623 6814 57777 6818
rect 57623 6813 57626 6814
rect 57654 6813 57666 6814
rect 57694 6813 57706 6814
rect 57734 6813 57746 6814
rect 57774 6813 57777 6814
rect 57654 6787 57655 6813
rect 57745 6787 57746 6813
rect 57623 6786 57626 6787
rect 57654 6786 57666 6787
rect 57694 6786 57706 6787
rect 57734 6786 57746 6787
rect 57774 6786 57777 6787
rect 57623 6781 57777 6786
rect 59120 6694 59146 6697
rect 59120 6665 59146 6668
rect 58706 6660 58732 6663
rect 58706 6631 58732 6634
rect 57556 6626 57582 6629
rect 57556 6597 57582 6600
rect 58476 6626 58502 6629
rect 58476 6597 58502 6600
rect 57510 6218 57536 6221
rect 57510 6189 57536 6192
rect 57470 6147 57530 6161
rect 57516 5881 57530 6147
rect 57510 5878 57536 5881
rect 57510 5849 57536 5852
rect 57562 5677 57576 6597
rect 57878 6592 57904 6595
rect 57878 6563 57904 6566
rect 57884 6459 57898 6563
rect 57878 6456 57904 6459
rect 57878 6427 57904 6430
rect 57832 6388 57858 6391
rect 57924 6388 57950 6391
rect 57832 6359 57858 6362
rect 57884 6362 57924 6365
rect 57884 6359 57950 6362
rect 58384 6388 58410 6391
rect 58384 6359 58410 6362
rect 57623 6270 57777 6274
rect 57623 6269 57626 6270
rect 57654 6269 57666 6270
rect 57694 6269 57706 6270
rect 57734 6269 57746 6270
rect 57774 6269 57777 6270
rect 57654 6243 57655 6269
rect 57745 6243 57746 6269
rect 57623 6242 57626 6243
rect 57654 6242 57666 6243
rect 57694 6242 57706 6243
rect 57734 6242 57746 6243
rect 57774 6242 57777 6243
rect 57623 6237 57777 6242
rect 57838 6051 57852 6359
rect 57884 6351 57944 6359
rect 57884 6187 57898 6351
rect 57924 6320 57950 6323
rect 57924 6291 57950 6294
rect 57878 6184 57904 6187
rect 57878 6155 57904 6158
rect 57832 6048 57858 6051
rect 57832 6019 57858 6022
rect 57838 5949 57852 6019
rect 57832 5946 57858 5949
rect 57832 5917 57858 5920
rect 57884 5889 57898 6155
rect 57838 5875 57898 5889
rect 57838 5847 57852 5875
rect 57832 5844 57858 5847
rect 57832 5815 57858 5818
rect 57878 5844 57904 5847
rect 57878 5815 57904 5818
rect 57623 5726 57777 5730
rect 57623 5725 57626 5726
rect 57654 5725 57666 5726
rect 57694 5725 57706 5726
rect 57734 5725 57746 5726
rect 57774 5725 57777 5726
rect 57654 5699 57655 5725
rect 57745 5699 57746 5725
rect 57623 5698 57626 5699
rect 57654 5698 57666 5699
rect 57694 5698 57706 5699
rect 57734 5698 57746 5699
rect 57774 5698 57777 5699
rect 57623 5693 57777 5698
rect 57556 5674 57582 5677
rect 57556 5645 57582 5648
rect 57884 5575 57898 5815
rect 57930 5575 57944 6291
rect 58200 6048 58226 6051
rect 58200 6019 58226 6022
rect 58206 5881 58220 6019
rect 58390 5949 58404 6359
rect 58482 6221 58496 6597
rect 58712 6493 58726 6631
rect 58844 6626 58870 6629
rect 58844 6597 58870 6600
rect 58706 6490 58732 6493
rect 58706 6461 58732 6464
rect 58660 6456 58686 6459
rect 58660 6427 58686 6430
rect 58476 6218 58502 6221
rect 58476 6189 58502 6192
rect 58666 5949 58680 6427
rect 58384 5946 58410 5949
rect 58384 5917 58410 5920
rect 58660 5946 58686 5949
rect 58660 5917 58686 5920
rect 58200 5878 58226 5881
rect 58200 5849 58226 5852
rect 57372 5572 57398 5575
rect 57372 5543 57398 5546
rect 57878 5572 57904 5575
rect 57878 5543 57904 5546
rect 57924 5572 57950 5575
rect 57924 5543 57950 5546
rect 56866 5538 56892 5541
rect 56866 5509 56892 5512
rect 57623 5182 57777 5186
rect 57623 5181 57626 5182
rect 57654 5181 57666 5182
rect 57694 5181 57706 5182
rect 57734 5181 57746 5182
rect 57774 5181 57777 5182
rect 57654 5155 57655 5181
rect 57745 5155 57746 5181
rect 57623 5154 57626 5155
rect 57654 5154 57666 5155
rect 57694 5154 57706 5155
rect 57734 5154 57746 5155
rect 57774 5154 57777 5155
rect 57623 5149 57777 5154
rect 58712 4963 58726 6461
rect 58850 5677 58864 6597
rect 59028 6592 59054 6595
rect 59028 6563 59054 6566
rect 59034 6425 59048 6563
rect 59126 6493 59140 6665
rect 59356 6493 59370 6827
rect 60644 6731 60658 7643
rect 62109 7600 62137 8000
rect 63673 7657 63701 8000
rect 63496 7643 63701 7657
rect 62116 6841 62130 7600
rect 62754 6898 62780 6901
rect 62754 6869 62780 6872
rect 62070 6827 62130 6841
rect 62070 6731 62084 6827
rect 59442 6728 59468 6731
rect 59442 6699 59468 6702
rect 60638 6728 60664 6731
rect 60638 6699 60664 6702
rect 62064 6728 62090 6731
rect 62064 6699 62090 6702
rect 59396 6660 59422 6663
rect 59396 6631 59422 6634
rect 59120 6490 59146 6493
rect 59120 6461 59146 6464
rect 59350 6490 59376 6493
rect 59350 6461 59376 6464
rect 59028 6422 59054 6425
rect 59028 6393 59054 6396
rect 59034 6119 59048 6393
rect 59028 6116 59054 6119
rect 59028 6087 59054 6090
rect 59126 6085 59140 6461
rect 59166 6116 59192 6119
rect 59166 6087 59192 6090
rect 59120 6082 59146 6085
rect 59120 6053 59146 6056
rect 59172 5881 59186 6087
rect 59402 5949 59416 6631
rect 59448 6153 59462 6699
rect 62760 6629 62774 6869
rect 62754 6626 62780 6629
rect 62754 6597 62780 6600
rect 59856 6592 59882 6595
rect 59856 6563 59882 6566
rect 63076 6592 63102 6595
rect 63076 6563 63102 6566
rect 63260 6592 63286 6595
rect 63260 6563 63286 6566
rect 59442 6150 59468 6153
rect 59442 6121 59468 6124
rect 59396 5946 59422 5949
rect 59396 5917 59422 5920
rect 59166 5878 59192 5881
rect 59166 5849 59192 5852
rect 58844 5674 58870 5677
rect 58844 5645 58870 5648
rect 59862 5575 59876 6563
rect 63082 6119 63096 6563
rect 63266 6459 63280 6563
rect 63496 6501 63510 7643
rect 63673 7600 63701 7643
rect 65191 7600 65219 8000
rect 66709 7657 66737 8000
rect 66709 7643 66914 7657
rect 66709 7600 66737 7643
rect 63720 6864 63746 6867
rect 63720 6835 63746 6838
rect 63766 6864 63792 6867
rect 63766 6835 63792 6838
rect 64870 6864 64896 6867
rect 64870 6835 64896 6838
rect 63450 6493 63510 6501
rect 63444 6490 63510 6493
rect 63470 6487 63510 6490
rect 63444 6461 63470 6464
rect 63260 6456 63286 6459
rect 63260 6427 63286 6430
rect 63726 6425 63740 6835
rect 63772 6731 63786 6835
rect 63766 6728 63792 6731
rect 63766 6699 63792 6702
rect 63766 6660 63792 6663
rect 63766 6631 63792 6634
rect 64686 6660 64712 6663
rect 64686 6631 64712 6634
rect 63720 6422 63746 6425
rect 63720 6393 63746 6396
rect 63772 6391 63786 6631
rect 63904 6626 63930 6629
rect 63904 6597 63930 6600
rect 63766 6388 63792 6391
rect 63766 6359 63792 6362
rect 63910 6221 63924 6597
rect 64042 6592 64068 6595
rect 64042 6563 64068 6566
rect 64594 6592 64620 6595
rect 64594 6563 64620 6566
rect 64048 6493 64062 6563
rect 64600 6493 64614 6563
rect 64042 6490 64068 6493
rect 64042 6461 64068 6464
rect 64318 6490 64344 6493
rect 64318 6461 64344 6464
rect 64594 6490 64620 6493
rect 64594 6461 64620 6464
rect 64180 6388 64206 6391
rect 64180 6359 64206 6362
rect 64042 6320 64068 6323
rect 64186 6297 64200 6359
rect 64068 6294 64200 6297
rect 64042 6291 64200 6294
rect 64048 6283 64200 6291
rect 63904 6218 63930 6221
rect 63904 6189 63930 6192
rect 63076 6116 63102 6119
rect 63076 6087 63102 6090
rect 64186 5881 64200 6283
rect 64324 6119 64338 6461
rect 64548 6422 64574 6425
rect 64548 6393 64574 6396
rect 64554 6221 64568 6393
rect 64548 6218 64574 6221
rect 64548 6189 64574 6192
rect 64318 6116 64344 6119
rect 64318 6087 64344 6090
rect 64692 5949 64706 6631
rect 64876 6391 64890 6835
rect 65146 6694 65172 6697
rect 65146 6665 65172 6668
rect 65152 6425 65166 6665
rect 65146 6422 65172 6425
rect 65146 6393 65172 6396
rect 64870 6388 64896 6391
rect 64870 6359 64896 6362
rect 64686 5946 64712 5949
rect 64686 5917 64712 5920
rect 64180 5878 64206 5881
rect 64180 5849 64206 5852
rect 64876 5847 64890 6359
rect 65146 6354 65172 6357
rect 65146 6325 65172 6328
rect 65152 5949 65166 6325
rect 65146 5946 65172 5949
rect 65146 5917 65172 5920
rect 65146 5878 65172 5881
rect 65146 5849 65172 5852
rect 64870 5844 64896 5847
rect 64870 5815 64896 5818
rect 65152 5609 65166 5849
rect 65198 5677 65212 7600
rect 65928 6898 65954 6901
rect 65928 6869 65954 6872
rect 65606 6626 65632 6629
rect 65606 6597 65632 6600
rect 65560 6388 65586 6391
rect 65560 6359 65586 6362
rect 65468 6218 65494 6221
rect 65468 6189 65494 6192
rect 65238 6116 65264 6119
rect 65238 6087 65264 6090
rect 65192 5674 65218 5677
rect 65192 5645 65218 5648
rect 65146 5606 65172 5609
rect 65146 5577 65172 5580
rect 59856 5572 59882 5575
rect 59856 5543 59882 5546
rect 65152 5337 65166 5577
rect 65244 5405 65258 6087
rect 65474 5949 65488 6189
rect 65514 6150 65540 6153
rect 65514 6121 65540 6124
rect 65468 5946 65494 5949
rect 65468 5917 65494 5920
rect 65474 5575 65488 5917
rect 65520 5847 65534 6121
rect 65566 5949 65580 6359
rect 65560 5946 65586 5949
rect 65560 5917 65586 5920
rect 65514 5844 65540 5847
rect 65514 5815 65540 5818
rect 65612 5677 65626 6597
rect 65790 6592 65816 6595
rect 65790 6563 65816 6566
rect 65796 6051 65810 6563
rect 65790 6048 65816 6051
rect 65790 6019 65816 6022
rect 65796 5881 65810 6019
rect 65790 5878 65816 5881
rect 65790 5849 65816 5852
rect 65934 5779 65948 6869
rect 66802 6864 66828 6867
rect 66802 6835 66828 6838
rect 66434 6626 66460 6629
rect 66434 6597 66460 6600
rect 66664 6626 66690 6629
rect 66664 6597 66690 6600
rect 66204 6456 66230 6459
rect 66204 6427 66230 6430
rect 66210 6221 66224 6427
rect 66296 6388 66322 6391
rect 66296 6359 66322 6362
rect 66204 6218 66230 6221
rect 66204 6189 66230 6192
rect 66302 6161 66316 6359
rect 66210 6147 66316 6161
rect 66210 6119 66224 6147
rect 66204 6116 66230 6119
rect 66204 6087 66230 6090
rect 66296 6116 66322 6119
rect 66296 6087 66322 6090
rect 66250 6082 66276 6085
rect 66250 6053 66276 6056
rect 66256 5881 66270 6053
rect 66250 5878 66276 5881
rect 66250 5849 66276 5852
rect 65928 5776 65954 5779
rect 65928 5747 65954 5750
rect 65606 5674 65632 5677
rect 65606 5645 65632 5648
rect 66302 5609 66316 6087
rect 66440 5677 66454 6597
rect 66670 6493 66684 6597
rect 66664 6490 66690 6493
rect 66664 6461 66690 6464
rect 66808 6459 66822 6835
rect 66900 6637 66914 7643
rect 68273 7600 68301 8000
rect 69791 7600 69819 8000
rect 71355 7657 71383 8000
rect 71355 7643 71468 7657
rect 71355 7600 71383 7643
rect 68280 6841 68294 7600
rect 68412 6864 68438 6867
rect 68280 6827 68340 6841
rect 68412 6835 68438 6838
rect 68326 6731 68340 6827
rect 68320 6728 68346 6731
rect 68320 6699 68346 6702
rect 68418 6663 68432 6835
rect 69798 6731 69812 7600
rect 71454 6765 71468 7643
rect 72873 7600 72901 8000
rect 74391 7657 74419 8000
rect 74260 7643 74419 7657
rect 72880 6765 72894 7600
rect 74070 6864 74096 6867
rect 74070 6835 74096 6838
rect 74076 6765 74090 6835
rect 71448 6762 71474 6765
rect 71448 6733 71474 6736
rect 72874 6762 72900 6765
rect 72874 6733 72900 6736
rect 74070 6762 74096 6765
rect 74070 6733 74096 6736
rect 69792 6728 69818 6731
rect 69792 6699 69818 6702
rect 71034 6694 71060 6697
rect 71034 6665 71060 6668
rect 68412 6660 68438 6663
rect 66900 6623 66960 6637
rect 68412 6631 68438 6634
rect 66848 6592 66874 6595
rect 66848 6563 66874 6566
rect 66802 6456 66828 6459
rect 66802 6427 66828 6430
rect 66854 6425 66868 6563
rect 66946 6493 66960 6623
rect 67078 6592 67104 6595
rect 67078 6563 67104 6566
rect 66940 6490 66966 6493
rect 66940 6461 66966 6464
rect 67084 6459 67098 6563
rect 67078 6456 67104 6459
rect 67078 6427 67104 6430
rect 66848 6422 66874 6425
rect 66848 6393 66874 6396
rect 66854 6357 66960 6365
rect 66848 6354 66966 6357
rect 66874 6351 66940 6354
rect 66848 6325 66874 6328
rect 66940 6325 66966 6328
rect 66572 6320 66598 6323
rect 66572 6291 66598 6294
rect 66618 6320 66644 6323
rect 66618 6291 66644 6294
rect 66434 5674 66460 5677
rect 66434 5645 66460 5648
rect 66296 5606 66322 5609
rect 66296 5577 66322 5580
rect 66578 5575 66592 6291
rect 66624 6153 66638 6291
rect 70988 6184 71014 6187
rect 70988 6155 71014 6158
rect 66618 6150 66644 6153
rect 66618 6121 66644 6124
rect 68872 6116 68898 6119
rect 68872 6087 68898 6090
rect 68878 5949 68892 6087
rect 69010 6082 69036 6085
rect 69010 6053 69036 6056
rect 68872 5946 68898 5949
rect 68872 5917 68898 5920
rect 68878 5847 68892 5917
rect 69016 5915 69030 6053
rect 69010 5912 69036 5915
rect 69010 5883 69036 5886
rect 68872 5844 68898 5847
rect 68872 5815 68898 5818
rect 65468 5572 65494 5575
rect 65468 5543 65494 5546
rect 66572 5572 66598 5575
rect 66572 5543 66598 5546
rect 70344 5538 70370 5541
rect 70344 5509 70370 5512
rect 65238 5402 65264 5405
rect 65238 5373 65264 5376
rect 70350 5371 70364 5509
rect 70994 5405 71008 6155
rect 71040 5575 71054 6665
rect 71540 6660 71566 6663
rect 71540 6631 71566 6634
rect 72874 6660 72900 6663
rect 72874 6631 72900 6634
rect 71546 6459 71560 6631
rect 71540 6456 71566 6459
rect 71540 6427 71566 6430
rect 71632 6388 71658 6391
rect 71632 6359 71658 6362
rect 71638 5813 71652 6359
rect 72880 6357 72894 6631
rect 72966 6626 72992 6629
rect 72966 6597 72992 6600
rect 73012 6626 73038 6629
rect 73012 6597 73038 6600
rect 73794 6626 73820 6629
rect 73794 6597 73820 6600
rect 72920 6592 72946 6595
rect 72920 6563 72946 6566
rect 72926 6425 72940 6563
rect 72972 6459 72986 6597
rect 72966 6456 72992 6459
rect 72966 6427 72992 6430
rect 72920 6422 72946 6425
rect 72920 6393 72946 6396
rect 72874 6354 72900 6357
rect 72874 6325 72900 6328
rect 71632 5810 71658 5813
rect 71632 5781 71658 5784
rect 71638 5609 71652 5781
rect 71632 5606 71658 5609
rect 71632 5577 71658 5580
rect 72880 5575 72894 6325
rect 73018 5813 73032 6597
rect 73748 6592 73774 6595
rect 73748 6563 73774 6566
rect 73656 6422 73682 6425
rect 73656 6393 73682 6396
rect 73012 5810 73038 5813
rect 73012 5781 73038 5784
rect 73662 5779 73676 6393
rect 73702 6388 73728 6391
rect 73702 6359 73728 6362
rect 73656 5776 73682 5779
rect 73656 5747 73682 5750
rect 73708 5643 73722 6359
rect 73702 5640 73728 5643
rect 73702 5611 73728 5614
rect 73754 5609 73768 6563
rect 73800 6187 73814 6597
rect 73840 6490 73866 6493
rect 73840 6461 73866 6464
rect 73794 6184 73820 6187
rect 73794 6155 73820 6158
rect 73846 5881 73860 6461
rect 73886 6388 73912 6391
rect 73886 6359 73912 6362
rect 73892 6221 73906 6359
rect 74260 6323 74274 7643
rect 74391 7600 74419 7643
rect 75955 7657 75983 8000
rect 75955 7643 76022 7657
rect 75955 7600 75983 7643
rect 75220 6864 75246 6867
rect 75220 6835 75246 6838
rect 75226 6629 75240 6835
rect 75404 6762 75430 6765
rect 75404 6733 75430 6736
rect 75220 6626 75246 6629
rect 75220 6597 75246 6600
rect 74622 6592 74648 6595
rect 74622 6563 74648 6566
rect 74628 6391 74642 6563
rect 75226 6425 75240 6597
rect 74668 6422 74694 6425
rect 74668 6393 74694 6396
rect 75220 6422 75246 6425
rect 75220 6393 75246 6396
rect 74484 6388 74510 6391
rect 74622 6388 74648 6391
rect 74484 6359 74510 6362
rect 74536 6368 74622 6382
rect 74254 6320 74280 6323
rect 74254 6291 74280 6294
rect 73886 6218 73912 6221
rect 73886 6189 73912 6192
rect 74024 6116 74050 6119
rect 74024 6087 74050 6090
rect 73840 5878 73866 5881
rect 73840 5849 73866 5852
rect 74030 5677 74044 6087
rect 74162 5844 74188 5847
rect 74162 5815 74188 5818
rect 74300 5844 74326 5847
rect 74300 5815 74326 5818
rect 74024 5674 74050 5677
rect 74024 5645 74050 5648
rect 73748 5606 73774 5609
rect 73748 5577 73774 5580
rect 71034 5572 71060 5575
rect 71034 5543 71060 5546
rect 72874 5572 72900 5575
rect 72874 5543 72900 5546
rect 70988 5402 71014 5405
rect 70988 5373 71014 5376
rect 70344 5368 70370 5371
rect 70344 5339 70370 5342
rect 65146 5334 65172 5337
rect 65146 5305 65172 5308
rect 70350 5031 70364 5339
rect 70344 5028 70370 5031
rect 70344 4999 70370 5002
rect 58706 4960 58732 4963
rect 58706 4931 58732 4934
rect 70350 4827 70364 4999
rect 70344 4824 70370 4827
rect 70344 4795 70370 4798
rect 74168 4691 74182 5815
rect 74306 5405 74320 5815
rect 74490 5405 74504 6359
rect 74536 6153 74550 6368
rect 74622 6359 74648 6362
rect 74530 6150 74556 6153
rect 74530 6121 74556 6124
rect 74536 5507 74550 6121
rect 74674 6119 74688 6393
rect 75174 6354 75200 6357
rect 75174 6325 75200 6328
rect 74990 6320 75016 6323
rect 74990 6291 75016 6294
rect 74668 6116 74694 6119
rect 74668 6087 74694 6090
rect 74714 6116 74740 6119
rect 74714 6087 74740 6090
rect 74530 5504 74556 5507
rect 74530 5475 74556 5478
rect 74300 5402 74326 5405
rect 74300 5373 74326 5376
rect 74484 5402 74510 5405
rect 74484 5373 74510 5376
rect 52128 4688 52154 4691
rect 52128 4659 52154 4662
rect 74162 4688 74188 4691
rect 74162 4659 74188 4662
rect 19524 4638 19678 4642
rect 19524 4637 19527 4638
rect 19555 4637 19567 4638
rect 19595 4637 19607 4638
rect 19635 4637 19647 4638
rect 19675 4637 19678 4638
rect 19555 4611 19556 4637
rect 19646 4611 19647 4637
rect 19524 4610 19527 4611
rect 19555 4610 19567 4611
rect 19595 4610 19607 4611
rect 19635 4610 19647 4611
rect 19675 4610 19678 4611
rect 19524 4605 19678 4610
rect 57623 4638 57777 4642
rect 57623 4637 57626 4638
rect 57654 4637 57666 4638
rect 57694 4637 57706 4638
rect 57734 4637 57746 4638
rect 57774 4637 57777 4638
rect 57654 4611 57655 4637
rect 57745 4611 57746 4637
rect 57623 4610 57626 4611
rect 57654 4610 57666 4611
rect 57694 4610 57706 4611
rect 57734 4610 57746 4611
rect 57774 4610 57777 4611
rect 57623 4605 57777 4610
rect 38574 4366 38728 4370
rect 38574 4365 38577 4366
rect 38605 4365 38617 4366
rect 38645 4365 38657 4366
rect 38685 4365 38697 4366
rect 38725 4365 38728 4366
rect 38605 4339 38606 4365
rect 38696 4339 38697 4365
rect 38574 4338 38577 4339
rect 38605 4338 38617 4339
rect 38645 4338 38657 4339
rect 38685 4338 38697 4339
rect 38725 4338 38728 4339
rect 38574 4333 38728 4338
rect 700 4178 726 4181
rect 700 4149 726 4152
rect 706 4064 720 4149
rect 19524 4094 19678 4098
rect 19524 4093 19527 4094
rect 19555 4093 19567 4094
rect 19595 4093 19607 4094
rect 19635 4093 19647 4094
rect 19675 4093 19678 4094
rect 19555 4067 19556 4093
rect 19646 4067 19647 4093
rect 19524 4066 19527 4067
rect 19555 4066 19567 4067
rect 19595 4066 19607 4067
rect 19635 4066 19647 4067
rect 19675 4066 19678 4067
rect 699 4060 727 4064
rect 19524 4061 19678 4066
rect 57623 4094 57777 4098
rect 57623 4093 57626 4094
rect 57654 4093 57666 4094
rect 57694 4093 57706 4094
rect 57734 4093 57746 4094
rect 57774 4093 57777 4094
rect 57654 4067 57655 4093
rect 57745 4067 57746 4093
rect 57623 4066 57626 4067
rect 57654 4066 57666 4067
rect 57694 4066 57706 4067
rect 57734 4066 57746 4067
rect 57774 4066 57777 4067
rect 57623 4061 57777 4066
rect 699 4027 727 4032
rect 38574 3822 38728 3826
rect 38574 3821 38577 3822
rect 38605 3821 38617 3822
rect 38645 3821 38657 3822
rect 38685 3821 38697 3822
rect 38725 3821 38728 3822
rect 38605 3795 38606 3821
rect 38696 3795 38697 3821
rect 38574 3794 38577 3795
rect 38605 3794 38617 3795
rect 38645 3794 38657 3795
rect 38685 3794 38697 3795
rect 38725 3794 38728 3795
rect 38574 3789 38728 3794
rect 19524 3550 19678 3554
rect 19524 3549 19527 3550
rect 19555 3549 19567 3550
rect 19595 3549 19607 3550
rect 19635 3549 19647 3550
rect 19675 3549 19678 3550
rect 19555 3523 19556 3549
rect 19646 3523 19647 3549
rect 19524 3522 19527 3523
rect 19555 3522 19567 3523
rect 19595 3522 19607 3523
rect 19635 3522 19647 3523
rect 19675 3522 19678 3523
rect 19524 3517 19678 3522
rect 57623 3550 57777 3554
rect 57623 3549 57626 3550
rect 57654 3549 57666 3550
rect 57694 3549 57706 3550
rect 57734 3549 57746 3550
rect 57774 3549 57777 3550
rect 57654 3523 57655 3549
rect 57745 3523 57746 3549
rect 57623 3522 57626 3523
rect 57654 3522 57666 3523
rect 57694 3522 57706 3523
rect 57734 3522 57746 3523
rect 57774 3522 57777 3523
rect 57623 3517 57777 3522
rect 38574 3278 38728 3282
rect 38574 3277 38577 3278
rect 38605 3277 38617 3278
rect 38645 3277 38657 3278
rect 38685 3277 38697 3278
rect 38725 3277 38728 3278
rect 38605 3251 38606 3277
rect 38696 3251 38697 3277
rect 38574 3250 38577 3251
rect 38605 3250 38617 3251
rect 38645 3250 38657 3251
rect 38685 3250 38697 3251
rect 38725 3250 38728 3251
rect 38574 3245 38728 3250
rect 19524 3006 19678 3010
rect 19524 3005 19527 3006
rect 19555 3005 19567 3006
rect 19595 3005 19607 3006
rect 19635 3005 19647 3006
rect 19675 3005 19678 3006
rect 19555 2979 19556 3005
rect 19646 2979 19647 3005
rect 19524 2978 19527 2979
rect 19555 2978 19567 2979
rect 19595 2978 19607 2979
rect 19635 2978 19647 2979
rect 19675 2978 19678 2979
rect 19524 2973 19678 2978
rect 57623 3006 57777 3010
rect 57623 3005 57626 3006
rect 57654 3005 57666 3006
rect 57694 3005 57706 3006
rect 57734 3005 57746 3006
rect 57774 3005 57777 3006
rect 57654 2979 57655 3005
rect 57745 2979 57746 3005
rect 57623 2978 57626 2979
rect 57654 2978 57666 2979
rect 57694 2978 57706 2979
rect 57734 2978 57746 2979
rect 57774 2978 57777 2979
rect 57623 2973 57777 2978
rect 38574 2734 38728 2738
rect 38574 2733 38577 2734
rect 38605 2733 38617 2734
rect 38645 2733 38657 2734
rect 38685 2733 38697 2734
rect 38725 2733 38728 2734
rect 38605 2707 38606 2733
rect 38696 2707 38697 2733
rect 38574 2706 38577 2707
rect 38605 2706 38617 2707
rect 38645 2706 38657 2707
rect 38685 2706 38697 2707
rect 38725 2706 38728 2707
rect 38574 2701 38728 2706
rect 19524 2462 19678 2466
rect 19524 2461 19527 2462
rect 19555 2461 19567 2462
rect 19595 2461 19607 2462
rect 19635 2461 19647 2462
rect 19675 2461 19678 2462
rect 19555 2435 19556 2461
rect 19646 2435 19647 2461
rect 19524 2434 19527 2435
rect 19555 2434 19567 2435
rect 19595 2434 19607 2435
rect 19635 2434 19647 2435
rect 19675 2434 19678 2435
rect 19524 2429 19678 2434
rect 57623 2462 57777 2466
rect 57623 2461 57626 2462
rect 57654 2461 57666 2462
rect 57694 2461 57706 2462
rect 57734 2461 57746 2462
rect 57774 2461 57777 2462
rect 57654 2435 57655 2461
rect 57745 2435 57746 2461
rect 57623 2434 57626 2435
rect 57654 2434 57666 2435
rect 57694 2434 57706 2435
rect 57734 2434 57746 2435
rect 57774 2434 57777 2435
rect 57623 2429 57777 2434
rect 38574 2190 38728 2194
rect 38574 2189 38577 2190
rect 38605 2189 38617 2190
rect 38645 2189 38657 2190
rect 38685 2189 38697 2190
rect 38725 2189 38728 2190
rect 38605 2163 38606 2189
rect 38696 2163 38697 2189
rect 38574 2162 38577 2163
rect 38605 2162 38617 2163
rect 38645 2162 38657 2163
rect 38685 2162 38697 2163
rect 38725 2162 38728 2163
rect 38574 2157 38728 2162
rect 19524 1918 19678 1922
rect 19524 1917 19527 1918
rect 19555 1917 19567 1918
rect 19595 1917 19607 1918
rect 19635 1917 19647 1918
rect 19675 1917 19678 1918
rect 19555 1891 19556 1917
rect 19646 1891 19647 1917
rect 19524 1890 19527 1891
rect 19555 1890 19567 1891
rect 19595 1890 19607 1891
rect 19635 1890 19647 1891
rect 19675 1890 19678 1891
rect 19524 1885 19678 1890
rect 57623 1918 57777 1922
rect 57623 1917 57626 1918
rect 57654 1917 57666 1918
rect 57694 1917 57706 1918
rect 57734 1917 57746 1918
rect 57774 1917 57777 1918
rect 57654 1891 57655 1917
rect 57745 1891 57746 1917
rect 57623 1890 57626 1891
rect 57654 1890 57666 1891
rect 57694 1890 57706 1891
rect 57734 1890 57746 1891
rect 57774 1890 57777 1891
rect 57623 1885 57777 1890
rect 38574 1646 38728 1650
rect 38574 1645 38577 1646
rect 38605 1645 38617 1646
rect 38645 1645 38657 1646
rect 38685 1645 38697 1646
rect 38725 1645 38728 1646
rect 38605 1619 38606 1645
rect 38696 1619 38697 1645
rect 38574 1618 38577 1619
rect 38605 1618 38617 1619
rect 38645 1618 38657 1619
rect 38685 1618 38697 1619
rect 38725 1618 38728 1619
rect 38574 1613 38728 1618
rect 19524 1374 19678 1378
rect 19524 1373 19527 1374
rect 19555 1373 19567 1374
rect 19595 1373 19607 1374
rect 19635 1373 19647 1374
rect 19675 1373 19678 1374
rect 19555 1347 19556 1373
rect 19646 1347 19647 1373
rect 19524 1346 19527 1347
rect 19555 1346 19567 1347
rect 19595 1346 19607 1347
rect 19635 1346 19647 1347
rect 19675 1346 19678 1347
rect 19524 1341 19678 1346
rect 57623 1374 57777 1378
rect 57623 1373 57626 1374
rect 57654 1373 57666 1374
rect 57694 1373 57706 1374
rect 57734 1373 57746 1374
rect 57774 1373 57777 1374
rect 57654 1347 57655 1373
rect 57745 1347 57746 1373
rect 57623 1346 57626 1347
rect 57654 1346 57666 1347
rect 57694 1346 57706 1347
rect 57734 1346 57746 1347
rect 57774 1346 57777 1347
rect 57623 1341 57777 1346
rect 74720 1325 74734 6087
rect 74760 6048 74786 6051
rect 74760 6019 74786 6022
rect 74766 5507 74780 6019
rect 74996 5915 75010 6291
rect 74990 5912 75016 5915
rect 74990 5883 75016 5886
rect 74760 5504 74786 5507
rect 74760 5475 74786 5478
rect 75180 5337 75194 6325
rect 75410 5677 75424 6733
rect 75542 6626 75568 6629
rect 75542 6597 75568 6600
rect 75548 5949 75562 6597
rect 75772 6388 75798 6391
rect 75772 6359 75798 6362
rect 75634 6320 75660 6323
rect 75634 6291 75660 6294
rect 75680 6320 75706 6323
rect 75680 6291 75706 6294
rect 75542 5946 75568 5949
rect 75542 5917 75568 5920
rect 75640 5881 75654 6291
rect 75686 6119 75700 6291
rect 75680 6116 75706 6119
rect 75680 6087 75706 6090
rect 75778 6093 75792 6359
rect 75818 6354 75844 6357
rect 75818 6325 75844 6328
rect 75824 6187 75838 6325
rect 75818 6184 75844 6187
rect 75818 6155 75844 6158
rect 75634 5878 75660 5881
rect 75634 5849 75660 5852
rect 75404 5674 75430 5677
rect 75404 5645 75430 5648
rect 75686 5609 75700 6087
rect 75778 6079 75884 6093
rect 75870 6051 75884 6079
rect 75818 6048 75844 6051
rect 75818 6019 75844 6022
rect 75864 6048 75890 6051
rect 75864 6019 75890 6022
rect 75680 5606 75706 5609
rect 75680 5577 75706 5580
rect 75824 5371 75838 6019
rect 75870 5779 75884 6019
rect 76008 5949 76022 7643
rect 77473 7600 77501 8000
rect 78991 7600 79019 8000
rect 80555 7657 80583 8000
rect 80555 7643 80668 7657
rect 80555 7600 80583 7643
rect 77480 6731 77494 7600
rect 78578 6864 78604 6867
rect 78578 6835 78604 6838
rect 77474 6728 77500 6731
rect 77474 6699 77500 6702
rect 77612 6660 77638 6663
rect 77612 6631 77638 6634
rect 77934 6660 77960 6663
rect 77934 6631 77960 6634
rect 78210 6660 78236 6663
rect 78210 6631 78236 6634
rect 76232 6626 76258 6629
rect 76232 6597 76258 6600
rect 76876 6626 76902 6629
rect 76876 6597 76902 6600
rect 77106 6626 77132 6629
rect 77106 6597 77132 6600
rect 76238 6221 76252 6597
rect 76324 6592 76350 6595
rect 76324 6563 76350 6566
rect 76330 6493 76344 6563
rect 76673 6542 76827 6546
rect 76673 6541 76676 6542
rect 76704 6541 76716 6542
rect 76744 6541 76756 6542
rect 76784 6541 76796 6542
rect 76824 6541 76827 6542
rect 76704 6515 76705 6541
rect 76795 6515 76796 6541
rect 76673 6514 76676 6515
rect 76704 6514 76716 6515
rect 76744 6514 76756 6515
rect 76784 6514 76796 6515
rect 76824 6514 76827 6515
rect 76673 6509 76827 6514
rect 76324 6490 76350 6493
rect 76324 6461 76350 6464
rect 76416 6490 76442 6493
rect 76416 6461 76442 6464
rect 76330 6416 76344 6461
rect 76284 6402 76344 6416
rect 76232 6218 76258 6221
rect 76232 6189 76258 6192
rect 76284 6051 76298 6402
rect 76370 6388 76396 6391
rect 76370 6359 76396 6362
rect 76376 6187 76390 6359
rect 76422 6357 76436 6461
rect 76416 6354 76442 6357
rect 76416 6325 76442 6328
rect 76554 6354 76580 6357
rect 76554 6325 76580 6328
rect 76370 6184 76396 6187
rect 76370 6155 76396 6158
rect 76094 6048 76120 6051
rect 76094 6019 76120 6022
rect 76278 6048 76304 6051
rect 76278 6019 76304 6022
rect 76002 5946 76028 5949
rect 76002 5917 76028 5920
rect 76100 5881 76114 6019
rect 76376 5881 76390 6155
rect 76094 5878 76120 5881
rect 76094 5849 76120 5852
rect 76370 5878 76396 5881
rect 76370 5849 76396 5852
rect 75864 5776 75890 5779
rect 75864 5747 75890 5750
rect 76560 5575 76574 6325
rect 76882 6221 76896 6597
rect 77060 6320 77086 6323
rect 77060 6291 77086 6294
rect 76876 6218 76902 6221
rect 76876 6189 76902 6192
rect 77066 6153 77080 6291
rect 77060 6150 77086 6153
rect 77060 6121 77086 6124
rect 76673 5998 76827 6002
rect 76673 5997 76676 5998
rect 76704 5997 76716 5998
rect 76744 5997 76756 5998
rect 76784 5997 76796 5998
rect 76824 5997 76827 5998
rect 76704 5971 76705 5997
rect 76795 5971 76796 5997
rect 76673 5970 76676 5971
rect 76704 5970 76716 5971
rect 76744 5970 76756 5971
rect 76784 5970 76796 5971
rect 76824 5970 76827 5971
rect 76673 5965 76827 5970
rect 77112 5949 77126 6597
rect 77618 6595 77632 6631
rect 77612 6592 77638 6595
rect 77612 6563 77638 6566
rect 77519 6440 77547 6444
rect 77940 6425 77954 6631
rect 77519 6407 77547 6412
rect 77934 6422 77960 6425
rect 77526 6391 77540 6407
rect 77934 6393 77960 6396
rect 77520 6388 77546 6391
rect 77520 6359 77546 6362
rect 77526 6187 77540 6359
rect 77520 6184 77546 6187
rect 77520 6155 77546 6158
rect 77940 6085 77954 6393
rect 78216 6085 78230 6631
rect 78302 6626 78328 6629
rect 78302 6597 78328 6600
rect 78308 6459 78322 6597
rect 78584 6493 78598 6835
rect 78998 6765 79012 7600
rect 78624 6762 78650 6765
rect 78624 6733 78650 6736
rect 78992 6762 79018 6765
rect 78992 6733 79018 6736
rect 79728 6762 79754 6765
rect 79728 6733 79754 6736
rect 78578 6490 78604 6493
rect 78578 6461 78604 6464
rect 78302 6456 78328 6459
rect 78302 6427 78328 6430
rect 78630 6221 78644 6733
rect 78900 6660 78926 6663
rect 78900 6631 78926 6634
rect 79314 6660 79340 6663
rect 79314 6631 79340 6634
rect 78906 6425 78920 6631
rect 79320 6493 79334 6631
rect 79452 6626 79478 6629
rect 79452 6597 79478 6600
rect 79314 6490 79340 6493
rect 79314 6461 79340 6464
rect 78900 6422 78926 6425
rect 78900 6393 78926 6396
rect 78946 6320 78972 6323
rect 78945 6304 78946 6308
rect 78972 6304 78973 6308
rect 78945 6271 78973 6276
rect 78624 6218 78650 6221
rect 78624 6189 78650 6192
rect 77934 6082 77960 6085
rect 77934 6053 77960 6056
rect 78210 6082 78236 6085
rect 78210 6053 78236 6056
rect 77106 5946 77132 5949
rect 77106 5917 77132 5920
rect 78216 5643 78230 6053
rect 78630 5677 78644 6189
rect 78624 5674 78650 5677
rect 78624 5645 78650 5648
rect 78210 5640 78236 5643
rect 78210 5611 78236 5614
rect 76554 5572 76580 5575
rect 76554 5543 76580 5546
rect 78072 5538 78098 5541
rect 78072 5509 78098 5512
rect 76673 5454 76827 5458
rect 76673 5453 76676 5454
rect 76704 5453 76716 5454
rect 76744 5453 76756 5454
rect 76784 5453 76796 5454
rect 76824 5453 76827 5454
rect 76704 5427 76705 5453
rect 76795 5427 76796 5453
rect 76673 5426 76676 5427
rect 76704 5426 76716 5427
rect 76744 5426 76756 5427
rect 76784 5426 76796 5427
rect 76824 5426 76827 5427
rect 76673 5421 76827 5426
rect 78078 5371 78092 5509
rect 75818 5368 75844 5371
rect 75818 5339 75844 5342
rect 78072 5368 78098 5371
rect 78072 5339 78098 5342
rect 75174 5334 75200 5337
rect 75174 5305 75200 5308
rect 78078 5031 78092 5339
rect 78072 5028 78098 5031
rect 78072 4999 78098 5002
rect 76673 4910 76827 4914
rect 76673 4909 76676 4910
rect 76704 4909 76716 4910
rect 76744 4909 76756 4910
rect 76784 4909 76796 4910
rect 76824 4909 76827 4910
rect 76704 4883 76705 4909
rect 76795 4883 76796 4909
rect 76673 4882 76676 4883
rect 76704 4882 76716 4883
rect 76744 4882 76756 4883
rect 76784 4882 76796 4883
rect 76824 4882 76827 4883
rect 76673 4877 76827 4882
rect 78078 4827 78092 4999
rect 79320 4827 79334 6461
rect 79406 6354 79432 6357
rect 79406 6325 79432 6328
rect 79412 6119 79426 6325
rect 79458 6187 79472 6597
rect 79734 6391 79748 6733
rect 80464 6694 80490 6697
rect 80464 6665 80490 6668
rect 79774 6592 79800 6595
rect 79774 6563 79800 6566
rect 80188 6592 80214 6595
rect 80188 6563 80214 6566
rect 79780 6391 79794 6563
rect 80194 6459 80208 6563
rect 80188 6456 80214 6459
rect 80188 6427 80214 6430
rect 79728 6388 79754 6391
rect 79728 6359 79754 6362
rect 79774 6388 79800 6391
rect 79774 6359 79800 6362
rect 80142 6320 80168 6323
rect 80141 6304 80142 6308
rect 80168 6304 80169 6308
rect 80141 6271 80169 6276
rect 79452 6184 79478 6187
rect 79452 6155 79478 6158
rect 80194 6153 80208 6427
rect 80470 6221 80484 6665
rect 80602 6626 80628 6629
rect 80602 6597 80628 6600
rect 80464 6218 80490 6221
rect 80464 6189 80490 6192
rect 80188 6150 80214 6153
rect 80188 6121 80214 6124
rect 79406 6116 79432 6119
rect 79406 6087 79432 6090
rect 80556 6048 80582 6051
rect 80556 6019 80582 6022
rect 80562 5881 80576 6019
rect 80556 5878 80582 5881
rect 80556 5849 80582 5852
rect 80608 5813 80622 6597
rect 80654 5813 80668 7643
rect 82073 7600 82101 8000
rect 83591 7600 83619 8000
rect 85155 7657 85183 8000
rect 86673 7657 86701 8000
rect 85155 7643 85222 7657
rect 85155 7600 85183 7643
rect 80832 6898 80858 6901
rect 80832 6869 80858 6872
rect 80786 6762 80812 6765
rect 80746 6742 80786 6756
rect 80746 6153 80760 6742
rect 80786 6733 80812 6736
rect 80838 6425 80852 6869
rect 81338 6762 81364 6765
rect 81338 6733 81364 6736
rect 81752 6762 81778 6765
rect 81752 6733 81778 6736
rect 81344 6663 81358 6733
rect 81758 6663 81772 6733
rect 81338 6660 81364 6663
rect 81338 6631 81364 6634
rect 81752 6660 81778 6663
rect 81752 6631 81778 6634
rect 81016 6592 81042 6595
rect 81016 6563 81042 6566
rect 81246 6592 81272 6595
rect 81246 6563 81272 6566
rect 80832 6422 80858 6425
rect 80832 6393 80858 6396
rect 80786 6388 80812 6391
rect 80786 6359 80812 6362
rect 80792 6221 80806 6359
rect 80786 6218 80812 6221
rect 80786 6189 80812 6192
rect 80740 6150 80766 6153
rect 80740 6121 80766 6124
rect 80878 6116 80904 6119
rect 80878 6087 80904 6090
rect 80884 5881 80898 6087
rect 81022 5949 81036 6563
rect 81062 6388 81088 6391
rect 81062 6359 81088 6362
rect 81016 5946 81042 5949
rect 81016 5917 81042 5920
rect 80878 5878 80904 5881
rect 80878 5849 80904 5852
rect 80602 5810 80628 5813
rect 80602 5781 80628 5784
rect 80648 5810 80674 5813
rect 80648 5781 80674 5784
rect 81068 5677 81082 6359
rect 81252 6153 81266 6563
rect 81344 6153 81358 6631
rect 81384 6626 81410 6629
rect 81384 6597 81410 6600
rect 81246 6150 81272 6153
rect 81246 6121 81272 6124
rect 81338 6150 81364 6153
rect 81338 6121 81364 6124
rect 81292 6082 81318 6085
rect 81292 6053 81318 6056
rect 81338 6082 81364 6085
rect 81338 6053 81364 6056
rect 81108 6048 81134 6051
rect 81108 6019 81134 6022
rect 81062 5674 81088 5677
rect 81062 5645 81088 5648
rect 81114 5575 81128 6019
rect 81298 5915 81312 6053
rect 81292 5912 81318 5915
rect 81292 5883 81318 5886
rect 81344 5677 81358 6053
rect 81390 5949 81404 6597
rect 81758 6493 81772 6631
rect 81890 6626 81916 6629
rect 81890 6597 81916 6600
rect 81752 6490 81778 6493
rect 81752 6461 81778 6464
rect 81706 6456 81732 6459
rect 81706 6427 81732 6430
rect 81430 6388 81456 6391
rect 81430 6359 81456 6362
rect 81436 6051 81450 6359
rect 81430 6048 81456 6051
rect 81430 6019 81456 6022
rect 81384 5946 81410 5949
rect 81384 5917 81410 5920
rect 81712 5677 81726 6427
rect 81844 6320 81870 6323
rect 81844 6291 81870 6294
rect 81797 6168 81825 6172
rect 81797 6135 81798 6140
rect 81824 6135 81825 6140
rect 81798 6121 81824 6124
rect 81752 5844 81778 5847
rect 81752 5815 81778 5818
rect 81338 5674 81364 5677
rect 81338 5645 81364 5648
rect 81706 5674 81732 5677
rect 81706 5645 81732 5648
rect 81758 5575 81772 5815
rect 81108 5572 81134 5575
rect 81108 5543 81134 5546
rect 81752 5572 81778 5575
rect 81752 5543 81778 5546
rect 81804 5065 81818 6121
rect 81850 5881 81864 6291
rect 81896 5949 81910 6597
rect 82080 6365 82094 7600
rect 83040 6898 83066 6901
rect 83040 6869 83066 6872
rect 82626 6694 82652 6697
rect 82626 6665 82652 6668
rect 82442 6660 82468 6663
rect 82632 6637 82646 6665
rect 82442 6631 82468 6634
rect 82304 6592 82330 6595
rect 82304 6563 82330 6566
rect 82310 6391 82324 6563
rect 82304 6388 82330 6391
rect 82080 6357 82140 6365
rect 82304 6359 82330 6362
rect 82080 6354 82146 6357
rect 82080 6351 82120 6354
rect 82120 6325 82146 6328
rect 82166 6082 82192 6085
rect 82166 6053 82192 6056
rect 82172 5949 82186 6053
rect 82448 5949 82462 6631
rect 82586 6629 82646 6637
rect 82580 6626 82646 6629
rect 82606 6623 82646 6626
rect 82580 6597 82606 6600
rect 82626 6592 82652 6595
rect 82626 6563 82652 6566
rect 82672 6592 82698 6595
rect 82672 6563 82698 6566
rect 82632 6493 82646 6563
rect 82626 6490 82652 6493
rect 82626 6461 82652 6464
rect 81890 5946 81916 5949
rect 81890 5917 81916 5920
rect 82166 5946 82192 5949
rect 82166 5917 82192 5920
rect 82442 5946 82468 5949
rect 82442 5917 82468 5920
rect 81844 5878 81870 5881
rect 81844 5849 81870 5852
rect 82678 5609 82692 6563
rect 82718 6422 82744 6425
rect 82718 6393 82744 6396
rect 82724 6187 82738 6393
rect 83046 6187 83060 6869
rect 83224 6728 83250 6731
rect 83224 6699 83250 6702
rect 83230 6595 83244 6699
rect 83224 6592 83250 6595
rect 83224 6563 83250 6566
rect 83086 6422 83112 6425
rect 83086 6393 83112 6396
rect 83092 6323 83106 6393
rect 83086 6320 83112 6323
rect 83086 6291 83112 6294
rect 83230 6221 83244 6563
rect 83598 6493 83612 7600
rect 83684 6898 83710 6901
rect 83684 6869 83710 6872
rect 83690 6629 83704 6869
rect 85208 6731 85222 7643
rect 86542 7643 86701 7657
rect 86542 6731 86556 7643
rect 86673 7600 86701 7643
rect 88237 7600 88265 8000
rect 89755 7600 89783 8000
rect 91273 7657 91301 8000
rect 92837 7657 92865 8000
rect 91273 7643 91386 7657
rect 91273 7600 91301 7643
rect 87088 6898 87114 6901
rect 87088 6869 87114 6872
rect 85202 6728 85228 6731
rect 85202 6699 85228 6702
rect 86536 6728 86562 6731
rect 86536 6699 86562 6702
rect 86904 6728 86930 6731
rect 86904 6699 86930 6702
rect 83684 6626 83710 6629
rect 83684 6597 83710 6600
rect 83592 6490 83618 6493
rect 83592 6461 83618 6464
rect 86910 6459 86924 6699
rect 87094 6663 87108 6869
rect 87922 6759 88028 6773
rect 87922 6663 87936 6759
rect 88014 6731 88028 6759
rect 88192 6762 88218 6765
rect 88192 6733 88218 6736
rect 87962 6728 87988 6731
rect 87962 6699 87988 6702
rect 88008 6728 88034 6731
rect 88008 6699 88034 6702
rect 87088 6660 87114 6663
rect 87088 6631 87114 6634
rect 87916 6660 87942 6663
rect 87916 6631 87942 6634
rect 87870 6626 87896 6629
rect 87870 6597 87896 6600
rect 87502 6592 87528 6595
rect 87502 6563 87528 6566
rect 87508 6493 87522 6563
rect 87876 6493 87890 6597
rect 87502 6490 87528 6493
rect 87502 6461 87528 6464
rect 87870 6490 87896 6493
rect 87870 6461 87896 6464
rect 87968 6459 87982 6699
rect 88198 6663 88212 6733
rect 88192 6660 88218 6663
rect 88192 6631 88218 6634
rect 88198 6493 88212 6631
rect 88192 6490 88218 6493
rect 88192 6461 88218 6464
rect 86904 6456 86930 6459
rect 86904 6427 86930 6430
rect 87962 6456 87988 6459
rect 87962 6427 87988 6430
rect 88198 6425 88212 6461
rect 83270 6422 83296 6425
rect 83270 6393 83296 6396
rect 88192 6422 88218 6425
rect 88192 6393 88218 6396
rect 83224 6218 83250 6221
rect 83224 6189 83250 6192
rect 82718 6184 82744 6187
rect 82718 6155 82744 6158
rect 83040 6184 83066 6187
rect 83040 6155 83066 6158
rect 82724 5643 82738 6155
rect 83276 6085 83290 6393
rect 83316 6320 83342 6323
rect 83316 6291 83342 6294
rect 82948 6082 82974 6085
rect 82948 6053 82974 6056
rect 83270 6082 83296 6085
rect 83270 6053 83296 6056
rect 82954 5813 82968 6053
rect 83322 5881 83336 6291
rect 88244 6221 88258 7600
rect 88882 6898 88908 6901
rect 88882 6869 88908 6872
rect 88888 6731 88902 6869
rect 88882 6728 88908 6731
rect 88882 6699 88908 6702
rect 88836 6626 88862 6629
rect 88836 6597 88862 6600
rect 88468 6456 88494 6459
rect 88468 6427 88494 6430
rect 88376 6388 88402 6391
rect 88376 6359 88402 6362
rect 88238 6218 88264 6221
rect 88238 6189 88264 6192
rect 88330 6048 88356 6051
rect 88330 6019 88356 6022
rect 88336 5881 88350 6019
rect 88382 5949 88396 6359
rect 88474 6229 88488 6427
rect 88698 6320 88724 6323
rect 88698 6291 88724 6294
rect 88474 6215 88580 6229
rect 88566 6153 88580 6215
rect 88560 6150 88586 6153
rect 88560 6121 88586 6124
rect 88376 5946 88402 5949
rect 88376 5917 88402 5920
rect 83316 5878 83342 5881
rect 83316 5849 83342 5852
rect 88330 5878 88356 5881
rect 88330 5849 88356 5852
rect 88566 5847 88580 6121
rect 88704 5949 88718 6291
rect 88698 5946 88724 5949
rect 88698 5917 88724 5920
rect 88560 5844 88586 5847
rect 88560 5815 88586 5818
rect 82948 5810 82974 5813
rect 82948 5781 82974 5784
rect 82954 5677 82968 5781
rect 82948 5674 82974 5677
rect 82948 5645 82974 5648
rect 82718 5640 82744 5643
rect 82718 5611 82744 5614
rect 88842 5609 88856 6597
rect 88888 6187 88902 6699
rect 88974 6456 89000 6459
rect 88974 6427 89000 6430
rect 88928 6320 88954 6323
rect 88928 6291 88954 6294
rect 88882 6184 88908 6187
rect 88882 6155 88908 6158
rect 88934 6119 88948 6291
rect 88928 6116 88954 6119
rect 88928 6087 88954 6090
rect 88934 5949 88948 6087
rect 88928 5946 88954 5949
rect 88928 5917 88954 5920
rect 88980 5609 88994 6427
rect 89762 6221 89776 7600
rect 90952 6898 90978 6901
rect 90952 6869 90978 6872
rect 90216 6728 90242 6731
rect 90216 6699 90242 6702
rect 89986 6626 90012 6629
rect 89986 6597 90012 6600
rect 89940 6320 89966 6323
rect 89940 6291 89966 6294
rect 89756 6218 89782 6221
rect 89756 6189 89782 6192
rect 89572 6116 89598 6119
rect 89572 6087 89598 6090
rect 89020 6048 89046 6051
rect 89020 6019 89046 6022
rect 82672 5606 82698 5609
rect 82672 5577 82698 5580
rect 88836 5606 88862 5609
rect 88836 5577 88862 5580
rect 88974 5606 89000 5609
rect 88974 5577 89000 5580
rect 89026 5575 89040 6019
rect 89020 5572 89046 5575
rect 89020 5543 89046 5546
rect 89578 5235 89592 6087
rect 89710 6082 89736 6085
rect 89710 6053 89736 6056
rect 89716 5541 89730 6053
rect 89946 5949 89960 6291
rect 89992 5949 90006 6597
rect 90078 6490 90104 6493
rect 90078 6461 90104 6464
rect 90124 6490 90150 6493
rect 90124 6461 90150 6464
rect 90084 6391 90098 6461
rect 90078 6388 90104 6391
rect 90078 6359 90104 6362
rect 90130 6357 90144 6461
rect 90170 6422 90196 6425
rect 90170 6393 90196 6396
rect 90124 6354 90150 6357
rect 90124 6325 90150 6328
rect 90078 6048 90104 6051
rect 90078 6019 90104 6022
rect 90084 5949 90098 6019
rect 89940 5946 89966 5949
rect 89940 5917 89966 5920
rect 89986 5946 90012 5949
rect 89986 5917 90012 5920
rect 90078 5946 90104 5949
rect 90078 5917 90104 5920
rect 89940 5878 89966 5881
rect 90032 5878 90058 5881
rect 89966 5858 90032 5872
rect 89940 5849 89966 5852
rect 90032 5849 90058 5852
rect 90176 5813 90190 6393
rect 90170 5810 90196 5813
rect 90170 5781 90196 5784
rect 90222 5575 90236 6699
rect 90958 6697 90972 6869
rect 91372 6765 91386 7643
rect 92837 7643 92904 7657
rect 92837 7600 92865 7643
rect 92890 6765 92904 7643
rect 94355 7600 94383 8000
rect 95873 7657 95901 8000
rect 95650 7643 95901 7657
rect 91366 6762 91392 6765
rect 91366 6733 91392 6736
rect 92884 6762 92910 6765
rect 92884 6733 92910 6736
rect 90952 6694 90978 6697
rect 90952 6665 90978 6668
rect 91044 6694 91070 6697
rect 91044 6665 91070 6668
rect 94264 6694 94290 6697
rect 94264 6665 94290 6668
rect 90308 6660 90334 6663
rect 90308 6631 90334 6634
rect 90262 6354 90288 6357
rect 90262 6325 90288 6328
rect 90268 5779 90282 6325
rect 90314 6323 90328 6631
rect 90446 6626 90472 6629
rect 90446 6597 90472 6600
rect 90354 6592 90380 6595
rect 90354 6563 90380 6566
rect 90308 6320 90334 6323
rect 90308 6291 90334 6294
rect 90360 6119 90374 6563
rect 90452 6187 90466 6597
rect 90768 6422 90794 6425
rect 90768 6393 90794 6396
rect 90722 6320 90748 6323
rect 90722 6291 90748 6294
rect 90446 6184 90472 6187
rect 90446 6155 90472 6158
rect 90354 6116 90380 6119
rect 90354 6087 90380 6090
rect 90308 5878 90334 5881
rect 90360 5872 90374 6087
rect 90728 6085 90742 6291
rect 90722 6082 90748 6085
rect 90722 6053 90748 6056
rect 90334 5858 90374 5872
rect 90308 5849 90334 5852
rect 90774 5847 90788 6393
rect 91050 6357 91064 6665
rect 93896 6592 93922 6595
rect 93896 6563 93922 6566
rect 93988 6592 94014 6595
rect 93988 6563 94014 6566
rect 94172 6592 94198 6595
rect 94172 6563 94198 6566
rect 91044 6354 91070 6357
rect 91044 6325 91070 6328
rect 93902 6323 93916 6563
rect 93896 6320 93922 6323
rect 93896 6291 93922 6294
rect 93994 6153 94008 6563
rect 94178 6493 94192 6563
rect 94172 6490 94198 6493
rect 94172 6461 94198 6464
rect 94270 6459 94284 6665
rect 94264 6456 94290 6459
rect 94264 6427 94290 6430
rect 94172 6422 94198 6425
rect 94172 6393 94198 6396
rect 93988 6150 94014 6153
rect 93988 6121 94014 6124
rect 94178 5949 94192 6393
rect 94310 6354 94336 6357
rect 94362 6348 94376 7600
rect 94954 6932 94980 6935
rect 94954 6903 94980 6906
rect 94678 6898 94704 6901
rect 94678 6869 94704 6872
rect 94684 6765 94698 6869
rect 94678 6762 94704 6765
rect 94678 6733 94704 6736
rect 94402 6728 94428 6731
rect 94402 6699 94428 6702
rect 94408 6425 94422 6699
rect 94684 6425 94698 6733
rect 94770 6728 94796 6731
rect 94796 6708 94836 6722
rect 94770 6699 94796 6702
rect 94770 6660 94796 6663
rect 94770 6631 94796 6634
rect 94776 6595 94790 6631
rect 94770 6592 94796 6595
rect 94770 6563 94796 6566
rect 94402 6422 94428 6425
rect 94402 6393 94428 6396
rect 94678 6422 94704 6425
rect 94678 6393 94704 6396
rect 94776 6391 94790 6563
rect 94770 6388 94796 6391
rect 94770 6359 94796 6362
rect 94336 6334 94376 6348
rect 94586 6354 94612 6357
rect 94310 6325 94336 6328
rect 94586 6325 94612 6328
rect 94494 6320 94520 6323
rect 94494 6291 94520 6294
rect 94172 5946 94198 5949
rect 94172 5917 94198 5920
rect 90400 5844 90426 5847
rect 90400 5815 90426 5818
rect 90768 5844 90794 5847
rect 90768 5815 90794 5818
rect 90262 5776 90288 5779
rect 90262 5747 90288 5750
rect 90406 5609 90420 5815
rect 90400 5606 90426 5609
rect 90400 5577 90426 5580
rect 94500 5575 94514 6291
rect 94592 6221 94606 6325
rect 94822 6221 94836 6708
rect 94960 6697 94974 6903
rect 95460 6762 95486 6765
rect 95460 6733 95486 6736
rect 94954 6694 94980 6697
rect 94954 6665 94980 6668
rect 95466 6459 95480 6733
rect 95460 6456 95486 6459
rect 95460 6427 95486 6430
rect 95276 6320 95302 6323
rect 95276 6291 95302 6294
rect 94586 6218 94612 6221
rect 94586 6189 94612 6192
rect 94816 6218 94842 6221
rect 94816 6189 94842 6192
rect 94770 6116 94796 6119
rect 94770 6087 94796 6090
rect 94776 5915 94790 6087
rect 94770 5912 94796 5915
rect 94770 5883 94796 5886
rect 94815 5896 94843 5900
rect 94815 5863 94816 5868
rect 94842 5863 94843 5868
rect 94816 5849 94842 5852
rect 94724 5776 94750 5779
rect 94724 5747 94750 5750
rect 90216 5572 90242 5575
rect 90216 5543 90242 5546
rect 94494 5572 94520 5575
rect 94494 5543 94520 5546
rect 94730 5541 94744 5747
rect 89710 5538 89736 5541
rect 89710 5509 89736 5512
rect 94724 5538 94750 5541
rect 94724 5509 94750 5512
rect 95282 5337 95296 6291
rect 95414 6218 95440 6221
rect 95414 6189 95440 6192
rect 95420 6085 95434 6189
rect 95414 6082 95440 6085
rect 95414 6053 95440 6056
rect 95552 6082 95578 6085
rect 95552 6053 95578 6056
rect 95598 6082 95624 6085
rect 95598 6053 95624 6056
rect 95414 5878 95440 5881
rect 95414 5849 95440 5852
rect 95420 5575 95434 5849
rect 95322 5572 95348 5575
rect 95322 5543 95348 5546
rect 95414 5572 95440 5575
rect 95414 5543 95440 5546
rect 95276 5334 95302 5337
rect 95276 5305 95302 5308
rect 93758 5300 93784 5303
rect 93758 5271 93784 5274
rect 89572 5232 89598 5235
rect 89572 5203 89598 5206
rect 81798 5062 81824 5065
rect 81798 5033 81824 5036
rect 78072 4824 78098 4827
rect 78072 4795 78098 4798
rect 79314 4824 79340 4827
rect 79314 4795 79340 4798
rect 76673 4366 76827 4370
rect 76673 4365 76676 4366
rect 76704 4365 76716 4366
rect 76744 4365 76756 4366
rect 76784 4365 76796 4366
rect 76824 4365 76827 4366
rect 76704 4339 76705 4365
rect 76795 4339 76796 4365
rect 76673 4338 76676 4339
rect 76704 4338 76716 4339
rect 76744 4338 76756 4339
rect 76784 4338 76796 4339
rect 76824 4338 76827 4339
rect 76673 4333 76827 4338
rect 93764 4181 93778 5271
rect 95328 4827 95342 5543
rect 95558 5405 95572 6053
rect 95604 5609 95618 6053
rect 95598 5606 95624 5609
rect 95598 5577 95624 5580
rect 95552 5402 95578 5405
rect 95552 5373 95578 5376
rect 95650 5133 95664 7643
rect 95873 7600 95901 7643
rect 97437 7657 97465 8000
rect 98955 7657 98983 8000
rect 100519 7657 100547 8000
rect 97437 7643 97642 7657
rect 97437 7600 97465 7643
rect 96610 6898 96636 6901
rect 96610 6869 96636 6872
rect 95722 6814 95876 6818
rect 95722 6813 95725 6814
rect 95753 6813 95765 6814
rect 95793 6813 95805 6814
rect 95833 6813 95845 6814
rect 95873 6813 95876 6814
rect 95753 6787 95754 6813
rect 95844 6787 95845 6813
rect 95722 6786 95725 6787
rect 95753 6786 95765 6787
rect 95793 6786 95805 6787
rect 95833 6786 95845 6787
rect 95873 6786 95876 6787
rect 95722 6781 95876 6786
rect 95920 6728 95946 6731
rect 95920 6699 95946 6702
rect 95690 6592 95716 6595
rect 95690 6563 95716 6566
rect 95696 6493 95710 6563
rect 95690 6490 95716 6493
rect 95690 6461 95716 6464
rect 95874 6456 95900 6459
rect 95874 6427 95900 6430
rect 95880 6357 95894 6427
rect 95874 6354 95900 6357
rect 95874 6325 95900 6328
rect 95926 6308 95940 6699
rect 96196 6626 96222 6629
rect 96196 6597 96222 6600
rect 95966 6354 95992 6357
rect 95966 6325 95992 6328
rect 96018 6351 96170 6365
rect 95919 6304 95947 6308
rect 95722 6270 95876 6274
rect 95919 6271 95947 6276
rect 95722 6269 95725 6270
rect 95753 6269 95765 6270
rect 95793 6269 95805 6270
rect 95833 6269 95845 6270
rect 95873 6269 95876 6270
rect 95753 6243 95754 6269
rect 95844 6243 95845 6269
rect 95722 6242 95725 6243
rect 95753 6242 95765 6243
rect 95793 6242 95805 6243
rect 95833 6242 95845 6243
rect 95873 6242 95876 6243
rect 95722 6237 95876 6242
rect 95972 6217 95986 6325
rect 96018 6323 96032 6351
rect 96012 6320 96038 6323
rect 96012 6291 96038 6294
rect 96058 6320 96084 6323
rect 96058 6291 96084 6294
rect 96103 6304 96131 6308
rect 96064 6217 96078 6291
rect 96103 6271 96131 6276
rect 95880 6203 95986 6217
rect 96018 6203 96078 6217
rect 95880 5949 95894 6203
rect 95920 6150 95946 6153
rect 95920 6121 95946 6124
rect 95926 5949 95940 6121
rect 95874 5946 95900 5949
rect 95874 5917 95900 5920
rect 95920 5946 95946 5949
rect 95920 5917 95946 5920
rect 95926 5881 95940 5917
rect 95920 5878 95946 5881
rect 95920 5849 95946 5852
rect 95722 5726 95876 5730
rect 95722 5725 95725 5726
rect 95753 5725 95765 5726
rect 95793 5725 95805 5726
rect 95833 5725 95845 5726
rect 95873 5725 95876 5726
rect 95753 5699 95754 5725
rect 95844 5699 95845 5725
rect 95722 5698 95725 5699
rect 95753 5698 95765 5699
rect 95793 5698 95805 5699
rect 95833 5698 95845 5699
rect 95873 5698 95876 5699
rect 95722 5693 95876 5698
rect 95926 5609 95940 5849
rect 96018 5617 96032 6203
rect 96058 5844 96084 5847
rect 96058 5815 96084 5818
rect 95920 5606 95946 5609
rect 95920 5577 95946 5580
rect 95972 5603 96032 5617
rect 95972 5575 95986 5603
rect 95966 5572 95992 5575
rect 95966 5543 95992 5546
rect 96064 5269 96078 5815
rect 96110 5371 96124 6271
rect 96104 5368 96130 5371
rect 96104 5339 96130 5342
rect 96156 5337 96170 6351
rect 96202 6217 96216 6597
rect 96242 6490 96268 6493
rect 96242 6461 96268 6464
rect 96248 6357 96262 6461
rect 96288 6422 96314 6425
rect 96288 6393 96314 6396
rect 96242 6354 96268 6357
rect 96242 6325 96268 6328
rect 96202 6203 96262 6217
rect 96150 5334 96176 5337
rect 96150 5305 96176 5308
rect 96058 5266 96084 5269
rect 96058 5237 96084 5240
rect 95722 5182 95876 5186
rect 95722 5181 95725 5182
rect 95753 5181 95765 5182
rect 95793 5181 95805 5182
rect 95833 5181 95845 5182
rect 95873 5181 95876 5182
rect 95753 5155 95754 5181
rect 95844 5155 95845 5181
rect 95722 5154 95725 5155
rect 95753 5154 95765 5155
rect 95793 5154 95805 5155
rect 95833 5154 95845 5155
rect 95873 5154 95876 5155
rect 95722 5149 95876 5154
rect 96248 5133 96262 6203
rect 96294 6187 96308 6393
rect 96334 6388 96360 6391
rect 96334 6359 96360 6362
rect 96518 6388 96544 6391
rect 96518 6359 96544 6362
rect 96288 6184 96314 6187
rect 96288 6155 96314 6158
rect 95644 5130 95670 5133
rect 95644 5101 95670 5104
rect 96242 5130 96268 5133
rect 96242 5101 96268 5104
rect 96294 5031 96308 6155
rect 96340 6153 96354 6359
rect 96524 6323 96538 6359
rect 96518 6320 96544 6323
rect 96518 6291 96544 6294
rect 96524 6172 96538 6291
rect 96517 6168 96545 6172
rect 96334 6150 96360 6153
rect 96517 6135 96545 6140
rect 96334 6121 96360 6124
rect 96518 6048 96544 6051
rect 96518 6019 96544 6022
rect 96524 5900 96538 6019
rect 96517 5896 96545 5900
rect 96517 5863 96545 5868
rect 96616 5371 96630 6869
rect 96748 6762 96774 6765
rect 96748 6733 96774 6736
rect 96702 6626 96728 6629
rect 96702 6597 96728 6600
rect 96708 6217 96722 6597
rect 96662 6203 96722 6217
rect 96662 5779 96676 6203
rect 96702 6082 96728 6085
rect 96702 6053 96728 6056
rect 96656 5776 96682 5779
rect 96656 5747 96682 5750
rect 96708 5685 96722 6053
rect 96754 6025 96768 6733
rect 96978 6626 97004 6629
rect 96978 6597 97004 6600
rect 97300 6626 97326 6629
rect 97300 6597 97326 6600
rect 97392 6626 97418 6629
rect 97392 6597 97418 6600
rect 96984 6493 96998 6597
rect 97306 6569 97320 6597
rect 97260 6555 97320 6569
rect 96978 6490 97004 6493
rect 96978 6461 97004 6464
rect 97208 6320 97234 6323
rect 97208 6291 97234 6294
rect 97024 6218 97050 6221
rect 97214 6217 97228 6291
rect 97050 6203 97228 6217
rect 97024 6189 97050 6192
rect 97208 6116 97234 6119
rect 97208 6087 97234 6090
rect 96840 6048 96866 6051
rect 96754 6022 96840 6025
rect 96754 6019 96866 6022
rect 96754 6011 96860 6019
rect 96754 5779 96768 6011
rect 97214 5949 97228 6087
rect 97208 5946 97234 5949
rect 97208 5917 97234 5920
rect 96932 5912 96958 5915
rect 96932 5883 96958 5886
rect 96748 5776 96774 5779
rect 96748 5747 96774 5750
rect 96708 5671 96768 5685
rect 96754 5609 96768 5671
rect 96748 5606 96774 5609
rect 96748 5577 96774 5580
rect 96656 5538 96682 5541
rect 96656 5509 96682 5512
rect 96610 5368 96636 5371
rect 96610 5339 96636 5342
rect 96288 5028 96314 5031
rect 96288 4999 96314 5002
rect 96662 4827 96676 5509
rect 96938 5405 96952 5883
rect 97162 5844 97188 5847
rect 97162 5815 97188 5818
rect 97208 5844 97234 5847
rect 97208 5815 97234 5818
rect 96932 5402 96958 5405
rect 96932 5373 96958 5376
rect 97070 5334 97096 5337
rect 97070 5305 97096 5308
rect 95322 4824 95348 4827
rect 95322 4795 95348 4798
rect 96656 4824 96682 4827
rect 96656 4795 96682 4798
rect 97076 4793 97090 5305
rect 97168 4963 97182 5815
rect 97214 5609 97228 5815
rect 97208 5606 97234 5609
rect 97208 5577 97234 5580
rect 97208 5504 97234 5507
rect 97208 5475 97234 5478
rect 97214 5031 97228 5475
rect 97208 5028 97234 5031
rect 97208 4999 97234 5002
rect 97162 4960 97188 4963
rect 97162 4931 97188 4934
rect 97070 4790 97096 4793
rect 97070 4761 97096 4764
rect 97260 4725 97274 6555
rect 97299 6440 97327 6444
rect 97299 6407 97327 6412
rect 97306 5609 97320 6407
rect 97398 6391 97412 6597
rect 97438 6490 97464 6493
rect 97438 6461 97464 6464
rect 97392 6388 97418 6391
rect 97392 6359 97418 6362
rect 97346 6082 97372 6085
rect 97346 6053 97372 6056
rect 97352 5949 97366 6053
rect 97346 5946 97372 5949
rect 97346 5917 97372 5920
rect 97300 5606 97326 5609
rect 97300 5577 97326 5580
rect 97444 5575 97458 6461
rect 97530 6422 97556 6425
rect 97530 6393 97556 6396
rect 97536 6376 97550 6393
rect 97529 6372 97557 6376
rect 97529 6339 97557 6344
rect 97484 6048 97510 6051
rect 97484 6019 97510 6022
rect 97438 5572 97464 5575
rect 97438 5543 97464 5546
rect 97490 5337 97504 6019
rect 97536 5371 97550 6339
rect 97628 5541 97642 7643
rect 98955 7643 99114 7657
rect 98955 7600 98983 7643
rect 97990 6898 98016 6901
rect 97990 6869 98016 6872
rect 97996 6493 98010 6869
rect 98818 6694 98844 6697
rect 98818 6665 98844 6668
rect 98220 6626 98246 6629
rect 98220 6597 98246 6600
rect 98680 6626 98706 6629
rect 98680 6597 98706 6600
rect 97990 6490 98016 6493
rect 97990 6461 98016 6464
rect 97897 6440 97925 6444
rect 97897 6407 97925 6412
rect 97904 6391 97918 6407
rect 97898 6388 97924 6391
rect 97898 6359 97924 6362
rect 97990 6320 98016 6323
rect 97990 6291 98016 6294
rect 97898 5776 97924 5779
rect 97898 5747 97924 5750
rect 97944 5776 97970 5779
rect 97944 5747 97970 5750
rect 97904 5575 97918 5747
rect 97898 5572 97924 5575
rect 97898 5543 97924 5546
rect 97622 5538 97648 5541
rect 97622 5509 97648 5512
rect 97530 5368 97556 5371
rect 97530 5339 97556 5342
rect 97484 5334 97510 5337
rect 97484 5305 97510 5308
rect 97950 5065 97964 5747
rect 97944 5062 97970 5065
rect 97944 5033 97970 5036
rect 97996 4759 98010 6291
rect 98226 5609 98240 6597
rect 98686 6444 98700 6597
rect 98679 6440 98707 6444
rect 98679 6407 98680 6412
rect 98706 6407 98707 6412
rect 98726 6422 98752 6425
rect 98680 6393 98706 6396
rect 98726 6393 98752 6396
rect 98732 6187 98746 6393
rect 98824 6391 98838 6665
rect 98864 6592 98890 6595
rect 98864 6563 98890 6566
rect 98956 6592 98982 6595
rect 98956 6563 98982 6566
rect 98870 6493 98884 6563
rect 98864 6490 98890 6493
rect 98864 6461 98890 6464
rect 98818 6388 98844 6391
rect 98818 6359 98844 6362
rect 98726 6184 98752 6187
rect 98726 6155 98752 6158
rect 98726 6116 98752 6119
rect 98726 6087 98752 6090
rect 98404 6048 98430 6051
rect 98404 6019 98430 6022
rect 98496 6048 98522 6051
rect 98496 6019 98522 6022
rect 98680 6048 98706 6051
rect 98680 6019 98706 6022
rect 98410 5915 98424 6019
rect 98404 5912 98430 5915
rect 98404 5883 98430 5886
rect 98502 5779 98516 6019
rect 98686 5847 98700 6019
rect 98680 5844 98706 5847
rect 98680 5815 98706 5818
rect 98732 5813 98746 6087
rect 98962 5881 98976 6563
rect 99100 6323 99114 7643
rect 100519 7643 100586 7657
rect 100519 7600 100547 7643
rect 100427 6644 100455 6648
rect 100427 6611 100455 6616
rect 100434 6595 100448 6611
rect 99278 6592 99304 6595
rect 99278 6563 99304 6566
rect 100244 6592 100270 6595
rect 100244 6563 100270 6566
rect 100428 6592 100454 6595
rect 100428 6563 100454 6566
rect 99186 6422 99212 6425
rect 99186 6393 99212 6396
rect 99094 6320 99120 6323
rect 99094 6291 99120 6294
rect 99192 6119 99206 6393
rect 99284 6391 99298 6563
rect 99278 6388 99304 6391
rect 99278 6359 99304 6362
rect 100198 6388 100224 6391
rect 100198 6359 100224 6362
rect 100204 6308 100218 6359
rect 100197 6304 100225 6308
rect 100197 6271 100225 6276
rect 100250 6153 100264 6563
rect 100336 6422 100362 6425
rect 100336 6393 100362 6396
rect 100342 6217 100356 6393
rect 100572 6323 100586 7643
rect 102037 7600 102065 8000
rect 103555 7657 103583 8000
rect 105119 7657 105147 8000
rect 106637 7657 106665 8000
rect 108155 7657 108183 8000
rect 103555 7643 103668 7657
rect 103555 7600 103583 7643
rect 100980 6728 101006 6731
rect 100980 6699 101006 6702
rect 101716 6728 101742 6731
rect 101716 6699 101742 6702
rect 100750 6660 100776 6663
rect 100750 6631 100776 6634
rect 100658 6592 100684 6595
rect 100658 6563 100684 6566
rect 100664 6425 100678 6563
rect 100658 6422 100684 6425
rect 100658 6393 100684 6396
rect 100566 6320 100592 6323
rect 100566 6291 100592 6294
rect 100296 6203 100356 6217
rect 100244 6150 100270 6153
rect 100244 6121 100270 6124
rect 100296 6119 100310 6203
rect 99186 6116 99212 6119
rect 99186 6087 99212 6090
rect 100290 6116 100316 6119
rect 100290 6087 100316 6090
rect 100520 6116 100546 6119
rect 100520 6087 100546 6090
rect 100526 5881 100540 6087
rect 98956 5878 98982 5881
rect 98956 5849 98982 5852
rect 100520 5878 100546 5881
rect 100520 5849 100546 5852
rect 98726 5810 98752 5813
rect 98726 5781 98752 5784
rect 98496 5776 98522 5779
rect 98496 5747 98522 5750
rect 100526 5609 100540 5849
rect 100664 5847 100678 6393
rect 100658 5844 100684 5847
rect 100658 5815 100684 5818
rect 100756 5779 100770 6631
rect 100986 6323 101000 6699
rect 101026 6694 101052 6697
rect 101026 6665 101052 6668
rect 100980 6320 101006 6323
rect 100980 6291 101006 6294
rect 101032 6153 101046 6665
rect 101072 6660 101098 6663
rect 101722 6648 101736 6699
rect 101072 6631 101098 6634
rect 101715 6644 101743 6648
rect 101078 6357 101092 6631
rect 101210 6626 101236 6629
rect 101210 6597 101236 6600
rect 101578 6626 101604 6629
rect 101715 6611 101743 6616
rect 101578 6597 101604 6600
rect 101072 6354 101098 6357
rect 101072 6325 101098 6328
rect 101216 6221 101230 6597
rect 101486 6456 101512 6459
rect 101486 6427 101512 6430
rect 101492 6391 101506 6427
rect 101440 6388 101466 6391
rect 101440 6359 101466 6362
rect 101486 6388 101512 6391
rect 101486 6359 101512 6362
rect 101210 6218 101236 6221
rect 101210 6189 101236 6192
rect 101026 6150 101052 6153
rect 101026 6121 101052 6124
rect 101446 5949 101460 6359
rect 101532 6048 101558 6051
rect 101532 6019 101558 6022
rect 101440 5946 101466 5949
rect 101440 5917 101466 5920
rect 101538 5881 101552 6019
rect 101584 5915 101598 6597
rect 101670 6456 101696 6459
rect 101670 6427 101696 6430
rect 101578 5912 101604 5915
rect 101578 5883 101604 5886
rect 101532 5878 101558 5881
rect 101532 5849 101558 5852
rect 101440 5844 101466 5847
rect 101440 5815 101466 5818
rect 100750 5776 100776 5779
rect 100750 5747 100776 5750
rect 98220 5606 98246 5609
rect 98220 5577 98246 5580
rect 100520 5606 100546 5609
rect 100520 5577 100546 5580
rect 100526 5303 100540 5577
rect 101348 5572 101374 5575
rect 101446 5549 101460 5815
rect 101676 5609 101690 6427
rect 101722 6051 101736 6611
rect 101762 6150 101788 6153
rect 101762 6121 101788 6124
rect 101716 6048 101742 6051
rect 101716 6019 101742 6022
rect 101722 5813 101736 6019
rect 101768 5847 101782 6121
rect 101762 5844 101788 5847
rect 101762 5815 101788 5818
rect 101716 5810 101742 5813
rect 101716 5781 101742 5784
rect 101670 5606 101696 5609
rect 101670 5577 101696 5580
rect 101374 5546 101460 5549
rect 101348 5543 101460 5546
rect 101354 5535 101460 5543
rect 100520 5300 100546 5303
rect 100520 5271 100546 5274
rect 101768 5235 101782 5815
rect 102044 5541 102058 7600
rect 103555 6780 103583 6784
rect 103555 6747 103556 6752
rect 103582 6747 103583 6752
rect 103556 6733 103582 6736
rect 103004 6728 103030 6731
rect 102826 6702 103004 6705
rect 102826 6699 103030 6702
rect 102826 6691 103024 6699
rect 102773 6644 102801 6648
rect 102130 6626 102156 6629
rect 102130 6597 102156 6600
rect 102728 6626 102754 6629
rect 102773 6611 102801 6616
rect 102728 6597 102754 6600
rect 102084 6388 102110 6391
rect 102084 6359 102110 6362
rect 102090 6217 102104 6359
rect 102136 6323 102150 6597
rect 102544 6388 102570 6391
rect 102544 6359 102570 6362
rect 102590 6388 102616 6391
rect 102590 6359 102616 6362
rect 102130 6320 102156 6323
rect 102130 6291 102156 6294
rect 102268 6320 102294 6323
rect 102268 6291 102294 6294
rect 102090 6203 102150 6217
rect 102136 6051 102150 6203
rect 102274 6119 102288 6291
rect 102268 6116 102294 6119
rect 102268 6087 102294 6090
rect 102130 6048 102156 6051
rect 102130 6019 102156 6022
rect 102274 5949 102288 6087
rect 102498 6082 102524 6085
rect 102498 6053 102524 6056
rect 102268 5946 102294 5949
rect 102268 5917 102294 5920
rect 102452 5810 102478 5813
rect 102452 5781 102478 5784
rect 102406 5776 102432 5779
rect 102406 5747 102432 5750
rect 102038 5538 102064 5541
rect 102038 5509 102064 5512
rect 102412 5337 102426 5747
rect 102458 5575 102472 5781
rect 102504 5609 102518 6053
rect 102498 5606 102524 5609
rect 102498 5577 102524 5580
rect 102452 5572 102478 5575
rect 102452 5543 102478 5546
rect 102550 5405 102564 6359
rect 102596 6323 102610 6359
rect 102590 6320 102616 6323
rect 102636 6320 102662 6323
rect 102590 6291 102616 6294
rect 102635 6304 102636 6308
rect 102662 6304 102663 6308
rect 102635 6271 102663 6276
rect 102734 5541 102748 6597
rect 102780 5915 102794 6611
rect 102826 6595 102840 6691
rect 103602 6660 103628 6663
rect 102865 6644 102893 6648
rect 103601 6644 103602 6648
rect 103628 6644 103629 6648
rect 102865 6611 102893 6616
rect 103188 6626 103214 6629
rect 102872 6595 102886 6611
rect 103601 6611 103629 6616
rect 103188 6597 103214 6600
rect 102820 6592 102846 6595
rect 102820 6563 102846 6566
rect 102866 6592 102892 6595
rect 102866 6563 102892 6566
rect 102820 6456 102846 6459
rect 102820 6427 102846 6430
rect 102826 6221 102840 6427
rect 102820 6218 102846 6221
rect 102820 6189 102846 6192
rect 102774 5912 102800 5915
rect 102774 5883 102800 5886
rect 103194 5881 103208 6597
rect 103280 6490 103306 6493
rect 103280 6461 103306 6464
rect 103286 5949 103300 6461
rect 103654 6357 103668 7643
rect 105119 7643 105186 7657
rect 105119 7600 105147 7643
rect 104015 6780 104043 6784
rect 105172 6765 105186 7643
rect 106637 7643 106704 7657
rect 106637 7600 106665 7643
rect 106690 6765 106704 7643
rect 108155 7643 108222 7657
rect 108155 7600 108183 7643
rect 104015 6747 104043 6752
rect 105166 6762 105192 6765
rect 104022 6731 104036 6747
rect 105166 6733 105192 6736
rect 106684 6762 106710 6765
rect 106684 6733 106710 6736
rect 108208 6731 108222 7643
rect 109719 7600 109747 8000
rect 111237 7657 111265 8000
rect 112801 7657 112829 8000
rect 114319 7657 114347 8000
rect 115837 7657 115865 8000
rect 117401 7657 117429 8000
rect 111237 7643 111396 7657
rect 111237 7600 111265 7643
rect 109726 6731 109740 7600
rect 103878 6728 103904 6731
rect 103878 6699 103904 6702
rect 104016 6728 104042 6731
rect 106638 6728 106664 6731
rect 104016 6699 104042 6702
rect 106637 6712 106638 6716
rect 108202 6728 108228 6731
rect 106664 6712 106665 6716
rect 103786 6626 103812 6629
rect 103812 6606 103852 6620
rect 103786 6597 103812 6600
rect 103694 6592 103720 6595
rect 103694 6563 103720 6566
rect 103700 6493 103714 6563
rect 103694 6490 103720 6493
rect 103694 6461 103720 6464
rect 103838 6425 103852 6606
rect 103832 6422 103858 6425
rect 103832 6393 103858 6396
rect 103648 6354 103674 6357
rect 103648 6325 103674 6328
rect 103838 6221 103852 6393
rect 103832 6218 103858 6221
rect 103884 6217 103898 6699
rect 108202 6699 108228 6702
rect 109720 6728 109746 6731
rect 109720 6699 109746 6702
rect 109903 6712 109931 6716
rect 106637 6679 106665 6684
rect 109903 6679 109931 6684
rect 103970 6660 103996 6663
rect 103969 6644 103970 6648
rect 106776 6660 106802 6663
rect 103996 6644 103997 6648
rect 106776 6631 106802 6634
rect 108294 6660 108320 6663
rect 108294 6631 108320 6634
rect 103969 6611 103997 6616
rect 106782 6595 106796 6631
rect 106776 6592 106802 6595
rect 106776 6563 106802 6566
rect 103924 6490 103950 6493
rect 103924 6461 103950 6464
rect 103930 6376 103944 6461
rect 105304 6456 105330 6459
rect 105304 6427 105330 6430
rect 103923 6372 103951 6376
rect 103923 6339 103951 6344
rect 105310 6323 105324 6427
rect 108300 6425 108314 6631
rect 109910 6493 109924 6679
rect 111382 6595 111396 7643
rect 112801 7643 112868 7657
rect 112801 7600 112829 7643
rect 112026 6759 112224 6773
rect 112026 6697 112040 6759
rect 112066 6728 112092 6731
rect 112066 6699 112092 6702
rect 112020 6694 112046 6697
rect 112020 6665 112046 6668
rect 112026 6595 112040 6665
rect 112072 6595 112086 6699
rect 112210 6697 112224 6759
rect 112204 6694 112230 6697
rect 112204 6665 112230 6668
rect 112118 6629 112224 6637
rect 112112 6626 112230 6629
rect 112138 6623 112204 6626
rect 112112 6597 112138 6600
rect 112204 6597 112230 6600
rect 112854 6595 112868 7643
rect 114319 7643 114432 7657
rect 114319 7600 114347 7643
rect 113222 6759 113604 6773
rect 113222 6731 113236 6759
rect 113216 6728 113242 6731
rect 113216 6699 113242 6702
rect 113308 6728 113334 6731
rect 113308 6699 113334 6702
rect 113446 6728 113472 6731
rect 113446 6699 113472 6702
rect 113537 6712 113565 6716
rect 111376 6592 111402 6595
rect 111376 6563 111402 6566
rect 111836 6592 111862 6595
rect 111836 6563 111862 6566
rect 112020 6592 112046 6595
rect 112020 6563 112046 6566
rect 112066 6592 112092 6595
rect 112710 6592 112736 6595
rect 112066 6563 112092 6566
rect 112709 6576 112710 6580
rect 112848 6592 112874 6595
rect 112736 6576 112737 6580
rect 109904 6490 109930 6493
rect 109904 6461 109930 6464
rect 111842 6425 111856 6563
rect 112848 6563 112874 6566
rect 112709 6543 112737 6548
rect 113314 6433 113328 6699
rect 113314 6425 113420 6433
rect 108294 6422 108320 6425
rect 108294 6393 108320 6396
rect 109904 6422 109930 6425
rect 109904 6393 109930 6396
rect 111836 6422 111862 6425
rect 113314 6422 113426 6425
rect 113314 6419 113400 6422
rect 111836 6393 111862 6396
rect 113400 6393 113426 6396
rect 109910 6357 109924 6393
rect 109904 6354 109930 6357
rect 109904 6325 109930 6328
rect 113452 6323 113466 6699
rect 113590 6697 113604 6759
rect 113952 6728 113978 6731
rect 113978 6702 114018 6705
rect 113952 6699 114018 6702
rect 113537 6679 113538 6684
rect 113564 6679 113565 6684
rect 113584 6694 113610 6697
rect 113538 6665 113564 6668
rect 113958 6691 114018 6699
rect 113584 6665 113610 6668
rect 113538 6592 113564 6595
rect 113537 6576 113538 6580
rect 113564 6576 113565 6580
rect 113590 6569 113604 6665
rect 113860 6660 113886 6663
rect 113860 6631 113886 6634
rect 114004 6637 114018 6691
rect 113814 6592 113840 6595
rect 113590 6555 113650 6569
rect 113814 6563 113840 6566
rect 113537 6543 113565 6548
rect 105304 6320 105330 6323
rect 105304 6291 105330 6294
rect 113446 6320 113472 6323
rect 113446 6291 113472 6294
rect 103884 6203 103944 6217
rect 103832 6189 103858 6192
rect 103280 5946 103306 5949
rect 103280 5917 103306 5920
rect 103188 5878 103214 5881
rect 103188 5849 103214 5852
rect 103930 5847 103944 6203
rect 113636 5847 113650 6555
rect 113820 6365 113834 6563
rect 113866 6433 113880 6631
rect 114004 6629 114064 6637
rect 114004 6626 114070 6629
rect 114004 6623 114044 6626
rect 114044 6597 114070 6600
rect 113952 6592 113978 6595
rect 113952 6563 113978 6566
rect 113866 6419 113926 6433
rect 113958 6425 113972 6563
rect 114136 6456 114162 6459
rect 114136 6427 114162 6430
rect 113820 6351 113880 6365
rect 113866 5915 113880 6351
rect 113912 5949 113926 6419
rect 113952 6422 113978 6425
rect 113952 6393 113978 6396
rect 114142 6391 114156 6427
rect 114136 6388 114162 6391
rect 114136 6359 114162 6362
rect 114418 6187 114432 7643
rect 115837 7643 115904 7657
rect 115837 7600 115865 7643
rect 115890 6841 115904 7643
rect 117401 7643 117468 7657
rect 117401 7600 117429 7643
rect 115890 6827 116042 6841
rect 114596 6728 114622 6731
rect 114595 6712 114596 6716
rect 114622 6712 114623 6716
rect 114595 6679 114623 6684
rect 115890 6697 115996 6705
rect 115890 6694 116002 6697
rect 115890 6691 115976 6694
rect 115194 6660 115220 6663
rect 115193 6644 115194 6648
rect 115220 6644 115221 6648
rect 115193 6611 115221 6616
rect 115378 6626 115404 6629
rect 115378 6597 115404 6600
rect 114772 6542 114926 6546
rect 114772 6541 114775 6542
rect 114803 6541 114815 6542
rect 114843 6541 114855 6542
rect 114883 6541 114895 6542
rect 114923 6541 114926 6542
rect 114803 6515 114804 6541
rect 114894 6515 114895 6541
rect 114772 6514 114775 6515
rect 114803 6514 114815 6515
rect 114843 6514 114855 6515
rect 114883 6514 114895 6515
rect 114923 6514 114926 6515
rect 114772 6509 114926 6514
rect 115194 6456 115220 6459
rect 115194 6427 115220 6430
rect 115148 6422 115174 6425
rect 115148 6393 115174 6396
rect 115102 6388 115128 6391
rect 115102 6359 115128 6362
rect 115108 6323 115122 6359
rect 114780 6320 114806 6323
rect 114780 6291 114806 6294
rect 115056 6320 115082 6323
rect 115056 6291 115082 6294
rect 115102 6320 115128 6323
rect 115102 6291 115128 6294
rect 114412 6184 114438 6187
rect 114412 6155 114438 6158
rect 114412 6048 114438 6051
rect 114786 6042 114800 6291
rect 115062 6221 115076 6291
rect 115056 6218 115082 6221
rect 115056 6189 115082 6192
rect 114964 6116 114990 6119
rect 114964 6087 114990 6090
rect 114412 6019 114438 6022
rect 114740 6028 114800 6042
rect 114418 5949 114432 6019
rect 113906 5946 113932 5949
rect 113906 5917 113932 5920
rect 114412 5946 114438 5949
rect 114412 5917 114438 5920
rect 113860 5912 113886 5915
rect 114740 5889 114754 6028
rect 114772 5998 114926 6002
rect 114772 5997 114775 5998
rect 114803 5997 114815 5998
rect 114843 5997 114855 5998
rect 114883 5997 114895 5998
rect 114923 5997 114926 5998
rect 114803 5971 114804 5997
rect 114894 5971 114895 5997
rect 114772 5970 114775 5971
rect 114803 5970 114815 5971
rect 114843 5970 114855 5971
rect 114883 5970 114895 5971
rect 114923 5970 114926 5971
rect 114772 5965 114926 5970
rect 114970 5949 114984 6087
rect 114964 5946 114990 5949
rect 114964 5917 114990 5920
rect 113860 5883 113886 5886
rect 114694 5881 114754 5889
rect 114688 5878 114754 5881
rect 114714 5875 114754 5878
rect 114688 5849 114714 5852
rect 103924 5844 103950 5847
rect 103924 5815 103950 5818
rect 113630 5844 113656 5847
rect 113630 5815 113656 5818
rect 115154 5813 115168 6393
rect 115200 5949 115214 6427
rect 115194 5946 115220 5949
rect 115194 5917 115220 5920
rect 115148 5810 115174 5813
rect 115148 5781 115174 5784
rect 114688 5776 114714 5779
rect 114688 5747 114714 5750
rect 114694 5575 114708 5747
rect 114688 5572 114714 5575
rect 114688 5543 114714 5546
rect 115384 5541 115398 6597
rect 115516 6456 115542 6459
rect 115516 6427 115542 6430
rect 115424 6082 115450 6085
rect 115424 6053 115450 6056
rect 115430 5915 115444 6053
rect 115522 5949 115536 6427
rect 115562 6184 115588 6187
rect 115562 6155 115588 6158
rect 115568 6085 115582 6155
rect 115838 6150 115864 6153
rect 115838 6121 115864 6124
rect 115654 6116 115680 6119
rect 115654 6087 115680 6090
rect 115562 6082 115588 6085
rect 115562 6053 115588 6056
rect 115608 6048 115634 6051
rect 115660 6042 115674 6087
rect 115700 6048 115726 6051
rect 115660 6028 115700 6042
rect 115608 6019 115634 6022
rect 115700 6019 115726 6022
rect 115516 5946 115542 5949
rect 115516 5917 115542 5920
rect 115424 5912 115450 5915
rect 115424 5883 115450 5886
rect 115614 5881 115628 6019
rect 115844 5949 115858 6121
rect 115890 6051 115904 6691
rect 115976 6665 116002 6668
rect 116028 6663 116042 6827
rect 116574 6694 116600 6697
rect 116574 6665 116600 6668
rect 116666 6694 116692 6697
rect 116666 6665 116692 6668
rect 115930 6660 115956 6663
rect 115930 6631 115956 6634
rect 116022 6660 116048 6663
rect 116528 6660 116554 6663
rect 116022 6631 116048 6634
rect 116067 6644 116095 6648
rect 115936 6221 115950 6631
rect 116528 6631 116554 6634
rect 116067 6611 116095 6616
rect 116074 6595 116088 6611
rect 116068 6592 116094 6595
rect 116068 6563 116094 6566
rect 116160 6456 116186 6459
rect 116160 6427 116186 6430
rect 116166 6323 116180 6427
rect 116534 6425 116548 6631
rect 116580 6586 116594 6665
rect 116620 6592 116646 6595
rect 116580 6572 116620 6586
rect 116620 6563 116646 6566
rect 116672 6501 116686 6665
rect 117454 6595 117468 7643
rect 118919 7600 118947 8000
rect 120437 7657 120465 8000
rect 122001 7657 122029 8000
rect 123519 7657 123547 8000
rect 125037 7657 125065 8000
rect 120437 7643 120642 7657
rect 120437 7600 120465 7643
rect 117448 6592 117474 6595
rect 117448 6563 117474 6566
rect 118506 6592 118532 6595
rect 118506 6563 118532 6566
rect 116580 6487 116686 6501
rect 116528 6422 116554 6425
rect 116528 6393 116554 6396
rect 116160 6320 116186 6323
rect 116160 6291 116186 6294
rect 116252 6320 116278 6323
rect 116252 6291 116278 6294
rect 115930 6218 115956 6221
rect 115930 6189 115956 6192
rect 116258 6187 116272 6291
rect 116252 6184 116278 6187
rect 116252 6155 116278 6158
rect 116534 6119 116548 6393
rect 116580 6323 116594 6487
rect 118512 6425 118526 6563
rect 118506 6422 118532 6425
rect 118506 6393 118532 6396
rect 118926 6357 118940 7600
rect 119748 6728 119774 6731
rect 119057 6712 119085 6716
rect 118966 6694 118992 6697
rect 119057 6679 119058 6684
rect 118966 6665 118992 6668
rect 119084 6679 119085 6684
rect 119747 6712 119748 6716
rect 119774 6712 119775 6716
rect 119747 6679 119775 6684
rect 119058 6665 119084 6668
rect 118972 6357 118986 6665
rect 119104 6660 119130 6663
rect 119104 6631 119130 6634
rect 119110 6493 119124 6631
rect 119242 6626 119268 6629
rect 119242 6597 119268 6600
rect 119104 6490 119130 6493
rect 119104 6461 119130 6464
rect 119150 6456 119176 6459
rect 119150 6427 119176 6430
rect 119156 6376 119170 6427
rect 119196 6422 119222 6425
rect 119196 6393 119222 6396
rect 119149 6372 119177 6376
rect 118920 6354 118946 6357
rect 118920 6325 118946 6328
rect 118966 6354 118992 6357
rect 119149 6339 119177 6344
rect 118966 6325 118992 6328
rect 116574 6320 116600 6323
rect 116574 6291 116600 6294
rect 119202 6119 119216 6393
rect 119248 6323 119262 6597
rect 119518 6456 119544 6459
rect 119518 6427 119544 6430
rect 119242 6320 119268 6323
rect 119242 6291 119268 6294
rect 119426 6320 119452 6323
rect 119426 6291 119452 6294
rect 119432 6153 119446 6291
rect 119524 6221 119538 6427
rect 119564 6320 119590 6323
rect 119564 6291 119590 6294
rect 119518 6218 119544 6221
rect 119518 6189 119544 6192
rect 119426 6150 119452 6153
rect 119426 6121 119452 6124
rect 119570 6119 119584 6291
rect 119656 6150 119682 6153
rect 119656 6121 119682 6124
rect 116068 6116 116094 6119
rect 116068 6087 116094 6090
rect 116528 6116 116554 6119
rect 116528 6087 116554 6090
rect 119012 6116 119038 6119
rect 119012 6087 119038 6090
rect 119196 6116 119222 6119
rect 119196 6087 119222 6090
rect 119564 6116 119590 6119
rect 119564 6087 119590 6090
rect 115884 6048 115910 6051
rect 115884 6019 115910 6022
rect 115838 5946 115864 5949
rect 115838 5917 115864 5920
rect 115608 5878 115634 5881
rect 115608 5849 115634 5852
rect 115844 5779 115858 5917
rect 116074 5813 116088 6087
rect 116534 6051 116548 6087
rect 116528 6048 116554 6051
rect 116528 6019 116554 6022
rect 116068 5810 116094 5813
rect 116068 5781 116094 5784
rect 115838 5776 115864 5779
rect 115838 5747 115864 5750
rect 119018 5609 119032 6087
rect 119662 5847 119676 6121
rect 119754 6119 119768 6679
rect 119886 6660 119912 6663
rect 119886 6631 119912 6634
rect 119748 6116 119774 6119
rect 119748 6087 119774 6090
rect 119656 5844 119682 5847
rect 119656 5815 119682 5818
rect 119702 5776 119728 5779
rect 119702 5747 119728 5750
rect 119708 5677 119722 5747
rect 119892 5677 119906 6631
rect 120530 6626 120556 6629
rect 120530 6597 120556 6600
rect 120024 6456 120050 6459
rect 120024 6427 120050 6430
rect 120484 6456 120510 6459
rect 120484 6427 120510 6430
rect 119978 6150 120004 6153
rect 119978 6121 120004 6124
rect 119984 5847 119998 6121
rect 119978 5844 120004 5847
rect 119978 5815 120004 5818
rect 120030 5677 120044 6427
rect 120162 6320 120188 6323
rect 120162 6291 120188 6294
rect 120070 6218 120096 6221
rect 120070 6189 120096 6192
rect 120076 5915 120090 6189
rect 120168 5949 120182 6291
rect 120438 6048 120464 6051
rect 120438 6019 120464 6022
rect 120162 5946 120188 5949
rect 120162 5917 120188 5920
rect 120070 5912 120096 5915
rect 120070 5883 120096 5886
rect 119702 5674 119728 5677
rect 119702 5645 119728 5648
rect 119886 5674 119912 5677
rect 119886 5645 119912 5648
rect 120024 5674 120050 5677
rect 120024 5645 120050 5648
rect 119012 5606 119038 5609
rect 119012 5577 119038 5580
rect 120444 5575 120458 6019
rect 120490 5677 120504 6427
rect 120536 5949 120550 6597
rect 120530 5946 120556 5949
rect 120530 5917 120556 5920
rect 120628 5779 120642 7643
rect 122001 7643 122114 7657
rect 122001 7600 122029 7643
rect 122048 6694 122074 6697
rect 122048 6665 122074 6668
rect 120898 6626 120924 6629
rect 120898 6597 120924 6600
rect 121818 6626 121844 6629
rect 121818 6597 121844 6600
rect 120760 6048 120786 6051
rect 120760 6019 120786 6022
rect 120766 5915 120780 6019
rect 120904 5949 120918 6597
rect 121266 6592 121292 6595
rect 121266 6563 121292 6566
rect 121036 6422 121062 6425
rect 121036 6393 121062 6396
rect 121128 6422 121154 6425
rect 121128 6393 121154 6396
rect 120898 5946 120924 5949
rect 120898 5917 120924 5920
rect 120760 5912 120786 5915
rect 120760 5883 120786 5886
rect 120990 5844 121016 5847
rect 120990 5815 121016 5818
rect 120622 5776 120648 5779
rect 120622 5747 120648 5750
rect 120484 5674 120510 5677
rect 120484 5645 120510 5648
rect 120996 5575 121010 5815
rect 121042 5677 121056 6393
rect 121081 6372 121109 6376
rect 121081 6339 121082 6344
rect 121108 6339 121109 6344
rect 121082 6325 121108 6328
rect 121134 6187 121148 6393
rect 121220 6320 121246 6323
rect 121220 6291 121246 6294
rect 121128 6184 121154 6187
rect 121128 6155 121154 6158
rect 121226 6153 121240 6291
rect 121220 6150 121246 6153
rect 121220 6121 121246 6124
rect 121082 6116 121108 6119
rect 121226 6093 121240 6121
rect 121108 6090 121240 6093
rect 121082 6087 121240 6090
rect 121088 6079 121240 6087
rect 121272 6051 121286 6563
rect 121450 6320 121476 6323
rect 121450 6291 121476 6294
rect 121456 6153 121470 6291
rect 121824 6221 121838 6597
rect 121818 6218 121844 6221
rect 121818 6189 121844 6192
rect 121496 6184 121522 6187
rect 121522 6158 121608 6161
rect 121496 6155 121608 6158
rect 121502 6153 121608 6155
rect 121450 6150 121476 6153
rect 121502 6150 121614 6153
rect 121502 6147 121588 6150
rect 121450 6121 121476 6124
rect 121588 6121 121614 6124
rect 122054 6051 122068 6665
rect 122100 6221 122114 7643
rect 123519 7643 123586 7657
rect 123519 7600 123547 7643
rect 123572 6731 123586 7643
rect 125037 7643 125104 7657
rect 125037 7600 125065 7643
rect 122324 6728 122350 6731
rect 122324 6699 122350 6702
rect 122692 6728 122718 6731
rect 122692 6699 122718 6702
rect 123566 6728 123592 6731
rect 123566 6699 123592 6702
rect 122330 6501 122344 6699
rect 122462 6626 122488 6629
rect 122462 6597 122488 6600
rect 122284 6487 122344 6501
rect 122284 6425 122298 6487
rect 122468 6459 122482 6597
rect 122698 6459 122712 6699
rect 122324 6456 122350 6459
rect 122324 6427 122350 6430
rect 122462 6456 122488 6459
rect 122462 6427 122488 6430
rect 122692 6456 122718 6459
rect 122692 6427 122718 6430
rect 122278 6422 122304 6425
rect 122278 6393 122304 6396
rect 122094 6218 122120 6221
rect 122094 6189 122120 6192
rect 121266 6048 121292 6051
rect 121266 6019 121292 6022
rect 122048 6048 122074 6051
rect 122048 6019 122074 6022
rect 121272 5881 121286 6019
rect 121266 5878 121292 5881
rect 121266 5849 121292 5852
rect 122284 5847 122298 6393
rect 122330 6357 122344 6427
rect 122416 6422 122442 6425
rect 122416 6393 122442 6396
rect 122324 6354 122350 6357
rect 122324 6325 122350 6328
rect 122422 5915 122436 6393
rect 125090 6357 125104 7643
rect 126601 7600 126629 8000
rect 128119 7600 128147 8000
rect 129683 7600 129711 8000
rect 131201 7657 131229 8000
rect 131201 7643 131268 7657
rect 131201 7600 131229 7643
rect 125504 6759 125748 6773
rect 125504 6697 125518 6759
rect 125544 6728 125570 6731
rect 125570 6702 125656 6705
rect 125544 6699 125656 6702
rect 125498 6694 125524 6697
rect 125550 6691 125656 6699
rect 125498 6665 125524 6668
rect 125544 6660 125570 6663
rect 125544 6631 125570 6634
rect 125550 6493 125564 6631
rect 125590 6592 125616 6595
rect 125590 6563 125616 6566
rect 125544 6490 125570 6493
rect 125544 6461 125570 6464
rect 125596 6425 125610 6563
rect 125590 6422 125616 6425
rect 125590 6393 125616 6396
rect 124164 6354 124190 6357
rect 124164 6325 124190 6328
rect 125084 6354 125110 6357
rect 125084 6325 125110 6328
rect 124170 6153 124184 6325
rect 124164 6150 124190 6153
rect 124164 6121 124190 6124
rect 124624 6150 124650 6153
rect 124624 6121 124650 6124
rect 124630 6085 124644 6121
rect 125642 6119 125656 6691
rect 125682 6626 125708 6629
rect 125682 6597 125708 6600
rect 125688 6221 125702 6597
rect 125682 6218 125708 6221
rect 125682 6189 125708 6192
rect 125734 6187 125748 6759
rect 126234 6728 126260 6731
rect 126234 6699 126260 6702
rect 126188 6626 126214 6629
rect 126188 6597 126214 6600
rect 125820 6456 125846 6459
rect 125820 6427 125846 6430
rect 125774 6422 125800 6425
rect 125774 6393 125800 6396
rect 125728 6184 125754 6187
rect 125728 6155 125754 6158
rect 125636 6116 125662 6119
rect 125636 6087 125662 6090
rect 124532 6082 124558 6085
rect 124532 6053 124558 6056
rect 124624 6082 124650 6085
rect 124624 6053 124650 6056
rect 122416 5912 122442 5915
rect 122416 5883 122442 5886
rect 121358 5844 121384 5847
rect 121358 5815 121384 5818
rect 122278 5844 122304 5847
rect 122278 5815 122304 5818
rect 121036 5674 121062 5677
rect 121036 5645 121062 5648
rect 121364 5609 121378 5815
rect 124538 5779 124552 6053
rect 124532 5776 124558 5779
rect 124532 5747 124558 5750
rect 121358 5606 121384 5609
rect 121358 5577 121384 5580
rect 120438 5572 120464 5575
rect 120438 5543 120464 5546
rect 120990 5572 121016 5575
rect 120990 5543 121016 5546
rect 102728 5538 102754 5541
rect 102728 5509 102754 5512
rect 115378 5538 115404 5541
rect 115378 5509 115404 5512
rect 114772 5454 114926 5458
rect 114772 5453 114775 5454
rect 114803 5453 114815 5454
rect 114843 5453 114855 5454
rect 114883 5453 114895 5454
rect 114923 5453 114926 5454
rect 114803 5427 114804 5453
rect 114894 5427 114895 5453
rect 114772 5426 114775 5427
rect 114803 5426 114815 5427
rect 114843 5426 114855 5427
rect 114883 5426 114895 5427
rect 114923 5426 114926 5427
rect 114772 5421 114926 5426
rect 102544 5402 102570 5405
rect 102544 5373 102570 5376
rect 102406 5334 102432 5337
rect 102406 5305 102432 5308
rect 101762 5232 101788 5235
rect 101762 5203 101788 5206
rect 114772 4910 114926 4914
rect 114772 4909 114775 4910
rect 114803 4909 114815 4910
rect 114843 4909 114855 4910
rect 114883 4909 114895 4910
rect 114923 4909 114926 4910
rect 114803 4883 114804 4909
rect 114894 4883 114895 4909
rect 114772 4882 114775 4883
rect 114803 4882 114815 4883
rect 114843 4882 114855 4883
rect 114883 4882 114895 4883
rect 114923 4882 114926 4883
rect 114772 4877 114926 4882
rect 97990 4756 98016 4759
rect 97990 4727 98016 4730
rect 97254 4722 97280 4725
rect 97254 4693 97280 4696
rect 95722 4638 95876 4642
rect 95722 4637 95725 4638
rect 95753 4637 95765 4638
rect 95793 4637 95805 4638
rect 95833 4637 95845 4638
rect 95873 4637 95876 4638
rect 95753 4611 95754 4637
rect 95844 4611 95845 4637
rect 95722 4610 95725 4611
rect 95753 4610 95765 4611
rect 95793 4610 95805 4611
rect 95833 4610 95845 4611
rect 95873 4610 95876 4611
rect 95722 4605 95876 4610
rect 114772 4366 114926 4370
rect 114772 4365 114775 4366
rect 114803 4365 114815 4366
rect 114843 4365 114855 4366
rect 114883 4365 114895 4366
rect 114923 4365 114926 4366
rect 114803 4339 114804 4365
rect 114894 4339 114895 4365
rect 114772 4338 114775 4339
rect 114803 4338 114815 4339
rect 114843 4338 114855 4339
rect 114883 4338 114895 4339
rect 114923 4338 114926 4339
rect 114772 4333 114926 4338
rect 93758 4178 93784 4181
rect 93758 4149 93784 4152
rect 95722 4094 95876 4098
rect 95722 4093 95725 4094
rect 95753 4093 95765 4094
rect 95793 4093 95805 4094
rect 95833 4093 95845 4094
rect 95873 4093 95876 4094
rect 95753 4067 95754 4093
rect 95844 4067 95845 4093
rect 95722 4066 95725 4067
rect 95753 4066 95765 4067
rect 95793 4066 95805 4067
rect 95833 4066 95845 4067
rect 95873 4066 95876 4067
rect 95722 4061 95876 4066
rect 76673 3822 76827 3826
rect 76673 3821 76676 3822
rect 76704 3821 76716 3822
rect 76744 3821 76756 3822
rect 76784 3821 76796 3822
rect 76824 3821 76827 3822
rect 76704 3795 76705 3821
rect 76795 3795 76796 3821
rect 76673 3794 76676 3795
rect 76704 3794 76716 3795
rect 76744 3794 76756 3795
rect 76784 3794 76796 3795
rect 76824 3794 76827 3795
rect 76673 3789 76827 3794
rect 114772 3822 114926 3826
rect 114772 3821 114775 3822
rect 114803 3821 114815 3822
rect 114843 3821 114855 3822
rect 114883 3821 114895 3822
rect 114923 3821 114926 3822
rect 114803 3795 114804 3821
rect 114894 3795 114895 3821
rect 114772 3794 114775 3795
rect 114803 3794 114815 3795
rect 114843 3794 114855 3795
rect 114883 3794 114895 3795
rect 114923 3794 114926 3795
rect 114772 3789 114926 3794
rect 95722 3550 95876 3554
rect 95722 3549 95725 3550
rect 95753 3549 95765 3550
rect 95793 3549 95805 3550
rect 95833 3549 95845 3550
rect 95873 3549 95876 3550
rect 95753 3523 95754 3549
rect 95844 3523 95845 3549
rect 95722 3522 95725 3523
rect 95753 3522 95765 3523
rect 95793 3522 95805 3523
rect 95833 3522 95845 3523
rect 95873 3522 95876 3523
rect 95722 3517 95876 3522
rect 76673 3278 76827 3282
rect 76673 3277 76676 3278
rect 76704 3277 76716 3278
rect 76744 3277 76756 3278
rect 76784 3277 76796 3278
rect 76824 3277 76827 3278
rect 76704 3251 76705 3277
rect 76795 3251 76796 3277
rect 76673 3250 76676 3251
rect 76704 3250 76716 3251
rect 76744 3250 76756 3251
rect 76784 3250 76796 3251
rect 76824 3250 76827 3251
rect 76673 3245 76827 3250
rect 114772 3278 114926 3282
rect 114772 3277 114775 3278
rect 114803 3277 114815 3278
rect 114843 3277 114855 3278
rect 114883 3277 114895 3278
rect 114923 3277 114926 3278
rect 114803 3251 114804 3277
rect 114894 3251 114895 3277
rect 114772 3250 114775 3251
rect 114803 3250 114815 3251
rect 114843 3250 114855 3251
rect 114883 3250 114895 3251
rect 114923 3250 114926 3251
rect 114772 3245 114926 3250
rect 124538 3127 124552 5747
rect 125780 5575 125794 6393
rect 125826 5813 125840 6427
rect 126050 6388 126076 6391
rect 126050 6359 126076 6362
rect 125912 6354 125938 6357
rect 125912 6325 125938 6328
rect 125918 6240 125932 6325
rect 125958 6320 125984 6323
rect 125957 6304 125958 6308
rect 126004 6320 126030 6323
rect 125984 6304 125985 6308
rect 126004 6291 126030 6294
rect 125957 6271 125985 6276
rect 125911 6236 125939 6240
rect 125911 6203 125939 6208
rect 125958 6218 125984 6221
rect 125958 6189 125984 6192
rect 125964 6119 125978 6189
rect 125958 6116 125984 6119
rect 125958 6087 125984 6090
rect 126010 5881 126024 6291
rect 126056 6187 126070 6359
rect 126194 6217 126208 6597
rect 126240 6459 126254 6699
rect 126510 6626 126536 6629
rect 126510 6597 126536 6600
rect 126234 6456 126260 6459
rect 126234 6427 126260 6430
rect 126516 6217 126530 6597
rect 126194 6203 126254 6217
rect 126050 6184 126076 6187
rect 126050 6155 126076 6158
rect 126004 5878 126030 5881
rect 126004 5849 126030 5852
rect 126056 5847 126070 6155
rect 126050 5844 126076 5847
rect 126050 5815 126076 5818
rect 125820 5810 125846 5813
rect 125820 5781 125846 5784
rect 126240 5677 126254 6203
rect 126470 6203 126530 6217
rect 126470 5949 126484 6203
rect 126556 6082 126582 6085
rect 126556 6053 126582 6056
rect 126464 5946 126490 5949
rect 126464 5917 126490 5920
rect 126372 5878 126398 5881
rect 126372 5849 126398 5852
rect 126510 5878 126536 5881
rect 126510 5849 126536 5852
rect 126234 5674 126260 5677
rect 126234 5645 126260 5648
rect 126378 5643 126392 5849
rect 126372 5640 126398 5643
rect 126372 5611 126398 5614
rect 125774 5572 125800 5575
rect 125774 5543 125800 5546
rect 126378 4997 126392 5611
rect 126516 5575 126530 5849
rect 126562 5677 126576 6053
rect 126556 5674 126582 5677
rect 126556 5645 126582 5648
rect 126608 5643 126622 7600
rect 127476 6728 127502 6731
rect 127344 6708 127476 6722
rect 126740 6592 126766 6595
rect 126740 6563 126766 6566
rect 126746 6382 126760 6563
rect 127344 6493 127358 6708
rect 127476 6699 127502 6702
rect 128126 6705 128140 7600
rect 129690 6841 129704 7600
rect 129690 6827 129750 6841
rect 129736 6731 129750 6827
rect 129730 6728 129756 6731
rect 128126 6691 128278 6705
rect 129730 6699 129756 6702
rect 128120 6660 128146 6663
rect 128120 6631 128146 6634
rect 127476 6626 127502 6629
rect 127476 6597 127502 6600
rect 127660 6626 127686 6629
rect 127660 6597 127686 6600
rect 127338 6490 127364 6493
rect 127338 6461 127364 6464
rect 126832 6388 126858 6391
rect 126746 6368 126832 6382
rect 126832 6359 126858 6362
rect 126970 6388 126996 6391
rect 126970 6359 126996 6362
rect 126976 6161 126990 6359
rect 127154 6184 127180 6187
rect 126976 6147 127036 6161
rect 127154 6155 127180 6158
rect 126648 5776 126674 5779
rect 126648 5747 126674 5750
rect 126602 5640 126628 5643
rect 126602 5611 126628 5614
rect 126654 5575 126668 5747
rect 127022 5677 127036 6147
rect 127160 5915 127174 6155
rect 127200 6048 127226 6051
rect 127200 6019 127226 6022
rect 127154 5912 127180 5915
rect 127154 5883 127180 5886
rect 127016 5674 127042 5677
rect 127016 5645 127042 5648
rect 127206 5575 127220 6019
rect 127344 5949 127358 6461
rect 127482 6217 127496 6597
rect 127666 6569 127680 6597
rect 127620 6555 127680 6569
rect 127568 6388 127594 6391
rect 127568 6359 127594 6362
rect 127522 6354 127548 6357
rect 127522 6325 127548 6328
rect 127390 6203 127496 6217
rect 127390 5949 127404 6203
rect 127528 6093 127542 6325
rect 127574 6119 127588 6359
rect 127620 6217 127634 6555
rect 128126 6493 128140 6631
rect 128166 6592 128192 6595
rect 128166 6563 128192 6566
rect 128120 6490 128146 6493
rect 128120 6461 128146 6464
rect 128172 6391 128186 6563
rect 128166 6388 128192 6391
rect 128166 6359 128192 6362
rect 128212 6388 128238 6391
rect 128212 6359 128238 6362
rect 127620 6203 127680 6217
rect 127614 6184 127640 6187
rect 127614 6155 127640 6158
rect 127482 6079 127542 6093
rect 127568 6116 127594 6119
rect 127568 6087 127594 6090
rect 127338 5946 127364 5949
rect 127338 5917 127364 5920
rect 127384 5946 127410 5949
rect 127384 5917 127410 5920
rect 127344 5575 127358 5917
rect 126510 5572 126536 5575
rect 126510 5543 126536 5546
rect 126648 5572 126674 5575
rect 126648 5543 126674 5546
rect 127200 5572 127226 5575
rect 127200 5543 127226 5546
rect 127338 5572 127364 5575
rect 127338 5543 127364 5546
rect 127482 5337 127496 6079
rect 127620 6051 127634 6155
rect 127522 6048 127548 6051
rect 127522 6019 127548 6022
rect 127614 6048 127640 6051
rect 127614 6019 127640 6022
rect 127528 5949 127542 6019
rect 127522 5946 127548 5949
rect 127522 5917 127548 5920
rect 127666 5838 127680 6203
rect 127798 6150 127824 6153
rect 127798 6121 127824 6124
rect 127804 5847 127818 6121
rect 128120 6116 128146 6119
rect 128120 6087 128146 6090
rect 128166 6116 128192 6119
rect 128166 6087 128192 6090
rect 128126 5881 128140 6087
rect 128172 6051 128186 6087
rect 128166 6048 128192 6051
rect 128166 6019 128192 6022
rect 128120 5878 128146 5881
rect 128120 5849 128146 5852
rect 128218 5847 128232 6359
rect 128264 6221 128278 6691
rect 128488 6626 128514 6629
rect 128488 6597 128514 6600
rect 130926 6626 130952 6629
rect 130926 6597 130952 6600
rect 128303 6508 128331 6512
rect 128303 6475 128331 6480
rect 128310 6425 128324 6475
rect 128304 6422 128330 6425
rect 128304 6393 128330 6396
rect 128258 6218 128284 6221
rect 128258 6189 128284 6192
rect 128494 6187 128508 6597
rect 128994 6592 129020 6595
rect 128994 6563 129020 6566
rect 129000 6512 129014 6563
rect 128993 6508 129021 6512
rect 128993 6475 129021 6480
rect 128626 6456 128652 6459
rect 128626 6427 128652 6430
rect 130880 6456 130906 6459
rect 130880 6427 130906 6430
rect 128580 6388 128606 6391
rect 128580 6359 128606 6362
rect 128534 6354 128560 6357
rect 128534 6325 128560 6328
rect 128540 6308 128554 6325
rect 128533 6304 128561 6308
rect 128533 6271 128561 6276
rect 128586 6240 128600 6359
rect 128579 6236 128607 6240
rect 128579 6203 128607 6208
rect 128488 6184 128514 6187
rect 128488 6155 128514 6158
rect 128632 5881 128646 6427
rect 128626 5878 128652 5881
rect 128626 5849 128652 5852
rect 127620 5824 127680 5838
rect 127798 5844 127824 5847
rect 127620 5405 127634 5824
rect 127798 5815 127824 5818
rect 128212 5844 128238 5847
rect 128212 5815 128238 5818
rect 130886 5779 130900 6427
rect 130932 6425 130946 6597
rect 130926 6422 130952 6425
rect 130926 6393 130952 6396
rect 130932 6153 130946 6393
rect 131156 6388 131182 6391
rect 131155 6372 131156 6376
rect 131182 6372 131183 6376
rect 131155 6339 131183 6344
rect 131110 6320 131136 6323
rect 131136 6300 131222 6314
rect 131110 6291 131136 6294
rect 131208 6153 131222 6300
rect 131254 6221 131268 7643
rect 132719 7600 132747 8000
rect 134283 7600 134311 8000
rect 135801 7657 135829 8000
rect 137319 7657 137347 8000
rect 138883 7657 138911 8000
rect 140401 7657 140429 8000
rect 141965 7657 141993 8000
rect 135801 7643 135914 7657
rect 135801 7600 135829 7643
rect 131754 6728 131780 6731
rect 131754 6699 131780 6702
rect 131707 6644 131735 6648
rect 131760 6629 131774 6699
rect 132076 6694 132102 6697
rect 132076 6665 132102 6668
rect 131707 6611 131708 6616
rect 131734 6611 131735 6616
rect 131754 6626 131780 6629
rect 131708 6597 131734 6600
rect 131754 6597 131780 6600
rect 131478 6592 131504 6595
rect 131662 6592 131688 6595
rect 131504 6572 131544 6586
rect 131478 6563 131504 6566
rect 131340 6354 131366 6357
rect 131340 6325 131366 6328
rect 131248 6218 131274 6221
rect 131248 6189 131274 6192
rect 130926 6150 130952 6153
rect 130926 6121 130952 6124
rect 131202 6150 131228 6153
rect 131202 6121 131228 6124
rect 131346 5779 131360 6325
rect 131530 6119 131544 6572
rect 131662 6563 131688 6566
rect 131668 6459 131682 6563
rect 131662 6456 131688 6459
rect 131662 6427 131688 6430
rect 131753 6372 131781 6376
rect 131753 6339 131754 6344
rect 131780 6339 131781 6344
rect 131754 6325 131780 6328
rect 131984 6320 132010 6323
rect 131984 6291 132010 6294
rect 131524 6116 131550 6119
rect 131524 6087 131550 6090
rect 131990 5847 132004 6291
rect 132082 6153 132096 6665
rect 132214 6626 132240 6629
rect 132214 6597 132240 6600
rect 132306 6626 132332 6629
rect 132306 6597 132332 6600
rect 132490 6626 132516 6629
rect 132490 6597 132516 6600
rect 132220 6425 132234 6597
rect 132312 6493 132326 6597
rect 132306 6490 132332 6493
rect 132306 6461 132332 6464
rect 132168 6422 132194 6425
rect 132168 6393 132194 6396
rect 132214 6422 132240 6425
rect 132214 6393 132240 6396
rect 132174 6376 132188 6393
rect 132167 6372 132195 6376
rect 132167 6339 132195 6344
rect 132496 6187 132510 6597
rect 132490 6184 132516 6187
rect 132490 6155 132516 6158
rect 132076 6150 132102 6153
rect 132076 6121 132102 6124
rect 132582 6150 132608 6153
rect 132582 6121 132608 6124
rect 132168 6116 132194 6119
rect 132168 6087 132194 6090
rect 132174 5881 132188 6087
rect 132588 6085 132602 6121
rect 132582 6082 132608 6085
rect 132582 6053 132608 6056
rect 132588 5957 132602 6053
rect 132588 5943 132648 5957
rect 132634 5881 132648 5943
rect 132168 5878 132194 5881
rect 132168 5849 132194 5852
rect 132582 5878 132608 5881
rect 132582 5849 132608 5852
rect 132628 5878 132654 5881
rect 132628 5849 132654 5852
rect 131984 5844 132010 5847
rect 131984 5815 132010 5818
rect 130880 5776 130906 5779
rect 130880 5747 130906 5750
rect 131340 5776 131366 5779
rect 131340 5747 131366 5750
rect 132174 5575 132188 5849
rect 132588 5643 132602 5849
rect 132726 5677 132740 7600
rect 133821 6814 133975 6818
rect 133821 6813 133824 6814
rect 133852 6813 133864 6814
rect 133892 6813 133904 6814
rect 133932 6813 133944 6814
rect 133972 6813 133975 6814
rect 133852 6787 133853 6813
rect 133943 6787 133944 6813
rect 133821 6786 133824 6787
rect 133852 6786 133864 6787
rect 133892 6786 133904 6787
rect 133932 6786 133944 6787
rect 133972 6786 133975 6787
rect 133821 6781 133975 6786
rect 132766 6728 132792 6731
rect 132766 6699 132792 6702
rect 132772 6648 132786 6699
rect 132765 6644 132793 6648
rect 132793 6623 132832 6637
rect 132765 6611 132793 6616
rect 132766 6456 132792 6459
rect 132766 6427 132792 6430
rect 132772 6221 132786 6427
rect 132766 6218 132792 6221
rect 132766 6189 132792 6192
rect 132818 6153 132832 6623
rect 133456 6626 133482 6629
rect 133456 6597 133482 6600
rect 133272 6456 133298 6459
rect 133272 6427 133298 6430
rect 132812 6150 132838 6153
rect 132812 6121 132838 6124
rect 132720 5674 132746 5677
rect 132720 5645 132746 5648
rect 132582 5640 132608 5643
rect 132582 5611 132608 5614
rect 132818 5575 132832 6121
rect 133134 5776 133160 5779
rect 133134 5747 133160 5750
rect 133180 5776 133206 5779
rect 133180 5747 133206 5750
rect 133140 5677 133154 5747
rect 133134 5674 133160 5677
rect 133134 5645 133160 5648
rect 132168 5572 132194 5575
rect 132168 5543 132194 5546
rect 132444 5572 132470 5575
rect 132444 5543 132470 5546
rect 132812 5572 132838 5575
rect 132812 5543 132838 5546
rect 127614 5402 127640 5405
rect 127614 5373 127640 5376
rect 132450 5371 132464 5543
rect 132444 5368 132470 5371
rect 132444 5339 132470 5342
rect 133186 5337 133200 5747
rect 133278 5405 133292 6427
rect 133410 6082 133436 6085
rect 133410 6053 133436 6056
rect 133416 5949 133430 6053
rect 133410 5946 133436 5949
rect 133410 5917 133436 5920
rect 133272 5402 133298 5405
rect 133272 5373 133298 5376
rect 127476 5334 127502 5337
rect 127476 5305 127502 5308
rect 133180 5334 133206 5337
rect 133180 5305 133206 5308
rect 133462 5133 133476 6597
rect 133824 6592 133850 6595
rect 133824 6563 133850 6566
rect 133502 6388 133528 6391
rect 133778 6388 133804 6391
rect 133502 6359 133528 6362
rect 133547 6372 133575 6376
rect 133508 6323 133522 6359
rect 133830 6376 133844 6563
rect 134192 6490 134218 6493
rect 134192 6461 134218 6464
rect 134146 6422 134172 6425
rect 134146 6393 134172 6396
rect 134008 6388 134034 6391
rect 133778 6359 133804 6362
rect 133823 6372 133851 6376
rect 133547 6339 133575 6344
rect 133554 6323 133568 6339
rect 133784 6323 133798 6359
rect 134008 6359 134034 6362
rect 134053 6372 134081 6376
rect 133823 6339 133851 6344
rect 133502 6320 133528 6323
rect 133502 6291 133528 6294
rect 133548 6320 133574 6323
rect 133548 6291 133574 6294
rect 133778 6320 133804 6323
rect 133778 6291 133804 6294
rect 133508 6051 133522 6291
rect 133821 6270 133975 6274
rect 133821 6269 133824 6270
rect 133852 6269 133864 6270
rect 133892 6269 133904 6270
rect 133932 6269 133944 6270
rect 133972 6269 133975 6270
rect 133852 6243 133853 6269
rect 133943 6243 133944 6269
rect 133821 6242 133824 6243
rect 133852 6242 133864 6243
rect 133892 6242 133904 6243
rect 133932 6242 133944 6243
rect 133972 6242 133975 6243
rect 133821 6237 133975 6242
rect 134014 6221 134028 6359
rect 134053 6339 134081 6344
rect 134008 6218 134034 6221
rect 134008 6189 134034 6192
rect 133640 6082 133666 6085
rect 133640 6053 133666 6056
rect 133502 6048 133528 6051
rect 133502 6019 133528 6022
rect 133646 5609 133660 6053
rect 134014 5813 134028 6189
rect 134060 6119 134074 6339
rect 134054 6116 134080 6119
rect 134054 6087 134080 6090
rect 134008 5810 134034 5813
rect 134008 5781 134034 5784
rect 133821 5726 133975 5730
rect 133821 5725 133824 5726
rect 133852 5725 133864 5726
rect 133892 5725 133904 5726
rect 133932 5725 133944 5726
rect 133972 5725 133975 5726
rect 133852 5699 133853 5725
rect 133943 5699 133944 5725
rect 133821 5698 133824 5699
rect 133852 5698 133864 5699
rect 133892 5698 133904 5699
rect 133932 5698 133944 5699
rect 133972 5698 133975 5699
rect 133821 5693 133975 5698
rect 134014 5609 134028 5781
rect 133640 5606 133666 5609
rect 133640 5577 133666 5580
rect 134008 5606 134034 5609
rect 134008 5577 134034 5580
rect 133821 5182 133975 5186
rect 133821 5181 133824 5182
rect 133852 5181 133864 5182
rect 133892 5181 133904 5182
rect 133932 5181 133944 5182
rect 133972 5181 133975 5182
rect 133852 5155 133853 5181
rect 133943 5155 133944 5181
rect 133821 5154 133824 5155
rect 133852 5154 133864 5155
rect 133892 5154 133904 5155
rect 133932 5154 133944 5155
rect 133972 5154 133975 5155
rect 133821 5149 133975 5154
rect 133456 5130 133482 5133
rect 133456 5101 133482 5104
rect 133870 5062 133896 5065
rect 133870 5033 133896 5036
rect 126372 4994 126398 4997
rect 126372 4965 126398 4968
rect 133876 4963 133890 5033
rect 134060 5031 134074 6087
rect 134100 6082 134126 6085
rect 134100 6053 134126 6056
rect 134106 5405 134120 6053
rect 134152 5915 134166 6393
rect 134198 6391 134212 6461
rect 134192 6388 134218 6391
rect 134192 6359 134218 6362
rect 134192 6218 134218 6221
rect 134192 6189 134218 6192
rect 134146 5912 134172 5915
rect 134146 5883 134172 5886
rect 134152 5541 134166 5883
rect 134146 5538 134172 5541
rect 134146 5509 134172 5512
rect 134100 5402 134126 5405
rect 134100 5373 134126 5376
rect 134198 5099 134212 6189
rect 134238 6048 134264 6051
rect 134238 6019 134264 6022
rect 134244 5881 134258 6019
rect 134238 5878 134264 5881
rect 134238 5849 134264 5852
rect 134244 5609 134258 5849
rect 134238 5606 134264 5609
rect 134238 5577 134264 5580
rect 134290 5133 134304 7600
rect 135900 6765 135914 7643
rect 137319 7643 137478 7657
rect 137319 7600 137347 7643
rect 137464 6765 137478 7643
rect 138883 7643 138950 7657
rect 138883 7600 138911 7643
rect 138936 6765 138950 7643
rect 140401 7643 140468 7657
rect 140401 7600 140429 7643
rect 140454 6765 140468 7643
rect 141965 7643 142124 7657
rect 141965 7600 141993 7643
rect 134468 6762 134494 6765
rect 134468 6733 134494 6736
rect 134790 6762 134816 6765
rect 134790 6733 134816 6736
rect 135894 6762 135920 6765
rect 135894 6733 135920 6736
rect 137458 6762 137484 6765
rect 137458 6733 137484 6736
rect 138930 6762 138956 6765
rect 138930 6733 138956 6736
rect 140448 6762 140474 6765
rect 142110 6756 142124 7643
rect 143483 7600 143511 8000
rect 145001 7657 145029 8000
rect 146565 7657 146593 8000
rect 148083 7657 148111 8000
rect 149601 7657 149629 8000
rect 151165 7657 151193 8000
rect 145001 7643 145068 7657
rect 145001 7600 145029 7643
rect 142150 6762 142176 6765
rect 142110 6742 142150 6756
rect 140448 6733 140474 6736
rect 143490 6756 143504 7600
rect 145054 6765 145068 7643
rect 146565 7643 146632 7657
rect 146565 7600 146593 7643
rect 146618 6765 146632 7643
rect 148083 7643 148150 7657
rect 148083 7600 148111 7643
rect 148136 6765 148150 7643
rect 149601 7643 149668 7657
rect 149601 7600 149629 7643
rect 149654 6765 149668 7643
rect 151165 7643 151324 7657
rect 151165 7600 151193 7643
rect 150706 6864 150732 6867
rect 150706 6835 150732 6838
rect 150712 6765 150726 6835
rect 143530 6762 143556 6765
rect 143490 6742 143530 6756
rect 142150 6733 142176 6736
rect 143530 6733 143556 6736
rect 145048 6762 145074 6765
rect 145048 6733 145074 6736
rect 146612 6762 146638 6765
rect 146612 6733 146638 6736
rect 148130 6762 148156 6765
rect 148130 6733 148156 6736
rect 149648 6762 149674 6765
rect 149648 6733 149674 6736
rect 150706 6762 150732 6765
rect 150706 6733 150732 6736
rect 134474 6716 134488 6733
rect 134467 6712 134495 6716
rect 134467 6679 134495 6684
rect 134474 6663 134488 6679
rect 134468 6660 134494 6663
rect 134468 6631 134494 6634
rect 134513 6644 134541 6648
rect 134376 6626 134402 6629
rect 134376 6597 134402 6600
rect 134330 6116 134356 6119
rect 134330 6087 134356 6090
rect 134336 6051 134350 6087
rect 134330 6048 134356 6051
rect 134330 6019 134356 6022
rect 134382 5269 134396 6597
rect 134474 5609 134488 6631
rect 134513 6611 134541 6616
rect 134520 6425 134534 6611
rect 134514 6422 134540 6425
rect 134514 6393 134540 6396
rect 134698 6388 134724 6391
rect 134658 6368 134698 6382
rect 134560 6320 134586 6323
rect 134586 6300 134626 6314
rect 134560 6291 134586 6294
rect 134560 6150 134586 6153
rect 134560 6121 134586 6124
rect 134566 5881 134580 6121
rect 134560 5878 134586 5881
rect 134560 5849 134586 5852
rect 134468 5606 134494 5609
rect 134468 5577 134494 5580
rect 134474 5541 134488 5577
rect 134468 5538 134494 5541
rect 134468 5509 134494 5512
rect 134422 5504 134448 5507
rect 134422 5475 134448 5478
rect 134376 5266 134402 5269
rect 134376 5237 134402 5240
rect 134284 5130 134310 5133
rect 134284 5101 134310 5104
rect 134192 5096 134218 5099
rect 134192 5067 134218 5070
rect 134428 5065 134442 5475
rect 134514 5334 134540 5337
rect 134514 5305 134540 5308
rect 134422 5062 134448 5065
rect 134422 5033 134448 5036
rect 134520 5031 134534 5305
rect 134612 5031 134626 6300
rect 134658 5677 134672 6368
rect 134698 6359 134724 6362
rect 134744 6082 134770 6085
rect 134744 6053 134770 6056
rect 134698 5844 134724 5847
rect 134698 5815 134724 5818
rect 134652 5674 134678 5677
rect 134652 5645 134678 5648
rect 134704 5405 134718 5815
rect 134698 5402 134724 5405
rect 134698 5373 134724 5376
rect 134750 5099 134764 6053
rect 134796 5235 134810 6733
rect 135204 6728 135230 6731
rect 136492 6728 136518 6731
rect 135204 6699 135230 6702
rect 136406 6702 136492 6705
rect 136406 6699 136518 6702
rect 136583 6712 136611 6716
rect 134836 6150 134862 6153
rect 134836 6121 134862 6124
rect 134842 5575 134856 6121
rect 135210 6093 135224 6699
rect 136406 6691 136512 6699
rect 135342 6626 135368 6629
rect 135342 6597 135368 6600
rect 135480 6626 135506 6629
rect 135480 6597 135506 6600
rect 135164 6079 135224 6093
rect 134928 5912 134954 5915
rect 134928 5883 134954 5886
rect 134836 5572 134862 5575
rect 134836 5543 134862 5546
rect 134790 5232 134816 5235
rect 134790 5203 134816 5206
rect 134744 5096 134770 5099
rect 134744 5067 134770 5070
rect 134054 5028 134080 5031
rect 134054 4999 134080 5002
rect 134514 5028 134540 5031
rect 134514 4999 134540 5002
rect 134606 5028 134632 5031
rect 134606 4999 134632 5002
rect 133870 4960 133896 4963
rect 133870 4931 133896 4934
rect 134060 4793 134074 4999
rect 134934 4827 134948 5883
rect 134974 5844 135000 5847
rect 134974 5815 135000 5818
rect 134980 5541 134994 5815
rect 134974 5538 135000 5541
rect 134974 5509 135000 5512
rect 135020 5504 135046 5507
rect 135020 5475 135046 5478
rect 135026 5371 135040 5475
rect 135020 5368 135046 5371
rect 135020 5339 135046 5342
rect 135164 5337 135178 6079
rect 135204 6048 135230 6051
rect 135204 6019 135230 6022
rect 135210 5575 135224 6019
rect 135348 5949 135362 6597
rect 135388 6592 135414 6595
rect 135388 6563 135414 6566
rect 135394 5949 135408 6563
rect 135434 6422 135460 6425
rect 135434 6393 135460 6396
rect 135440 6323 135454 6393
rect 135434 6320 135460 6323
rect 135434 6291 135460 6294
rect 135342 5946 135368 5949
rect 135342 5917 135368 5920
rect 135388 5946 135414 5949
rect 135388 5917 135414 5920
rect 135440 5575 135454 6291
rect 135204 5572 135230 5575
rect 135204 5543 135230 5546
rect 135434 5572 135460 5575
rect 135434 5543 135460 5546
rect 135158 5334 135184 5337
rect 135158 5305 135184 5308
rect 135486 4963 135500 6597
rect 135894 6592 135920 6595
rect 135894 6563 135920 6566
rect 135900 6459 135914 6563
rect 136406 6459 136420 6691
rect 136583 6679 136584 6684
rect 136610 6679 136611 6684
rect 136584 6665 136610 6668
rect 136630 6660 136656 6663
rect 136629 6644 136630 6648
rect 137550 6660 137576 6663
rect 136656 6644 136657 6648
rect 137550 6631 137576 6634
rect 140540 6660 140566 6663
rect 140540 6631 140566 6634
rect 142380 6660 142406 6663
rect 142380 6631 142406 6634
rect 145140 6660 145166 6663
rect 145140 6631 145166 6634
rect 149740 6660 149766 6663
rect 149740 6631 149766 6634
rect 136629 6611 136657 6616
rect 136446 6592 136472 6595
rect 136446 6563 136472 6566
rect 135526 6456 135552 6459
rect 135526 6427 135552 6430
rect 135894 6456 135920 6459
rect 135894 6427 135920 6430
rect 136400 6456 136426 6459
rect 136400 6427 136426 6430
rect 135532 6221 135546 6427
rect 136308 6422 136334 6425
rect 136308 6393 136334 6396
rect 136124 6388 136150 6391
rect 136124 6359 136150 6362
rect 135572 6320 135598 6323
rect 135572 6291 135598 6294
rect 135526 6218 135552 6221
rect 135526 6189 135552 6192
rect 135578 6153 135592 6291
rect 136130 6153 136144 6359
rect 136314 6323 136328 6393
rect 136452 6391 136466 6563
rect 136584 6456 136610 6459
rect 136584 6427 136610 6430
rect 136590 6391 136604 6427
rect 136446 6388 136472 6391
rect 136446 6359 136472 6362
rect 136584 6388 136610 6391
rect 136584 6359 136610 6362
rect 136400 6354 136426 6357
rect 136400 6325 136426 6328
rect 136262 6320 136288 6323
rect 136262 6291 136288 6294
rect 136308 6320 136334 6323
rect 136308 6291 136334 6294
rect 135572 6150 135598 6153
rect 135572 6121 135598 6124
rect 136124 6150 136150 6153
rect 136124 6121 136150 6124
rect 135664 6116 135690 6119
rect 135664 6087 135690 6090
rect 135670 5881 135684 6087
rect 135664 5878 135690 5881
rect 135664 5849 135690 5852
rect 136130 5609 136144 6121
rect 136124 5606 136150 5609
rect 136124 5577 136150 5580
rect 136268 5303 136282 6291
rect 136406 6153 136420 6325
rect 136400 6150 136426 6153
rect 136400 6121 136426 6124
rect 136452 6119 136466 6359
rect 136446 6116 136472 6119
rect 136446 6087 136472 6090
rect 136590 5847 136604 6359
rect 136584 5844 136610 5847
rect 136584 5815 136610 5818
rect 137556 5779 137570 6631
rect 140546 6323 140560 6631
rect 140540 6320 140566 6323
rect 140540 6291 140566 6294
rect 142386 6051 142400 6631
rect 145146 6425 145160 6631
rect 147946 6592 147972 6595
rect 147946 6563 147972 6566
rect 147952 6459 147966 6563
rect 147946 6456 147972 6459
rect 149746 6444 149760 6631
rect 151310 6493 151324 7643
rect 152683 7600 152711 8000
rect 151763 6984 151791 6988
rect 151763 6951 151791 6956
rect 151396 6898 151422 6901
rect 151396 6869 151422 6872
rect 151304 6490 151330 6493
rect 151304 6461 151330 6464
rect 147946 6427 147972 6430
rect 149739 6440 149767 6444
rect 145140 6422 145166 6425
rect 151402 6425 151416 6869
rect 151770 6663 151784 6951
rect 152500 6694 152526 6697
rect 152500 6665 152526 6668
rect 151764 6660 151790 6663
rect 151764 6631 151790 6634
rect 152506 6459 152520 6665
rect 152690 6493 152704 7600
rect 152684 6490 152710 6493
rect 152684 6461 152710 6464
rect 152500 6456 152526 6459
rect 152500 6427 152526 6430
rect 152730 6456 152756 6459
rect 152730 6427 152756 6430
rect 149739 6407 149767 6412
rect 151396 6422 151422 6425
rect 145140 6393 145166 6396
rect 151396 6393 151422 6396
rect 152736 6221 152750 6427
rect 152730 6218 152756 6221
rect 152730 6189 152756 6192
rect 142380 6048 142406 6051
rect 142380 6019 142406 6022
rect 137550 5776 137576 5779
rect 137550 5747 137576 5750
rect 136262 5300 136288 5303
rect 136262 5271 136288 5274
rect 152224 5028 152250 5031
rect 152223 5012 152224 5016
rect 152250 5012 152251 5016
rect 152223 4979 152251 4984
rect 135480 4960 135506 4963
rect 135480 4931 135506 4934
rect 134928 4824 134954 4827
rect 134928 4795 134954 4798
rect 134054 4790 134080 4793
rect 134054 4761 134080 4764
rect 133821 4638 133975 4642
rect 133821 4637 133824 4638
rect 133852 4637 133864 4638
rect 133892 4637 133904 4638
rect 133932 4637 133944 4638
rect 133972 4637 133975 4638
rect 133852 4611 133853 4637
rect 133943 4611 133944 4637
rect 133821 4610 133824 4611
rect 133852 4610 133864 4611
rect 133892 4610 133904 4611
rect 133932 4610 133944 4611
rect 133972 4610 133975 4611
rect 133821 4605 133975 4610
rect 133821 4094 133975 4098
rect 133821 4093 133824 4094
rect 133852 4093 133864 4094
rect 133892 4093 133904 4094
rect 133932 4093 133944 4094
rect 133972 4093 133975 4094
rect 133852 4067 133853 4093
rect 133943 4067 133944 4093
rect 133821 4066 133824 4067
rect 133852 4066 133864 4067
rect 133892 4066 133904 4067
rect 133932 4066 133944 4067
rect 133972 4066 133975 4067
rect 133821 4061 133975 4066
rect 133821 3550 133975 3554
rect 133821 3549 133824 3550
rect 133852 3549 133864 3550
rect 133892 3549 133904 3550
rect 133932 3549 133944 3550
rect 133972 3549 133975 3550
rect 133852 3523 133853 3549
rect 133943 3523 133944 3549
rect 133821 3522 133824 3523
rect 133852 3522 133864 3523
rect 133892 3522 133904 3523
rect 133932 3522 133944 3523
rect 133972 3522 133975 3523
rect 133821 3517 133975 3522
rect 151994 3158 152020 3161
rect 151994 3129 152020 3132
rect 124532 3124 124558 3127
rect 124532 3095 124558 3098
rect 95722 3006 95876 3010
rect 95722 3005 95725 3006
rect 95753 3005 95765 3006
rect 95793 3005 95805 3006
rect 95833 3005 95845 3006
rect 95873 3005 95876 3006
rect 95753 2979 95754 3005
rect 95844 2979 95845 3005
rect 95722 2978 95725 2979
rect 95753 2978 95765 2979
rect 95793 2978 95805 2979
rect 95833 2978 95845 2979
rect 95873 2978 95876 2979
rect 95722 2973 95876 2978
rect 133821 3006 133975 3010
rect 133821 3005 133824 3006
rect 133852 3005 133864 3006
rect 133892 3005 133904 3006
rect 133932 3005 133944 3006
rect 133972 3005 133975 3006
rect 133852 2979 133853 3005
rect 133943 2979 133944 3005
rect 133821 2978 133824 2979
rect 133852 2978 133864 2979
rect 133892 2978 133904 2979
rect 133932 2978 133944 2979
rect 133972 2978 133975 2979
rect 133821 2973 133975 2978
rect 152000 2976 152014 3129
rect 151993 2972 152021 2976
rect 151993 2939 152021 2944
rect 76673 2734 76827 2738
rect 76673 2733 76676 2734
rect 76704 2733 76716 2734
rect 76744 2733 76756 2734
rect 76784 2733 76796 2734
rect 76824 2733 76827 2734
rect 76704 2707 76705 2733
rect 76795 2707 76796 2733
rect 76673 2706 76676 2707
rect 76704 2706 76716 2707
rect 76744 2706 76756 2707
rect 76784 2706 76796 2707
rect 76824 2706 76827 2707
rect 76673 2701 76827 2706
rect 114772 2734 114926 2738
rect 114772 2733 114775 2734
rect 114803 2733 114815 2734
rect 114843 2733 114855 2734
rect 114883 2733 114895 2734
rect 114923 2733 114926 2734
rect 114803 2707 114804 2733
rect 114894 2707 114895 2733
rect 114772 2706 114775 2707
rect 114803 2706 114815 2707
rect 114843 2706 114855 2707
rect 114883 2706 114895 2707
rect 114923 2706 114926 2707
rect 114772 2701 114926 2706
rect 95722 2462 95876 2466
rect 95722 2461 95725 2462
rect 95753 2461 95765 2462
rect 95793 2461 95805 2462
rect 95833 2461 95845 2462
rect 95873 2461 95876 2462
rect 95753 2435 95754 2461
rect 95844 2435 95845 2461
rect 95722 2434 95725 2435
rect 95753 2434 95765 2435
rect 95793 2434 95805 2435
rect 95833 2434 95845 2435
rect 95873 2434 95876 2435
rect 95722 2429 95876 2434
rect 133821 2462 133975 2466
rect 133821 2461 133824 2462
rect 133852 2461 133864 2462
rect 133892 2461 133904 2462
rect 133932 2461 133944 2462
rect 133972 2461 133975 2462
rect 133852 2435 133853 2461
rect 133943 2435 133944 2461
rect 133821 2434 133824 2435
rect 133852 2434 133864 2435
rect 133892 2434 133904 2435
rect 133932 2434 133944 2435
rect 133972 2434 133975 2435
rect 133821 2429 133975 2434
rect 76673 2190 76827 2194
rect 76673 2189 76676 2190
rect 76704 2189 76716 2190
rect 76744 2189 76756 2190
rect 76784 2189 76796 2190
rect 76824 2189 76827 2190
rect 76704 2163 76705 2189
rect 76795 2163 76796 2189
rect 76673 2162 76676 2163
rect 76704 2162 76716 2163
rect 76744 2162 76756 2163
rect 76784 2162 76796 2163
rect 76824 2162 76827 2163
rect 76673 2157 76827 2162
rect 114772 2190 114926 2194
rect 114772 2189 114775 2190
rect 114803 2189 114815 2190
rect 114843 2189 114855 2190
rect 114883 2189 114895 2190
rect 114923 2189 114926 2190
rect 114803 2163 114804 2189
rect 114894 2163 114895 2189
rect 114772 2162 114775 2163
rect 114803 2162 114815 2163
rect 114843 2162 114855 2163
rect 114883 2162 114895 2163
rect 114923 2162 114926 2163
rect 114772 2157 114926 2162
rect 95722 1918 95876 1922
rect 95722 1917 95725 1918
rect 95753 1917 95765 1918
rect 95793 1917 95805 1918
rect 95833 1917 95845 1918
rect 95873 1917 95876 1918
rect 95753 1891 95754 1917
rect 95844 1891 95845 1917
rect 95722 1890 95725 1891
rect 95753 1890 95765 1891
rect 95793 1890 95805 1891
rect 95833 1890 95845 1891
rect 95873 1890 95876 1891
rect 95722 1885 95876 1890
rect 133821 1918 133975 1922
rect 133821 1917 133824 1918
rect 133852 1917 133864 1918
rect 133892 1917 133904 1918
rect 133932 1917 133944 1918
rect 133972 1917 133975 1918
rect 133852 1891 133853 1917
rect 133943 1891 133944 1917
rect 133821 1890 133824 1891
rect 133852 1890 133864 1891
rect 133892 1890 133904 1891
rect 133932 1890 133944 1891
rect 133972 1890 133975 1891
rect 133821 1885 133975 1890
rect 76673 1646 76827 1650
rect 76673 1645 76676 1646
rect 76704 1645 76716 1646
rect 76744 1645 76756 1646
rect 76784 1645 76796 1646
rect 76824 1645 76827 1646
rect 76704 1619 76705 1645
rect 76795 1619 76796 1645
rect 76673 1618 76676 1619
rect 76704 1618 76716 1619
rect 76744 1618 76756 1619
rect 76784 1618 76796 1619
rect 76824 1618 76827 1619
rect 76673 1613 76827 1618
rect 114772 1646 114926 1650
rect 114772 1645 114775 1646
rect 114803 1645 114815 1646
rect 114843 1645 114855 1646
rect 114883 1645 114895 1646
rect 114923 1645 114926 1646
rect 114803 1619 114804 1645
rect 114894 1619 114895 1645
rect 114772 1618 114775 1619
rect 114803 1618 114815 1619
rect 114843 1618 114855 1619
rect 114883 1618 114895 1619
rect 114923 1618 114926 1619
rect 114772 1613 114926 1618
rect 95722 1374 95876 1378
rect 95722 1373 95725 1374
rect 95753 1373 95765 1374
rect 95793 1373 95805 1374
rect 95833 1373 95845 1374
rect 95873 1373 95876 1374
rect 95753 1347 95754 1373
rect 95844 1347 95845 1373
rect 95722 1346 95725 1347
rect 95753 1346 95765 1347
rect 95793 1346 95805 1347
rect 95833 1346 95845 1347
rect 95873 1346 95876 1347
rect 95722 1341 95876 1346
rect 133821 1374 133975 1378
rect 133821 1373 133824 1374
rect 133852 1373 133864 1374
rect 133892 1373 133904 1374
rect 133932 1373 133944 1374
rect 133972 1373 133975 1374
rect 133852 1347 133853 1373
rect 133943 1347 133944 1373
rect 133821 1346 133824 1347
rect 133852 1346 133864 1347
rect 133892 1346 133904 1347
rect 133932 1346 133944 1347
rect 133972 1346 133975 1347
rect 133821 1341 133975 1346
rect 74714 1322 74740 1325
rect 74714 1293 74740 1296
rect 151120 1322 151146 1325
rect 151120 1293 151146 1296
rect 38574 1102 38728 1106
rect 38574 1101 38577 1102
rect 38605 1101 38617 1102
rect 38645 1101 38657 1102
rect 38685 1101 38697 1102
rect 38725 1101 38728 1102
rect 38605 1075 38606 1101
rect 38696 1075 38697 1101
rect 38574 1074 38577 1075
rect 38605 1074 38617 1075
rect 38645 1074 38657 1075
rect 38685 1074 38697 1075
rect 38725 1074 38728 1075
rect 38574 1069 38728 1074
rect 76673 1102 76827 1106
rect 76673 1101 76676 1102
rect 76704 1101 76716 1102
rect 76744 1101 76756 1102
rect 76784 1101 76796 1102
rect 76824 1101 76827 1102
rect 76704 1075 76705 1101
rect 76795 1075 76796 1101
rect 76673 1074 76676 1075
rect 76704 1074 76716 1075
rect 76744 1074 76756 1075
rect 76784 1074 76796 1075
rect 76824 1074 76827 1075
rect 76673 1069 76827 1074
rect 114772 1102 114926 1106
rect 114772 1101 114775 1102
rect 114803 1101 114815 1102
rect 114843 1101 114855 1102
rect 114883 1101 114895 1102
rect 114923 1101 114926 1102
rect 114803 1075 114804 1101
rect 114894 1075 114895 1101
rect 114772 1074 114775 1075
rect 114803 1074 114815 1075
rect 114843 1074 114855 1075
rect 114883 1074 114895 1075
rect 114923 1074 114926 1075
rect 114772 1069 114926 1074
rect 151126 1004 151140 1293
rect 151119 1000 151147 1004
rect 151119 967 151147 972
<< via2 >>
rect 14683 6090 14684 6100
rect 14684 6090 14710 6100
rect 14710 6090 14711 6100
rect 14683 6072 14711 6090
rect 15373 6072 15401 6100
rect 15695 6072 15723 6100
rect 19527 6813 19555 6814
rect 19567 6813 19595 6814
rect 19607 6813 19635 6814
rect 19647 6813 19675 6814
rect 19527 6787 19550 6813
rect 19550 6787 19555 6813
rect 19567 6787 19582 6813
rect 19582 6787 19588 6813
rect 19588 6787 19595 6813
rect 19607 6787 19614 6813
rect 19614 6787 19620 6813
rect 19620 6787 19635 6813
rect 19647 6787 19652 6813
rect 19652 6787 19675 6813
rect 19527 6786 19555 6787
rect 19567 6786 19595 6787
rect 19607 6786 19635 6787
rect 19647 6786 19675 6787
rect 19527 6269 19555 6270
rect 19567 6269 19595 6270
rect 19607 6269 19635 6270
rect 19647 6269 19675 6270
rect 19527 6243 19550 6269
rect 19550 6243 19555 6269
rect 19567 6243 19582 6269
rect 19582 6243 19588 6269
rect 19588 6243 19595 6269
rect 19607 6243 19614 6269
rect 19614 6243 19620 6269
rect 19620 6243 19635 6269
rect 19647 6243 19652 6269
rect 19652 6243 19675 6269
rect 19527 6242 19555 6243
rect 19567 6242 19595 6243
rect 19607 6242 19635 6243
rect 19647 6242 19675 6243
rect 19527 5725 19555 5726
rect 19567 5725 19595 5726
rect 19607 5725 19635 5726
rect 19647 5725 19675 5726
rect 19527 5699 19550 5725
rect 19550 5699 19555 5725
rect 19567 5699 19582 5725
rect 19582 5699 19588 5725
rect 19588 5699 19595 5725
rect 19607 5699 19614 5725
rect 19614 5699 19620 5725
rect 19620 5699 19635 5725
rect 19647 5699 19652 5725
rect 19652 5699 19675 5725
rect 19527 5698 19555 5699
rect 19567 5698 19595 5699
rect 19607 5698 19635 5699
rect 19647 5698 19675 5699
rect 20295 6090 20296 6100
rect 20296 6090 20322 6100
rect 20322 6090 20323 6100
rect 20295 6072 20323 6090
rect 21215 6072 21243 6100
rect 38577 6541 38605 6542
rect 38617 6541 38645 6542
rect 38657 6541 38685 6542
rect 38697 6541 38725 6542
rect 38577 6515 38600 6541
rect 38600 6515 38605 6541
rect 38617 6515 38632 6541
rect 38632 6515 38638 6541
rect 38638 6515 38645 6541
rect 38657 6515 38664 6541
rect 38664 6515 38670 6541
rect 38670 6515 38685 6541
rect 38697 6515 38702 6541
rect 38702 6515 38725 6541
rect 38577 6514 38605 6515
rect 38617 6514 38645 6515
rect 38657 6514 38685 6515
rect 38697 6514 38725 6515
rect 38577 5997 38605 5998
rect 38617 5997 38645 5998
rect 38657 5997 38685 5998
rect 38697 5997 38725 5998
rect 38577 5971 38600 5997
rect 38600 5971 38605 5997
rect 38617 5971 38632 5997
rect 38632 5971 38638 5997
rect 38638 5971 38645 5997
rect 38657 5971 38664 5997
rect 38664 5971 38670 5997
rect 38670 5971 38685 5997
rect 38697 5971 38702 5997
rect 38702 5971 38725 5997
rect 38577 5970 38605 5971
rect 38617 5970 38645 5971
rect 38657 5970 38685 5971
rect 38697 5970 38725 5971
rect 43479 6548 43507 6576
rect 43893 6344 43921 6372
rect 44077 6150 44105 6168
rect 44077 6140 44078 6150
rect 44078 6140 44104 6150
rect 44104 6140 44105 6150
rect 45917 6548 45945 6576
rect 44951 6140 44979 6168
rect 45365 6344 45393 6372
rect 38577 5453 38605 5454
rect 38617 5453 38645 5454
rect 38657 5453 38685 5454
rect 38697 5453 38725 5454
rect 38577 5427 38600 5453
rect 38600 5427 38605 5453
rect 38617 5427 38632 5453
rect 38632 5427 38638 5453
rect 38638 5427 38645 5453
rect 38657 5427 38664 5453
rect 38664 5427 38670 5453
rect 38670 5427 38685 5453
rect 38697 5427 38702 5453
rect 38702 5427 38725 5453
rect 38577 5426 38605 5427
rect 38617 5426 38645 5427
rect 38657 5426 38685 5427
rect 38697 5426 38725 5427
rect 19527 5181 19555 5182
rect 19567 5181 19595 5182
rect 19607 5181 19635 5182
rect 19647 5181 19675 5182
rect 19527 5155 19550 5181
rect 19550 5155 19555 5181
rect 19567 5155 19582 5181
rect 19582 5155 19588 5181
rect 19588 5155 19595 5181
rect 19607 5155 19614 5181
rect 19614 5155 19620 5181
rect 19620 5155 19635 5181
rect 19647 5155 19652 5181
rect 19652 5155 19675 5181
rect 19527 5154 19555 5155
rect 19567 5154 19595 5155
rect 19607 5154 19635 5155
rect 19647 5154 19675 5155
rect 38577 4909 38605 4910
rect 38617 4909 38645 4910
rect 38657 4909 38685 4910
rect 38697 4909 38725 4910
rect 38577 4883 38600 4909
rect 38600 4883 38605 4909
rect 38617 4883 38632 4909
rect 38632 4883 38638 4909
rect 38638 4883 38645 4909
rect 38657 4883 38664 4909
rect 38664 4883 38670 4909
rect 38670 4883 38685 4909
rect 38697 4883 38702 4909
rect 38702 4883 38725 4909
rect 38577 4882 38605 4883
rect 38617 4882 38645 4883
rect 38657 4882 38685 4883
rect 38697 4882 38725 4883
rect 57626 6813 57654 6814
rect 57666 6813 57694 6814
rect 57706 6813 57734 6814
rect 57746 6813 57774 6814
rect 57626 6787 57649 6813
rect 57649 6787 57654 6813
rect 57666 6787 57681 6813
rect 57681 6787 57687 6813
rect 57687 6787 57694 6813
rect 57706 6787 57713 6813
rect 57713 6787 57719 6813
rect 57719 6787 57734 6813
rect 57746 6787 57751 6813
rect 57751 6787 57774 6813
rect 57626 6786 57654 6787
rect 57666 6786 57694 6787
rect 57706 6786 57734 6787
rect 57746 6786 57774 6787
rect 57626 6269 57654 6270
rect 57666 6269 57694 6270
rect 57706 6269 57734 6270
rect 57746 6269 57774 6270
rect 57626 6243 57649 6269
rect 57649 6243 57654 6269
rect 57666 6243 57681 6269
rect 57681 6243 57687 6269
rect 57687 6243 57694 6269
rect 57706 6243 57713 6269
rect 57713 6243 57719 6269
rect 57719 6243 57734 6269
rect 57746 6243 57751 6269
rect 57751 6243 57774 6269
rect 57626 6242 57654 6243
rect 57666 6242 57694 6243
rect 57706 6242 57734 6243
rect 57746 6242 57774 6243
rect 57626 5725 57654 5726
rect 57666 5725 57694 5726
rect 57706 5725 57734 5726
rect 57746 5725 57774 5726
rect 57626 5699 57649 5725
rect 57649 5699 57654 5725
rect 57666 5699 57681 5725
rect 57681 5699 57687 5725
rect 57687 5699 57694 5725
rect 57706 5699 57713 5725
rect 57713 5699 57719 5725
rect 57719 5699 57734 5725
rect 57746 5699 57751 5725
rect 57751 5699 57774 5725
rect 57626 5698 57654 5699
rect 57666 5698 57694 5699
rect 57706 5698 57734 5699
rect 57746 5698 57774 5699
rect 57626 5181 57654 5182
rect 57666 5181 57694 5182
rect 57706 5181 57734 5182
rect 57746 5181 57774 5182
rect 57626 5155 57649 5181
rect 57649 5155 57654 5181
rect 57666 5155 57681 5181
rect 57681 5155 57687 5181
rect 57687 5155 57694 5181
rect 57706 5155 57713 5181
rect 57713 5155 57719 5181
rect 57719 5155 57734 5181
rect 57746 5155 57751 5181
rect 57751 5155 57774 5181
rect 57626 5154 57654 5155
rect 57666 5154 57694 5155
rect 57706 5154 57734 5155
rect 57746 5154 57774 5155
rect 19527 4637 19555 4638
rect 19567 4637 19595 4638
rect 19607 4637 19635 4638
rect 19647 4637 19675 4638
rect 19527 4611 19550 4637
rect 19550 4611 19555 4637
rect 19567 4611 19582 4637
rect 19582 4611 19588 4637
rect 19588 4611 19595 4637
rect 19607 4611 19614 4637
rect 19614 4611 19620 4637
rect 19620 4611 19635 4637
rect 19647 4611 19652 4637
rect 19652 4611 19675 4637
rect 19527 4610 19555 4611
rect 19567 4610 19595 4611
rect 19607 4610 19635 4611
rect 19647 4610 19675 4611
rect 57626 4637 57654 4638
rect 57666 4637 57694 4638
rect 57706 4637 57734 4638
rect 57746 4637 57774 4638
rect 57626 4611 57649 4637
rect 57649 4611 57654 4637
rect 57666 4611 57681 4637
rect 57681 4611 57687 4637
rect 57687 4611 57694 4637
rect 57706 4611 57713 4637
rect 57713 4611 57719 4637
rect 57719 4611 57734 4637
rect 57746 4611 57751 4637
rect 57751 4611 57774 4637
rect 57626 4610 57654 4611
rect 57666 4610 57694 4611
rect 57706 4610 57734 4611
rect 57746 4610 57774 4611
rect 38577 4365 38605 4366
rect 38617 4365 38645 4366
rect 38657 4365 38685 4366
rect 38697 4365 38725 4366
rect 38577 4339 38600 4365
rect 38600 4339 38605 4365
rect 38617 4339 38632 4365
rect 38632 4339 38638 4365
rect 38638 4339 38645 4365
rect 38657 4339 38664 4365
rect 38664 4339 38670 4365
rect 38670 4339 38685 4365
rect 38697 4339 38702 4365
rect 38702 4339 38725 4365
rect 38577 4338 38605 4339
rect 38617 4338 38645 4339
rect 38657 4338 38685 4339
rect 38697 4338 38725 4339
rect 19527 4093 19555 4094
rect 19567 4093 19595 4094
rect 19607 4093 19635 4094
rect 19647 4093 19675 4094
rect 19527 4067 19550 4093
rect 19550 4067 19555 4093
rect 19567 4067 19582 4093
rect 19582 4067 19588 4093
rect 19588 4067 19595 4093
rect 19607 4067 19614 4093
rect 19614 4067 19620 4093
rect 19620 4067 19635 4093
rect 19647 4067 19652 4093
rect 19652 4067 19675 4093
rect 19527 4066 19555 4067
rect 19567 4066 19595 4067
rect 19607 4066 19635 4067
rect 19647 4066 19675 4067
rect 57626 4093 57654 4094
rect 57666 4093 57694 4094
rect 57706 4093 57734 4094
rect 57746 4093 57774 4094
rect 57626 4067 57649 4093
rect 57649 4067 57654 4093
rect 57666 4067 57681 4093
rect 57681 4067 57687 4093
rect 57687 4067 57694 4093
rect 57706 4067 57713 4093
rect 57713 4067 57719 4093
rect 57719 4067 57734 4093
rect 57746 4067 57751 4093
rect 57751 4067 57774 4093
rect 57626 4066 57654 4067
rect 57666 4066 57694 4067
rect 57706 4066 57734 4067
rect 57746 4066 57774 4067
rect 699 4032 727 4060
rect 38577 3821 38605 3822
rect 38617 3821 38645 3822
rect 38657 3821 38685 3822
rect 38697 3821 38725 3822
rect 38577 3795 38600 3821
rect 38600 3795 38605 3821
rect 38617 3795 38632 3821
rect 38632 3795 38638 3821
rect 38638 3795 38645 3821
rect 38657 3795 38664 3821
rect 38664 3795 38670 3821
rect 38670 3795 38685 3821
rect 38697 3795 38702 3821
rect 38702 3795 38725 3821
rect 38577 3794 38605 3795
rect 38617 3794 38645 3795
rect 38657 3794 38685 3795
rect 38697 3794 38725 3795
rect 19527 3549 19555 3550
rect 19567 3549 19595 3550
rect 19607 3549 19635 3550
rect 19647 3549 19675 3550
rect 19527 3523 19550 3549
rect 19550 3523 19555 3549
rect 19567 3523 19582 3549
rect 19582 3523 19588 3549
rect 19588 3523 19595 3549
rect 19607 3523 19614 3549
rect 19614 3523 19620 3549
rect 19620 3523 19635 3549
rect 19647 3523 19652 3549
rect 19652 3523 19675 3549
rect 19527 3522 19555 3523
rect 19567 3522 19595 3523
rect 19607 3522 19635 3523
rect 19647 3522 19675 3523
rect 57626 3549 57654 3550
rect 57666 3549 57694 3550
rect 57706 3549 57734 3550
rect 57746 3549 57774 3550
rect 57626 3523 57649 3549
rect 57649 3523 57654 3549
rect 57666 3523 57681 3549
rect 57681 3523 57687 3549
rect 57687 3523 57694 3549
rect 57706 3523 57713 3549
rect 57713 3523 57719 3549
rect 57719 3523 57734 3549
rect 57746 3523 57751 3549
rect 57751 3523 57774 3549
rect 57626 3522 57654 3523
rect 57666 3522 57694 3523
rect 57706 3522 57734 3523
rect 57746 3522 57774 3523
rect 38577 3277 38605 3278
rect 38617 3277 38645 3278
rect 38657 3277 38685 3278
rect 38697 3277 38725 3278
rect 38577 3251 38600 3277
rect 38600 3251 38605 3277
rect 38617 3251 38632 3277
rect 38632 3251 38638 3277
rect 38638 3251 38645 3277
rect 38657 3251 38664 3277
rect 38664 3251 38670 3277
rect 38670 3251 38685 3277
rect 38697 3251 38702 3277
rect 38702 3251 38725 3277
rect 38577 3250 38605 3251
rect 38617 3250 38645 3251
rect 38657 3250 38685 3251
rect 38697 3250 38725 3251
rect 19527 3005 19555 3006
rect 19567 3005 19595 3006
rect 19607 3005 19635 3006
rect 19647 3005 19675 3006
rect 19527 2979 19550 3005
rect 19550 2979 19555 3005
rect 19567 2979 19582 3005
rect 19582 2979 19588 3005
rect 19588 2979 19595 3005
rect 19607 2979 19614 3005
rect 19614 2979 19620 3005
rect 19620 2979 19635 3005
rect 19647 2979 19652 3005
rect 19652 2979 19675 3005
rect 19527 2978 19555 2979
rect 19567 2978 19595 2979
rect 19607 2978 19635 2979
rect 19647 2978 19675 2979
rect 57626 3005 57654 3006
rect 57666 3005 57694 3006
rect 57706 3005 57734 3006
rect 57746 3005 57774 3006
rect 57626 2979 57649 3005
rect 57649 2979 57654 3005
rect 57666 2979 57681 3005
rect 57681 2979 57687 3005
rect 57687 2979 57694 3005
rect 57706 2979 57713 3005
rect 57713 2979 57719 3005
rect 57719 2979 57734 3005
rect 57746 2979 57751 3005
rect 57751 2979 57774 3005
rect 57626 2978 57654 2979
rect 57666 2978 57694 2979
rect 57706 2978 57734 2979
rect 57746 2978 57774 2979
rect 38577 2733 38605 2734
rect 38617 2733 38645 2734
rect 38657 2733 38685 2734
rect 38697 2733 38725 2734
rect 38577 2707 38600 2733
rect 38600 2707 38605 2733
rect 38617 2707 38632 2733
rect 38632 2707 38638 2733
rect 38638 2707 38645 2733
rect 38657 2707 38664 2733
rect 38664 2707 38670 2733
rect 38670 2707 38685 2733
rect 38697 2707 38702 2733
rect 38702 2707 38725 2733
rect 38577 2706 38605 2707
rect 38617 2706 38645 2707
rect 38657 2706 38685 2707
rect 38697 2706 38725 2707
rect 19527 2461 19555 2462
rect 19567 2461 19595 2462
rect 19607 2461 19635 2462
rect 19647 2461 19675 2462
rect 19527 2435 19550 2461
rect 19550 2435 19555 2461
rect 19567 2435 19582 2461
rect 19582 2435 19588 2461
rect 19588 2435 19595 2461
rect 19607 2435 19614 2461
rect 19614 2435 19620 2461
rect 19620 2435 19635 2461
rect 19647 2435 19652 2461
rect 19652 2435 19675 2461
rect 19527 2434 19555 2435
rect 19567 2434 19595 2435
rect 19607 2434 19635 2435
rect 19647 2434 19675 2435
rect 57626 2461 57654 2462
rect 57666 2461 57694 2462
rect 57706 2461 57734 2462
rect 57746 2461 57774 2462
rect 57626 2435 57649 2461
rect 57649 2435 57654 2461
rect 57666 2435 57681 2461
rect 57681 2435 57687 2461
rect 57687 2435 57694 2461
rect 57706 2435 57713 2461
rect 57713 2435 57719 2461
rect 57719 2435 57734 2461
rect 57746 2435 57751 2461
rect 57751 2435 57774 2461
rect 57626 2434 57654 2435
rect 57666 2434 57694 2435
rect 57706 2434 57734 2435
rect 57746 2434 57774 2435
rect 38577 2189 38605 2190
rect 38617 2189 38645 2190
rect 38657 2189 38685 2190
rect 38697 2189 38725 2190
rect 38577 2163 38600 2189
rect 38600 2163 38605 2189
rect 38617 2163 38632 2189
rect 38632 2163 38638 2189
rect 38638 2163 38645 2189
rect 38657 2163 38664 2189
rect 38664 2163 38670 2189
rect 38670 2163 38685 2189
rect 38697 2163 38702 2189
rect 38702 2163 38725 2189
rect 38577 2162 38605 2163
rect 38617 2162 38645 2163
rect 38657 2162 38685 2163
rect 38697 2162 38725 2163
rect 19527 1917 19555 1918
rect 19567 1917 19595 1918
rect 19607 1917 19635 1918
rect 19647 1917 19675 1918
rect 19527 1891 19550 1917
rect 19550 1891 19555 1917
rect 19567 1891 19582 1917
rect 19582 1891 19588 1917
rect 19588 1891 19595 1917
rect 19607 1891 19614 1917
rect 19614 1891 19620 1917
rect 19620 1891 19635 1917
rect 19647 1891 19652 1917
rect 19652 1891 19675 1917
rect 19527 1890 19555 1891
rect 19567 1890 19595 1891
rect 19607 1890 19635 1891
rect 19647 1890 19675 1891
rect 57626 1917 57654 1918
rect 57666 1917 57694 1918
rect 57706 1917 57734 1918
rect 57746 1917 57774 1918
rect 57626 1891 57649 1917
rect 57649 1891 57654 1917
rect 57666 1891 57681 1917
rect 57681 1891 57687 1917
rect 57687 1891 57694 1917
rect 57706 1891 57713 1917
rect 57713 1891 57719 1917
rect 57719 1891 57734 1917
rect 57746 1891 57751 1917
rect 57751 1891 57774 1917
rect 57626 1890 57654 1891
rect 57666 1890 57694 1891
rect 57706 1890 57734 1891
rect 57746 1890 57774 1891
rect 38577 1645 38605 1646
rect 38617 1645 38645 1646
rect 38657 1645 38685 1646
rect 38697 1645 38725 1646
rect 38577 1619 38600 1645
rect 38600 1619 38605 1645
rect 38617 1619 38632 1645
rect 38632 1619 38638 1645
rect 38638 1619 38645 1645
rect 38657 1619 38664 1645
rect 38664 1619 38670 1645
rect 38670 1619 38685 1645
rect 38697 1619 38702 1645
rect 38702 1619 38725 1645
rect 38577 1618 38605 1619
rect 38617 1618 38645 1619
rect 38657 1618 38685 1619
rect 38697 1618 38725 1619
rect 19527 1373 19555 1374
rect 19567 1373 19595 1374
rect 19607 1373 19635 1374
rect 19647 1373 19675 1374
rect 19527 1347 19550 1373
rect 19550 1347 19555 1373
rect 19567 1347 19582 1373
rect 19582 1347 19588 1373
rect 19588 1347 19595 1373
rect 19607 1347 19614 1373
rect 19614 1347 19620 1373
rect 19620 1347 19635 1373
rect 19647 1347 19652 1373
rect 19652 1347 19675 1373
rect 19527 1346 19555 1347
rect 19567 1346 19595 1347
rect 19607 1346 19635 1347
rect 19647 1346 19675 1347
rect 57626 1373 57654 1374
rect 57666 1373 57694 1374
rect 57706 1373 57734 1374
rect 57746 1373 57774 1374
rect 57626 1347 57649 1373
rect 57649 1347 57654 1373
rect 57666 1347 57681 1373
rect 57681 1347 57687 1373
rect 57687 1347 57694 1373
rect 57706 1347 57713 1373
rect 57713 1347 57719 1373
rect 57719 1347 57734 1373
rect 57746 1347 57751 1373
rect 57751 1347 57774 1373
rect 57626 1346 57654 1347
rect 57666 1346 57694 1347
rect 57706 1346 57734 1347
rect 57746 1346 57774 1347
rect 76676 6541 76704 6542
rect 76716 6541 76744 6542
rect 76756 6541 76784 6542
rect 76796 6541 76824 6542
rect 76676 6515 76699 6541
rect 76699 6515 76704 6541
rect 76716 6515 76731 6541
rect 76731 6515 76737 6541
rect 76737 6515 76744 6541
rect 76756 6515 76763 6541
rect 76763 6515 76769 6541
rect 76769 6515 76784 6541
rect 76796 6515 76801 6541
rect 76801 6515 76824 6541
rect 76676 6514 76704 6515
rect 76716 6514 76744 6515
rect 76756 6514 76784 6515
rect 76796 6514 76824 6515
rect 76676 5997 76704 5998
rect 76716 5997 76744 5998
rect 76756 5997 76784 5998
rect 76796 5997 76824 5998
rect 76676 5971 76699 5997
rect 76699 5971 76704 5997
rect 76716 5971 76731 5997
rect 76731 5971 76737 5997
rect 76737 5971 76744 5997
rect 76756 5971 76763 5997
rect 76763 5971 76769 5997
rect 76769 5971 76784 5997
rect 76796 5971 76801 5997
rect 76801 5971 76824 5997
rect 76676 5970 76704 5971
rect 76716 5970 76744 5971
rect 76756 5970 76784 5971
rect 76796 5970 76824 5971
rect 77519 6412 77547 6440
rect 78945 6294 78946 6304
rect 78946 6294 78972 6304
rect 78972 6294 78973 6304
rect 78945 6276 78973 6294
rect 76676 5453 76704 5454
rect 76716 5453 76744 5454
rect 76756 5453 76784 5454
rect 76796 5453 76824 5454
rect 76676 5427 76699 5453
rect 76699 5427 76704 5453
rect 76716 5427 76731 5453
rect 76731 5427 76737 5453
rect 76737 5427 76744 5453
rect 76756 5427 76763 5453
rect 76763 5427 76769 5453
rect 76769 5427 76784 5453
rect 76796 5427 76801 5453
rect 76801 5427 76824 5453
rect 76676 5426 76704 5427
rect 76716 5426 76744 5427
rect 76756 5426 76784 5427
rect 76796 5426 76824 5427
rect 76676 4909 76704 4910
rect 76716 4909 76744 4910
rect 76756 4909 76784 4910
rect 76796 4909 76824 4910
rect 76676 4883 76699 4909
rect 76699 4883 76704 4909
rect 76716 4883 76731 4909
rect 76731 4883 76737 4909
rect 76737 4883 76744 4909
rect 76756 4883 76763 4909
rect 76763 4883 76769 4909
rect 76769 4883 76784 4909
rect 76796 4883 76801 4909
rect 76801 4883 76824 4909
rect 76676 4882 76704 4883
rect 76716 4882 76744 4883
rect 76756 4882 76784 4883
rect 76796 4882 76824 4883
rect 80141 6294 80142 6304
rect 80142 6294 80168 6304
rect 80168 6294 80169 6304
rect 80141 6276 80169 6294
rect 81797 6150 81825 6168
rect 81797 6140 81798 6150
rect 81798 6140 81824 6150
rect 81824 6140 81825 6150
rect 94815 5878 94843 5896
rect 94815 5868 94816 5878
rect 94816 5868 94842 5878
rect 94842 5868 94843 5878
rect 76676 4365 76704 4366
rect 76716 4365 76744 4366
rect 76756 4365 76784 4366
rect 76796 4365 76824 4366
rect 76676 4339 76699 4365
rect 76699 4339 76704 4365
rect 76716 4339 76731 4365
rect 76731 4339 76737 4365
rect 76737 4339 76744 4365
rect 76756 4339 76763 4365
rect 76763 4339 76769 4365
rect 76769 4339 76784 4365
rect 76796 4339 76801 4365
rect 76801 4339 76824 4365
rect 76676 4338 76704 4339
rect 76716 4338 76744 4339
rect 76756 4338 76784 4339
rect 76796 4338 76824 4339
rect 95725 6813 95753 6814
rect 95765 6813 95793 6814
rect 95805 6813 95833 6814
rect 95845 6813 95873 6814
rect 95725 6787 95748 6813
rect 95748 6787 95753 6813
rect 95765 6787 95780 6813
rect 95780 6787 95786 6813
rect 95786 6787 95793 6813
rect 95805 6787 95812 6813
rect 95812 6787 95818 6813
rect 95818 6787 95833 6813
rect 95845 6787 95850 6813
rect 95850 6787 95873 6813
rect 95725 6786 95753 6787
rect 95765 6786 95793 6787
rect 95805 6786 95833 6787
rect 95845 6786 95873 6787
rect 95919 6276 95947 6304
rect 95725 6269 95753 6270
rect 95765 6269 95793 6270
rect 95805 6269 95833 6270
rect 95845 6269 95873 6270
rect 95725 6243 95748 6269
rect 95748 6243 95753 6269
rect 95765 6243 95780 6269
rect 95780 6243 95786 6269
rect 95786 6243 95793 6269
rect 95805 6243 95812 6269
rect 95812 6243 95818 6269
rect 95818 6243 95833 6269
rect 95845 6243 95850 6269
rect 95850 6243 95873 6269
rect 95725 6242 95753 6243
rect 95765 6242 95793 6243
rect 95805 6242 95833 6243
rect 95845 6242 95873 6243
rect 96103 6276 96131 6304
rect 95725 5725 95753 5726
rect 95765 5725 95793 5726
rect 95805 5725 95833 5726
rect 95845 5725 95873 5726
rect 95725 5699 95748 5725
rect 95748 5699 95753 5725
rect 95765 5699 95780 5725
rect 95780 5699 95786 5725
rect 95786 5699 95793 5725
rect 95805 5699 95812 5725
rect 95812 5699 95818 5725
rect 95818 5699 95833 5725
rect 95845 5699 95850 5725
rect 95850 5699 95873 5725
rect 95725 5698 95753 5699
rect 95765 5698 95793 5699
rect 95805 5698 95833 5699
rect 95845 5698 95873 5699
rect 95725 5181 95753 5182
rect 95765 5181 95793 5182
rect 95805 5181 95833 5182
rect 95845 5181 95873 5182
rect 95725 5155 95748 5181
rect 95748 5155 95753 5181
rect 95765 5155 95780 5181
rect 95780 5155 95786 5181
rect 95786 5155 95793 5181
rect 95805 5155 95812 5181
rect 95812 5155 95818 5181
rect 95818 5155 95833 5181
rect 95845 5155 95850 5181
rect 95850 5155 95873 5181
rect 95725 5154 95753 5155
rect 95765 5154 95793 5155
rect 95805 5154 95833 5155
rect 95845 5154 95873 5155
rect 96517 6140 96545 6168
rect 96517 5868 96545 5896
rect 97299 6412 97327 6440
rect 97529 6344 97557 6372
rect 97897 6412 97925 6440
rect 98679 6422 98707 6440
rect 98679 6412 98680 6422
rect 98680 6412 98706 6422
rect 98706 6412 98707 6422
rect 100427 6616 100455 6644
rect 100197 6276 100225 6304
rect 101715 6616 101743 6644
rect 103555 6762 103583 6780
rect 103555 6752 103556 6762
rect 103556 6752 103582 6762
rect 103582 6752 103583 6762
rect 102773 6616 102801 6644
rect 102635 6294 102636 6304
rect 102636 6294 102662 6304
rect 102662 6294 102663 6304
rect 102635 6276 102663 6294
rect 102865 6616 102893 6644
rect 103601 6634 103602 6644
rect 103602 6634 103628 6644
rect 103628 6634 103629 6644
rect 103601 6616 103629 6634
rect 104015 6752 104043 6780
rect 106637 6702 106638 6712
rect 106638 6702 106664 6712
rect 106664 6702 106665 6712
rect 106637 6684 106665 6702
rect 109903 6684 109931 6712
rect 103969 6634 103970 6644
rect 103970 6634 103996 6644
rect 103996 6634 103997 6644
rect 103969 6616 103997 6634
rect 103923 6344 103951 6372
rect 112709 6566 112710 6576
rect 112710 6566 112736 6576
rect 112736 6566 112737 6576
rect 112709 6548 112737 6566
rect 113537 6694 113565 6712
rect 113537 6684 113538 6694
rect 113538 6684 113564 6694
rect 113564 6684 113565 6694
rect 113537 6566 113538 6576
rect 113538 6566 113564 6576
rect 113564 6566 113565 6576
rect 113537 6548 113565 6566
rect 114595 6702 114596 6712
rect 114596 6702 114622 6712
rect 114622 6702 114623 6712
rect 114595 6684 114623 6702
rect 115193 6634 115194 6644
rect 115194 6634 115220 6644
rect 115220 6634 115221 6644
rect 115193 6616 115221 6634
rect 114775 6541 114803 6542
rect 114815 6541 114843 6542
rect 114855 6541 114883 6542
rect 114895 6541 114923 6542
rect 114775 6515 114798 6541
rect 114798 6515 114803 6541
rect 114815 6515 114830 6541
rect 114830 6515 114836 6541
rect 114836 6515 114843 6541
rect 114855 6515 114862 6541
rect 114862 6515 114868 6541
rect 114868 6515 114883 6541
rect 114895 6515 114900 6541
rect 114900 6515 114923 6541
rect 114775 6514 114803 6515
rect 114815 6514 114843 6515
rect 114855 6514 114883 6515
rect 114895 6514 114923 6515
rect 114775 5997 114803 5998
rect 114815 5997 114843 5998
rect 114855 5997 114883 5998
rect 114895 5997 114923 5998
rect 114775 5971 114798 5997
rect 114798 5971 114803 5997
rect 114815 5971 114830 5997
rect 114830 5971 114836 5997
rect 114836 5971 114843 5997
rect 114855 5971 114862 5997
rect 114862 5971 114868 5997
rect 114868 5971 114883 5997
rect 114895 5971 114900 5997
rect 114900 5971 114923 5997
rect 114775 5970 114803 5971
rect 114815 5970 114843 5971
rect 114855 5970 114883 5971
rect 114895 5970 114923 5971
rect 116067 6616 116095 6644
rect 119057 6694 119085 6712
rect 119057 6684 119058 6694
rect 119058 6684 119084 6694
rect 119084 6684 119085 6694
rect 119747 6702 119748 6712
rect 119748 6702 119774 6712
rect 119774 6702 119775 6712
rect 119747 6684 119775 6702
rect 119149 6344 119177 6372
rect 121081 6354 121109 6372
rect 121081 6344 121082 6354
rect 121082 6344 121108 6354
rect 121108 6344 121109 6354
rect 114775 5453 114803 5454
rect 114815 5453 114843 5454
rect 114855 5453 114883 5454
rect 114895 5453 114923 5454
rect 114775 5427 114798 5453
rect 114798 5427 114803 5453
rect 114815 5427 114830 5453
rect 114830 5427 114836 5453
rect 114836 5427 114843 5453
rect 114855 5427 114862 5453
rect 114862 5427 114868 5453
rect 114868 5427 114883 5453
rect 114895 5427 114900 5453
rect 114900 5427 114923 5453
rect 114775 5426 114803 5427
rect 114815 5426 114843 5427
rect 114855 5426 114883 5427
rect 114895 5426 114923 5427
rect 114775 4909 114803 4910
rect 114815 4909 114843 4910
rect 114855 4909 114883 4910
rect 114895 4909 114923 4910
rect 114775 4883 114798 4909
rect 114798 4883 114803 4909
rect 114815 4883 114830 4909
rect 114830 4883 114836 4909
rect 114836 4883 114843 4909
rect 114855 4883 114862 4909
rect 114862 4883 114868 4909
rect 114868 4883 114883 4909
rect 114895 4883 114900 4909
rect 114900 4883 114923 4909
rect 114775 4882 114803 4883
rect 114815 4882 114843 4883
rect 114855 4882 114883 4883
rect 114895 4882 114923 4883
rect 95725 4637 95753 4638
rect 95765 4637 95793 4638
rect 95805 4637 95833 4638
rect 95845 4637 95873 4638
rect 95725 4611 95748 4637
rect 95748 4611 95753 4637
rect 95765 4611 95780 4637
rect 95780 4611 95786 4637
rect 95786 4611 95793 4637
rect 95805 4611 95812 4637
rect 95812 4611 95818 4637
rect 95818 4611 95833 4637
rect 95845 4611 95850 4637
rect 95850 4611 95873 4637
rect 95725 4610 95753 4611
rect 95765 4610 95793 4611
rect 95805 4610 95833 4611
rect 95845 4610 95873 4611
rect 114775 4365 114803 4366
rect 114815 4365 114843 4366
rect 114855 4365 114883 4366
rect 114895 4365 114923 4366
rect 114775 4339 114798 4365
rect 114798 4339 114803 4365
rect 114815 4339 114830 4365
rect 114830 4339 114836 4365
rect 114836 4339 114843 4365
rect 114855 4339 114862 4365
rect 114862 4339 114868 4365
rect 114868 4339 114883 4365
rect 114895 4339 114900 4365
rect 114900 4339 114923 4365
rect 114775 4338 114803 4339
rect 114815 4338 114843 4339
rect 114855 4338 114883 4339
rect 114895 4338 114923 4339
rect 95725 4093 95753 4094
rect 95765 4093 95793 4094
rect 95805 4093 95833 4094
rect 95845 4093 95873 4094
rect 95725 4067 95748 4093
rect 95748 4067 95753 4093
rect 95765 4067 95780 4093
rect 95780 4067 95786 4093
rect 95786 4067 95793 4093
rect 95805 4067 95812 4093
rect 95812 4067 95818 4093
rect 95818 4067 95833 4093
rect 95845 4067 95850 4093
rect 95850 4067 95873 4093
rect 95725 4066 95753 4067
rect 95765 4066 95793 4067
rect 95805 4066 95833 4067
rect 95845 4066 95873 4067
rect 76676 3821 76704 3822
rect 76716 3821 76744 3822
rect 76756 3821 76784 3822
rect 76796 3821 76824 3822
rect 76676 3795 76699 3821
rect 76699 3795 76704 3821
rect 76716 3795 76731 3821
rect 76731 3795 76737 3821
rect 76737 3795 76744 3821
rect 76756 3795 76763 3821
rect 76763 3795 76769 3821
rect 76769 3795 76784 3821
rect 76796 3795 76801 3821
rect 76801 3795 76824 3821
rect 76676 3794 76704 3795
rect 76716 3794 76744 3795
rect 76756 3794 76784 3795
rect 76796 3794 76824 3795
rect 114775 3821 114803 3822
rect 114815 3821 114843 3822
rect 114855 3821 114883 3822
rect 114895 3821 114923 3822
rect 114775 3795 114798 3821
rect 114798 3795 114803 3821
rect 114815 3795 114830 3821
rect 114830 3795 114836 3821
rect 114836 3795 114843 3821
rect 114855 3795 114862 3821
rect 114862 3795 114868 3821
rect 114868 3795 114883 3821
rect 114895 3795 114900 3821
rect 114900 3795 114923 3821
rect 114775 3794 114803 3795
rect 114815 3794 114843 3795
rect 114855 3794 114883 3795
rect 114895 3794 114923 3795
rect 95725 3549 95753 3550
rect 95765 3549 95793 3550
rect 95805 3549 95833 3550
rect 95845 3549 95873 3550
rect 95725 3523 95748 3549
rect 95748 3523 95753 3549
rect 95765 3523 95780 3549
rect 95780 3523 95786 3549
rect 95786 3523 95793 3549
rect 95805 3523 95812 3549
rect 95812 3523 95818 3549
rect 95818 3523 95833 3549
rect 95845 3523 95850 3549
rect 95850 3523 95873 3549
rect 95725 3522 95753 3523
rect 95765 3522 95793 3523
rect 95805 3522 95833 3523
rect 95845 3522 95873 3523
rect 76676 3277 76704 3278
rect 76716 3277 76744 3278
rect 76756 3277 76784 3278
rect 76796 3277 76824 3278
rect 76676 3251 76699 3277
rect 76699 3251 76704 3277
rect 76716 3251 76731 3277
rect 76731 3251 76737 3277
rect 76737 3251 76744 3277
rect 76756 3251 76763 3277
rect 76763 3251 76769 3277
rect 76769 3251 76784 3277
rect 76796 3251 76801 3277
rect 76801 3251 76824 3277
rect 76676 3250 76704 3251
rect 76716 3250 76744 3251
rect 76756 3250 76784 3251
rect 76796 3250 76824 3251
rect 114775 3277 114803 3278
rect 114815 3277 114843 3278
rect 114855 3277 114883 3278
rect 114895 3277 114923 3278
rect 114775 3251 114798 3277
rect 114798 3251 114803 3277
rect 114815 3251 114830 3277
rect 114830 3251 114836 3277
rect 114836 3251 114843 3277
rect 114855 3251 114862 3277
rect 114862 3251 114868 3277
rect 114868 3251 114883 3277
rect 114895 3251 114900 3277
rect 114900 3251 114923 3277
rect 114775 3250 114803 3251
rect 114815 3250 114843 3251
rect 114855 3250 114883 3251
rect 114895 3250 114923 3251
rect 125957 6294 125958 6304
rect 125958 6294 125984 6304
rect 125984 6294 125985 6304
rect 125957 6276 125985 6294
rect 125911 6208 125939 6236
rect 128303 6480 128331 6508
rect 128993 6480 129021 6508
rect 128533 6276 128561 6304
rect 128579 6208 128607 6236
rect 131155 6362 131156 6372
rect 131156 6362 131182 6372
rect 131182 6362 131183 6372
rect 131155 6344 131183 6362
rect 131707 6626 131735 6644
rect 131707 6616 131708 6626
rect 131708 6616 131734 6626
rect 131734 6616 131735 6626
rect 131753 6354 131781 6372
rect 131753 6344 131754 6354
rect 131754 6344 131780 6354
rect 131780 6344 131781 6354
rect 132167 6344 132195 6372
rect 133824 6813 133852 6814
rect 133864 6813 133892 6814
rect 133904 6813 133932 6814
rect 133944 6813 133972 6814
rect 133824 6787 133847 6813
rect 133847 6787 133852 6813
rect 133864 6787 133879 6813
rect 133879 6787 133885 6813
rect 133885 6787 133892 6813
rect 133904 6787 133911 6813
rect 133911 6787 133917 6813
rect 133917 6787 133932 6813
rect 133944 6787 133949 6813
rect 133949 6787 133972 6813
rect 133824 6786 133852 6787
rect 133864 6786 133892 6787
rect 133904 6786 133932 6787
rect 133944 6786 133972 6787
rect 132765 6616 132793 6644
rect 133547 6344 133575 6372
rect 133823 6344 133851 6372
rect 133824 6269 133852 6270
rect 133864 6269 133892 6270
rect 133904 6269 133932 6270
rect 133944 6269 133972 6270
rect 133824 6243 133847 6269
rect 133847 6243 133852 6269
rect 133864 6243 133879 6269
rect 133879 6243 133885 6269
rect 133885 6243 133892 6269
rect 133904 6243 133911 6269
rect 133911 6243 133917 6269
rect 133917 6243 133932 6269
rect 133944 6243 133949 6269
rect 133949 6243 133972 6269
rect 133824 6242 133852 6243
rect 133864 6242 133892 6243
rect 133904 6242 133932 6243
rect 133944 6242 133972 6243
rect 134053 6344 134081 6372
rect 133824 5725 133852 5726
rect 133864 5725 133892 5726
rect 133904 5725 133932 5726
rect 133944 5725 133972 5726
rect 133824 5699 133847 5725
rect 133847 5699 133852 5725
rect 133864 5699 133879 5725
rect 133879 5699 133885 5725
rect 133885 5699 133892 5725
rect 133904 5699 133911 5725
rect 133911 5699 133917 5725
rect 133917 5699 133932 5725
rect 133944 5699 133949 5725
rect 133949 5699 133972 5725
rect 133824 5698 133852 5699
rect 133864 5698 133892 5699
rect 133904 5698 133932 5699
rect 133944 5698 133972 5699
rect 133824 5181 133852 5182
rect 133864 5181 133892 5182
rect 133904 5181 133932 5182
rect 133944 5181 133972 5182
rect 133824 5155 133847 5181
rect 133847 5155 133852 5181
rect 133864 5155 133879 5181
rect 133879 5155 133885 5181
rect 133885 5155 133892 5181
rect 133904 5155 133911 5181
rect 133911 5155 133917 5181
rect 133917 5155 133932 5181
rect 133944 5155 133949 5181
rect 133949 5155 133972 5181
rect 133824 5154 133852 5155
rect 133864 5154 133892 5155
rect 133904 5154 133932 5155
rect 133944 5154 133972 5155
rect 134467 6684 134495 6712
rect 134513 6616 134541 6644
rect 136583 6694 136611 6712
rect 136583 6684 136584 6694
rect 136584 6684 136610 6694
rect 136610 6684 136611 6694
rect 136629 6634 136630 6644
rect 136630 6634 136656 6644
rect 136656 6634 136657 6644
rect 136629 6616 136657 6634
rect 151763 6956 151791 6984
rect 149739 6412 149767 6440
rect 152223 5002 152224 5012
rect 152224 5002 152250 5012
rect 152250 5002 152251 5012
rect 152223 4984 152251 5002
rect 133824 4637 133852 4638
rect 133864 4637 133892 4638
rect 133904 4637 133932 4638
rect 133944 4637 133972 4638
rect 133824 4611 133847 4637
rect 133847 4611 133852 4637
rect 133864 4611 133879 4637
rect 133879 4611 133885 4637
rect 133885 4611 133892 4637
rect 133904 4611 133911 4637
rect 133911 4611 133917 4637
rect 133917 4611 133932 4637
rect 133944 4611 133949 4637
rect 133949 4611 133972 4637
rect 133824 4610 133852 4611
rect 133864 4610 133892 4611
rect 133904 4610 133932 4611
rect 133944 4610 133972 4611
rect 133824 4093 133852 4094
rect 133864 4093 133892 4094
rect 133904 4093 133932 4094
rect 133944 4093 133972 4094
rect 133824 4067 133847 4093
rect 133847 4067 133852 4093
rect 133864 4067 133879 4093
rect 133879 4067 133885 4093
rect 133885 4067 133892 4093
rect 133904 4067 133911 4093
rect 133911 4067 133917 4093
rect 133917 4067 133932 4093
rect 133944 4067 133949 4093
rect 133949 4067 133972 4093
rect 133824 4066 133852 4067
rect 133864 4066 133892 4067
rect 133904 4066 133932 4067
rect 133944 4066 133972 4067
rect 133824 3549 133852 3550
rect 133864 3549 133892 3550
rect 133904 3549 133932 3550
rect 133944 3549 133972 3550
rect 133824 3523 133847 3549
rect 133847 3523 133852 3549
rect 133864 3523 133879 3549
rect 133879 3523 133885 3549
rect 133885 3523 133892 3549
rect 133904 3523 133911 3549
rect 133911 3523 133917 3549
rect 133917 3523 133932 3549
rect 133944 3523 133949 3549
rect 133949 3523 133972 3549
rect 133824 3522 133852 3523
rect 133864 3522 133892 3523
rect 133904 3522 133932 3523
rect 133944 3522 133972 3523
rect 95725 3005 95753 3006
rect 95765 3005 95793 3006
rect 95805 3005 95833 3006
rect 95845 3005 95873 3006
rect 95725 2979 95748 3005
rect 95748 2979 95753 3005
rect 95765 2979 95780 3005
rect 95780 2979 95786 3005
rect 95786 2979 95793 3005
rect 95805 2979 95812 3005
rect 95812 2979 95818 3005
rect 95818 2979 95833 3005
rect 95845 2979 95850 3005
rect 95850 2979 95873 3005
rect 95725 2978 95753 2979
rect 95765 2978 95793 2979
rect 95805 2978 95833 2979
rect 95845 2978 95873 2979
rect 133824 3005 133852 3006
rect 133864 3005 133892 3006
rect 133904 3005 133932 3006
rect 133944 3005 133972 3006
rect 133824 2979 133847 3005
rect 133847 2979 133852 3005
rect 133864 2979 133879 3005
rect 133879 2979 133885 3005
rect 133885 2979 133892 3005
rect 133904 2979 133911 3005
rect 133911 2979 133917 3005
rect 133917 2979 133932 3005
rect 133944 2979 133949 3005
rect 133949 2979 133972 3005
rect 133824 2978 133852 2979
rect 133864 2978 133892 2979
rect 133904 2978 133932 2979
rect 133944 2978 133972 2979
rect 151993 2944 152021 2972
rect 76676 2733 76704 2734
rect 76716 2733 76744 2734
rect 76756 2733 76784 2734
rect 76796 2733 76824 2734
rect 76676 2707 76699 2733
rect 76699 2707 76704 2733
rect 76716 2707 76731 2733
rect 76731 2707 76737 2733
rect 76737 2707 76744 2733
rect 76756 2707 76763 2733
rect 76763 2707 76769 2733
rect 76769 2707 76784 2733
rect 76796 2707 76801 2733
rect 76801 2707 76824 2733
rect 76676 2706 76704 2707
rect 76716 2706 76744 2707
rect 76756 2706 76784 2707
rect 76796 2706 76824 2707
rect 114775 2733 114803 2734
rect 114815 2733 114843 2734
rect 114855 2733 114883 2734
rect 114895 2733 114923 2734
rect 114775 2707 114798 2733
rect 114798 2707 114803 2733
rect 114815 2707 114830 2733
rect 114830 2707 114836 2733
rect 114836 2707 114843 2733
rect 114855 2707 114862 2733
rect 114862 2707 114868 2733
rect 114868 2707 114883 2733
rect 114895 2707 114900 2733
rect 114900 2707 114923 2733
rect 114775 2706 114803 2707
rect 114815 2706 114843 2707
rect 114855 2706 114883 2707
rect 114895 2706 114923 2707
rect 95725 2461 95753 2462
rect 95765 2461 95793 2462
rect 95805 2461 95833 2462
rect 95845 2461 95873 2462
rect 95725 2435 95748 2461
rect 95748 2435 95753 2461
rect 95765 2435 95780 2461
rect 95780 2435 95786 2461
rect 95786 2435 95793 2461
rect 95805 2435 95812 2461
rect 95812 2435 95818 2461
rect 95818 2435 95833 2461
rect 95845 2435 95850 2461
rect 95850 2435 95873 2461
rect 95725 2434 95753 2435
rect 95765 2434 95793 2435
rect 95805 2434 95833 2435
rect 95845 2434 95873 2435
rect 133824 2461 133852 2462
rect 133864 2461 133892 2462
rect 133904 2461 133932 2462
rect 133944 2461 133972 2462
rect 133824 2435 133847 2461
rect 133847 2435 133852 2461
rect 133864 2435 133879 2461
rect 133879 2435 133885 2461
rect 133885 2435 133892 2461
rect 133904 2435 133911 2461
rect 133911 2435 133917 2461
rect 133917 2435 133932 2461
rect 133944 2435 133949 2461
rect 133949 2435 133972 2461
rect 133824 2434 133852 2435
rect 133864 2434 133892 2435
rect 133904 2434 133932 2435
rect 133944 2434 133972 2435
rect 76676 2189 76704 2190
rect 76716 2189 76744 2190
rect 76756 2189 76784 2190
rect 76796 2189 76824 2190
rect 76676 2163 76699 2189
rect 76699 2163 76704 2189
rect 76716 2163 76731 2189
rect 76731 2163 76737 2189
rect 76737 2163 76744 2189
rect 76756 2163 76763 2189
rect 76763 2163 76769 2189
rect 76769 2163 76784 2189
rect 76796 2163 76801 2189
rect 76801 2163 76824 2189
rect 76676 2162 76704 2163
rect 76716 2162 76744 2163
rect 76756 2162 76784 2163
rect 76796 2162 76824 2163
rect 114775 2189 114803 2190
rect 114815 2189 114843 2190
rect 114855 2189 114883 2190
rect 114895 2189 114923 2190
rect 114775 2163 114798 2189
rect 114798 2163 114803 2189
rect 114815 2163 114830 2189
rect 114830 2163 114836 2189
rect 114836 2163 114843 2189
rect 114855 2163 114862 2189
rect 114862 2163 114868 2189
rect 114868 2163 114883 2189
rect 114895 2163 114900 2189
rect 114900 2163 114923 2189
rect 114775 2162 114803 2163
rect 114815 2162 114843 2163
rect 114855 2162 114883 2163
rect 114895 2162 114923 2163
rect 95725 1917 95753 1918
rect 95765 1917 95793 1918
rect 95805 1917 95833 1918
rect 95845 1917 95873 1918
rect 95725 1891 95748 1917
rect 95748 1891 95753 1917
rect 95765 1891 95780 1917
rect 95780 1891 95786 1917
rect 95786 1891 95793 1917
rect 95805 1891 95812 1917
rect 95812 1891 95818 1917
rect 95818 1891 95833 1917
rect 95845 1891 95850 1917
rect 95850 1891 95873 1917
rect 95725 1890 95753 1891
rect 95765 1890 95793 1891
rect 95805 1890 95833 1891
rect 95845 1890 95873 1891
rect 133824 1917 133852 1918
rect 133864 1917 133892 1918
rect 133904 1917 133932 1918
rect 133944 1917 133972 1918
rect 133824 1891 133847 1917
rect 133847 1891 133852 1917
rect 133864 1891 133879 1917
rect 133879 1891 133885 1917
rect 133885 1891 133892 1917
rect 133904 1891 133911 1917
rect 133911 1891 133917 1917
rect 133917 1891 133932 1917
rect 133944 1891 133949 1917
rect 133949 1891 133972 1917
rect 133824 1890 133852 1891
rect 133864 1890 133892 1891
rect 133904 1890 133932 1891
rect 133944 1890 133972 1891
rect 76676 1645 76704 1646
rect 76716 1645 76744 1646
rect 76756 1645 76784 1646
rect 76796 1645 76824 1646
rect 76676 1619 76699 1645
rect 76699 1619 76704 1645
rect 76716 1619 76731 1645
rect 76731 1619 76737 1645
rect 76737 1619 76744 1645
rect 76756 1619 76763 1645
rect 76763 1619 76769 1645
rect 76769 1619 76784 1645
rect 76796 1619 76801 1645
rect 76801 1619 76824 1645
rect 76676 1618 76704 1619
rect 76716 1618 76744 1619
rect 76756 1618 76784 1619
rect 76796 1618 76824 1619
rect 114775 1645 114803 1646
rect 114815 1645 114843 1646
rect 114855 1645 114883 1646
rect 114895 1645 114923 1646
rect 114775 1619 114798 1645
rect 114798 1619 114803 1645
rect 114815 1619 114830 1645
rect 114830 1619 114836 1645
rect 114836 1619 114843 1645
rect 114855 1619 114862 1645
rect 114862 1619 114868 1645
rect 114868 1619 114883 1645
rect 114895 1619 114900 1645
rect 114900 1619 114923 1645
rect 114775 1618 114803 1619
rect 114815 1618 114843 1619
rect 114855 1618 114883 1619
rect 114895 1618 114923 1619
rect 95725 1373 95753 1374
rect 95765 1373 95793 1374
rect 95805 1373 95833 1374
rect 95845 1373 95873 1374
rect 95725 1347 95748 1373
rect 95748 1347 95753 1373
rect 95765 1347 95780 1373
rect 95780 1347 95786 1373
rect 95786 1347 95793 1373
rect 95805 1347 95812 1373
rect 95812 1347 95818 1373
rect 95818 1347 95833 1373
rect 95845 1347 95850 1373
rect 95850 1347 95873 1373
rect 95725 1346 95753 1347
rect 95765 1346 95793 1347
rect 95805 1346 95833 1347
rect 95845 1346 95873 1347
rect 133824 1373 133852 1374
rect 133864 1373 133892 1374
rect 133904 1373 133932 1374
rect 133944 1373 133972 1374
rect 133824 1347 133847 1373
rect 133847 1347 133852 1373
rect 133864 1347 133879 1373
rect 133879 1347 133885 1373
rect 133885 1347 133892 1373
rect 133904 1347 133911 1373
rect 133911 1347 133917 1373
rect 133917 1347 133932 1373
rect 133944 1347 133949 1373
rect 133949 1347 133972 1373
rect 133824 1346 133852 1347
rect 133864 1346 133892 1347
rect 133904 1346 133932 1347
rect 133944 1346 133972 1347
rect 38577 1101 38605 1102
rect 38617 1101 38645 1102
rect 38657 1101 38685 1102
rect 38697 1101 38725 1102
rect 38577 1075 38600 1101
rect 38600 1075 38605 1101
rect 38617 1075 38632 1101
rect 38632 1075 38638 1101
rect 38638 1075 38645 1101
rect 38657 1075 38664 1101
rect 38664 1075 38670 1101
rect 38670 1075 38685 1101
rect 38697 1075 38702 1101
rect 38702 1075 38725 1101
rect 38577 1074 38605 1075
rect 38617 1074 38645 1075
rect 38657 1074 38685 1075
rect 38697 1074 38725 1075
rect 76676 1101 76704 1102
rect 76716 1101 76744 1102
rect 76756 1101 76784 1102
rect 76796 1101 76824 1102
rect 76676 1075 76699 1101
rect 76699 1075 76704 1101
rect 76716 1075 76731 1101
rect 76731 1075 76737 1101
rect 76737 1075 76744 1101
rect 76756 1075 76763 1101
rect 76763 1075 76769 1101
rect 76769 1075 76784 1101
rect 76796 1075 76801 1101
rect 76801 1075 76824 1101
rect 76676 1074 76704 1075
rect 76716 1074 76744 1075
rect 76756 1074 76784 1075
rect 76796 1074 76824 1075
rect 114775 1101 114803 1102
rect 114815 1101 114843 1102
rect 114855 1101 114883 1102
rect 114895 1101 114923 1102
rect 114775 1075 114798 1101
rect 114798 1075 114803 1101
rect 114815 1075 114830 1101
rect 114830 1075 114836 1101
rect 114836 1075 114843 1101
rect 114855 1075 114862 1101
rect 114862 1075 114868 1101
rect 114868 1075 114883 1101
rect 114895 1075 114900 1101
rect 114900 1075 114923 1101
rect 114775 1074 114803 1075
rect 114815 1074 114843 1075
rect 114855 1074 114883 1075
rect 114895 1074 114923 1075
rect 151119 972 151147 1000
<< metal3 >>
rect 151760 6985 151793 6986
rect 153100 6985 153500 7000
rect 151760 6984 153500 6985
rect 151760 6956 151763 6984
rect 151791 6956 153500 6984
rect 151760 6955 153500 6956
rect 151760 6953 151793 6955
rect 153100 6940 153500 6955
rect 19522 6816 19680 6816
rect 19522 6784 19525 6816
rect 19557 6784 19565 6816
rect 19597 6784 19605 6816
rect 19637 6784 19645 6816
rect 19677 6784 19680 6816
rect 19522 6783 19680 6784
rect 57621 6816 57779 6816
rect 57621 6784 57624 6816
rect 57656 6784 57664 6816
rect 57696 6784 57704 6816
rect 57736 6784 57744 6816
rect 57776 6784 57779 6816
rect 57621 6783 57779 6784
rect 95720 6816 95878 6816
rect 95720 6784 95723 6816
rect 95755 6784 95763 6816
rect 95795 6784 95803 6816
rect 95835 6784 95843 6816
rect 95875 6784 95878 6816
rect 95720 6783 95878 6784
rect 133819 6816 133977 6816
rect 133819 6784 133822 6816
rect 133854 6784 133862 6816
rect 133894 6784 133902 6816
rect 133934 6784 133942 6816
rect 133974 6784 133977 6816
rect 133819 6783 133977 6784
rect 103552 6781 103585 6782
rect 104012 6781 104045 6782
rect 103552 6780 104045 6781
rect 103552 6752 103555 6780
rect 103583 6752 104015 6780
rect 104043 6752 104045 6780
rect 103552 6751 104045 6752
rect 103552 6749 103585 6751
rect 104012 6749 104045 6751
rect 106634 6713 106667 6714
rect 109900 6713 109933 6714
rect 106634 6712 109933 6713
rect 106634 6684 106637 6712
rect 106665 6684 109903 6712
rect 109931 6684 109933 6712
rect 106634 6683 109933 6684
rect 106634 6681 106667 6683
rect 109900 6681 109933 6683
rect 113534 6713 113567 6714
rect 114592 6713 114625 6714
rect 113534 6712 114625 6713
rect 113534 6684 113537 6712
rect 113565 6684 114595 6712
rect 114623 6684 114625 6712
rect 113534 6683 114625 6684
rect 113534 6681 113567 6683
rect 114592 6681 114625 6683
rect 119054 6713 119087 6714
rect 119744 6713 119777 6714
rect 119054 6712 119777 6713
rect 119054 6684 119057 6712
rect 119085 6684 119747 6712
rect 119775 6684 119777 6712
rect 119054 6683 119777 6684
rect 119054 6681 119087 6683
rect 119744 6681 119777 6683
rect 134464 6713 134497 6714
rect 136580 6713 136613 6714
rect 134464 6712 136613 6713
rect 134464 6684 134467 6712
rect 134495 6684 136583 6712
rect 136611 6684 136613 6712
rect 134464 6683 136613 6684
rect 134464 6681 134497 6683
rect 136580 6681 136613 6683
rect 100424 6645 100457 6646
rect 101712 6645 101745 6646
rect 100424 6644 101745 6645
rect 100424 6616 100427 6644
rect 100455 6616 101715 6644
rect 101743 6616 101745 6644
rect 100424 6615 101745 6616
rect 100424 6613 100457 6615
rect 101712 6613 101745 6615
rect 102770 6645 102803 6646
rect 102862 6645 102895 6646
rect 102770 6644 102895 6645
rect 102770 6616 102773 6644
rect 102801 6616 102865 6644
rect 102893 6616 102895 6644
rect 102770 6615 102895 6616
rect 102770 6613 102803 6615
rect 102862 6613 102895 6615
rect 103598 6645 103631 6646
rect 103966 6645 103999 6646
rect 103598 6644 103999 6645
rect 103598 6616 103601 6644
rect 103629 6616 103969 6644
rect 103997 6616 103999 6644
rect 103598 6615 103999 6616
rect 103598 6613 103631 6615
rect 103966 6613 103999 6615
rect 115190 6645 115223 6646
rect 116064 6645 116097 6646
rect 115190 6644 116097 6645
rect 115190 6616 115193 6644
rect 115221 6616 116067 6644
rect 116095 6616 116097 6644
rect 115190 6615 116097 6616
rect 115190 6613 115223 6615
rect 116064 6613 116097 6615
rect 131704 6645 131737 6646
rect 132762 6645 132795 6646
rect 131704 6644 132795 6645
rect 131704 6616 131707 6644
rect 131735 6616 132765 6644
rect 132793 6616 132795 6644
rect 131704 6615 132795 6616
rect 131704 6613 131737 6615
rect 132762 6613 132795 6615
rect 134510 6645 134543 6646
rect 136626 6645 136659 6646
rect 134510 6644 136659 6645
rect 134510 6616 134513 6644
rect 134541 6616 136629 6644
rect 136657 6616 136659 6644
rect 134510 6615 136659 6616
rect 134510 6613 134543 6615
rect 136626 6613 136659 6615
rect 43476 6577 43509 6578
rect 45914 6577 45947 6578
rect 43476 6576 45947 6577
rect 43476 6548 43479 6576
rect 43507 6548 45917 6576
rect 45945 6548 45947 6576
rect 43476 6547 45947 6548
rect 43476 6545 43509 6547
rect 45914 6545 45947 6547
rect 112706 6577 112739 6578
rect 113534 6577 113567 6578
rect 112706 6576 113567 6577
rect 112706 6548 112709 6576
rect 112737 6548 113537 6576
rect 113565 6548 113567 6576
rect 112706 6547 113567 6548
rect 112706 6545 112739 6547
rect 113534 6545 113567 6547
rect 38572 6544 38730 6544
rect 38572 6512 38575 6544
rect 38607 6512 38615 6544
rect 38647 6512 38655 6544
rect 38687 6512 38695 6544
rect 38727 6512 38730 6544
rect 38572 6511 38730 6512
rect 76671 6544 76829 6544
rect 76671 6512 76674 6544
rect 76706 6512 76714 6544
rect 76746 6512 76754 6544
rect 76786 6512 76794 6544
rect 76826 6512 76829 6544
rect 76671 6511 76829 6512
rect 114770 6544 114928 6544
rect 114770 6512 114773 6544
rect 114805 6512 114813 6544
rect 114845 6512 114853 6544
rect 114885 6512 114893 6544
rect 114925 6512 114928 6544
rect 114770 6511 114928 6512
rect 128300 6509 128333 6510
rect 128990 6509 129023 6510
rect 128300 6508 129023 6509
rect 128300 6480 128303 6508
rect 128331 6480 128993 6508
rect 129021 6480 129023 6508
rect 128300 6479 129023 6480
rect 128300 6477 128333 6479
rect 128990 6477 129023 6479
rect 77516 6441 77549 6442
rect 97296 6441 97329 6442
rect 97894 6441 97927 6442
rect 77516 6440 97927 6441
rect 77516 6412 77519 6440
rect 77547 6412 97299 6440
rect 97327 6412 97897 6440
rect 97925 6412 97927 6440
rect 77516 6411 97927 6412
rect 77516 6409 77549 6411
rect 97296 6409 97329 6411
rect 97894 6409 97927 6411
rect 98676 6441 98709 6442
rect 149736 6441 149769 6442
rect 98676 6440 149769 6441
rect 98676 6412 98679 6440
rect 98707 6412 149739 6440
rect 149767 6412 149769 6440
rect 98676 6411 149769 6412
rect 98676 6409 98709 6411
rect 149736 6409 149769 6411
rect 43890 6373 43923 6374
rect 45362 6373 45395 6374
rect 43890 6372 45395 6373
rect 43890 6344 43893 6372
rect 43921 6344 45365 6372
rect 45393 6344 45395 6372
rect 43890 6343 45395 6344
rect 43890 6341 43923 6343
rect 45362 6341 45395 6343
rect 97526 6373 97559 6374
rect 103920 6373 103953 6374
rect 97526 6372 103953 6373
rect 97526 6344 97529 6372
rect 97557 6344 103923 6372
rect 103951 6344 103953 6372
rect 97526 6343 103953 6344
rect 97526 6341 97559 6343
rect 103920 6341 103953 6343
rect 119146 6373 119179 6374
rect 121078 6373 121111 6374
rect 119146 6372 121111 6373
rect 119146 6344 119149 6372
rect 119177 6344 121081 6372
rect 121109 6344 121111 6372
rect 119146 6343 121111 6344
rect 119146 6341 119179 6343
rect 121078 6341 121111 6343
rect 131152 6373 131185 6374
rect 131750 6373 131783 6374
rect 131152 6372 131783 6373
rect 131152 6344 131155 6372
rect 131183 6344 131753 6372
rect 131781 6344 131783 6372
rect 131152 6343 131783 6344
rect 131152 6341 131185 6343
rect 131750 6341 131783 6343
rect 132164 6373 132197 6374
rect 133544 6373 133577 6374
rect 132164 6372 133577 6373
rect 132164 6344 132167 6372
rect 132195 6344 133547 6372
rect 133575 6344 133577 6372
rect 132164 6343 133577 6344
rect 132164 6341 132197 6343
rect 133544 6341 133577 6343
rect 133820 6373 133853 6374
rect 134050 6373 134083 6374
rect 133820 6372 134083 6373
rect 133820 6344 133823 6372
rect 133851 6344 134053 6372
rect 134081 6344 134083 6372
rect 133820 6343 134083 6344
rect 133820 6341 133853 6343
rect 134050 6341 134083 6343
rect 78942 6305 78975 6306
rect 80138 6305 80171 6306
rect 78942 6304 80171 6305
rect 78942 6276 78945 6304
rect 78973 6276 80141 6304
rect 80169 6276 80171 6304
rect 78942 6275 80171 6276
rect 78942 6273 78975 6275
rect 80138 6273 80171 6275
rect 95916 6305 95949 6306
rect 96100 6305 96133 6306
rect 95916 6304 96133 6305
rect 95916 6276 95919 6304
rect 95947 6276 96103 6304
rect 96131 6276 96133 6304
rect 95916 6275 96133 6276
rect 95916 6273 95949 6275
rect 96100 6273 96133 6275
rect 100194 6305 100227 6306
rect 102632 6305 102665 6306
rect 100194 6304 102665 6305
rect 100194 6276 100197 6304
rect 100225 6276 102635 6304
rect 102663 6276 102665 6304
rect 100194 6275 102665 6276
rect 100194 6273 100227 6275
rect 102632 6273 102665 6275
rect 125954 6305 125987 6306
rect 128530 6305 128563 6306
rect 125954 6304 128563 6305
rect 125954 6276 125957 6304
rect 125985 6276 128533 6304
rect 128561 6276 128563 6304
rect 125954 6275 128563 6276
rect 125954 6273 125987 6275
rect 128530 6273 128563 6275
rect 19522 6272 19680 6272
rect 19522 6240 19525 6272
rect 19557 6240 19565 6272
rect 19597 6240 19605 6272
rect 19637 6240 19645 6272
rect 19677 6240 19680 6272
rect 19522 6239 19680 6240
rect 57621 6272 57779 6272
rect 57621 6240 57624 6272
rect 57656 6240 57664 6272
rect 57696 6240 57704 6272
rect 57736 6240 57744 6272
rect 57776 6240 57779 6272
rect 57621 6239 57779 6240
rect 95720 6272 95878 6272
rect 95720 6240 95723 6272
rect 95755 6240 95763 6272
rect 95795 6240 95803 6272
rect 95835 6240 95843 6272
rect 95875 6240 95878 6272
rect 95720 6239 95878 6240
rect 133819 6272 133977 6272
rect 133819 6240 133822 6272
rect 133854 6240 133862 6272
rect 133894 6240 133902 6272
rect 133934 6240 133942 6272
rect 133974 6240 133977 6272
rect 133819 6239 133977 6240
rect 125908 6237 125941 6238
rect 128576 6237 128609 6238
rect 125908 6236 128609 6237
rect 125908 6208 125911 6236
rect 125939 6208 128579 6236
rect 128607 6208 128609 6236
rect 125908 6207 128609 6208
rect 125908 6205 125941 6207
rect 128576 6205 128609 6207
rect 44074 6169 44107 6170
rect 44948 6169 44981 6170
rect 44074 6168 44981 6169
rect 44074 6140 44077 6168
rect 44105 6140 44951 6168
rect 44979 6140 44981 6168
rect 44074 6139 44981 6140
rect 44074 6137 44107 6139
rect 44948 6137 44981 6139
rect 81794 6169 81827 6170
rect 96514 6169 96547 6170
rect 81794 6168 96547 6169
rect 81794 6140 81797 6168
rect 81825 6140 96517 6168
rect 96545 6140 96547 6168
rect 81794 6139 96547 6140
rect 81794 6137 81827 6139
rect 96514 6137 96547 6139
rect 14680 6101 14713 6102
rect 15370 6101 15403 6102
rect 15692 6101 15725 6102
rect 14680 6100 15725 6101
rect 14680 6072 14683 6100
rect 14711 6072 15373 6100
rect 15401 6072 15695 6100
rect 15723 6072 15725 6100
rect 14680 6071 15725 6072
rect 14680 6069 14713 6071
rect 15370 6069 15403 6071
rect 15692 6069 15725 6071
rect 20292 6101 20325 6102
rect 21212 6101 21245 6102
rect 20292 6100 21245 6101
rect 20292 6072 20295 6100
rect 20323 6072 21215 6100
rect 21243 6072 21245 6100
rect 20292 6071 21245 6072
rect 20292 6069 20325 6071
rect 21212 6069 21245 6071
rect 38572 6000 38730 6000
rect 38572 5968 38575 6000
rect 38607 5968 38615 6000
rect 38647 5968 38655 6000
rect 38687 5968 38695 6000
rect 38727 5968 38730 6000
rect 38572 5967 38730 5968
rect 76671 6000 76829 6000
rect 76671 5968 76674 6000
rect 76706 5968 76714 6000
rect 76746 5968 76754 6000
rect 76786 5968 76794 6000
rect 76826 5968 76829 6000
rect 76671 5967 76829 5968
rect 114770 6000 114928 6000
rect 114770 5968 114773 6000
rect 114805 5968 114813 6000
rect 114845 5968 114853 6000
rect 114885 5968 114893 6000
rect 114925 5968 114928 6000
rect 114770 5967 114928 5968
rect 94812 5897 94845 5898
rect 96514 5897 96547 5898
rect 94812 5896 96547 5897
rect 94812 5868 94815 5896
rect 94843 5868 96517 5896
rect 96545 5868 96547 5896
rect 94812 5867 96547 5868
rect 94812 5865 94845 5867
rect 96514 5865 96547 5867
rect 19522 5728 19680 5728
rect 19522 5696 19525 5728
rect 19557 5696 19565 5728
rect 19597 5696 19605 5728
rect 19637 5696 19645 5728
rect 19677 5696 19680 5728
rect 19522 5695 19680 5696
rect 57621 5728 57779 5728
rect 57621 5696 57624 5728
rect 57656 5696 57664 5728
rect 57696 5696 57704 5728
rect 57736 5696 57744 5728
rect 57776 5696 57779 5728
rect 57621 5695 57779 5696
rect 95720 5728 95878 5728
rect 95720 5696 95723 5728
rect 95755 5696 95763 5728
rect 95795 5696 95803 5728
rect 95835 5696 95843 5728
rect 95875 5696 95878 5728
rect 95720 5695 95878 5696
rect 133819 5728 133977 5728
rect 133819 5696 133822 5728
rect 133854 5696 133862 5728
rect 133894 5696 133902 5728
rect 133934 5696 133942 5728
rect 133974 5696 133977 5728
rect 133819 5695 133977 5696
rect 38572 5456 38730 5456
rect 38572 5424 38575 5456
rect 38607 5424 38615 5456
rect 38647 5424 38655 5456
rect 38687 5424 38695 5456
rect 38727 5424 38730 5456
rect 38572 5423 38730 5424
rect 76671 5456 76829 5456
rect 76671 5424 76674 5456
rect 76706 5424 76714 5456
rect 76746 5424 76754 5456
rect 76786 5424 76794 5456
rect 76826 5424 76829 5456
rect 76671 5423 76829 5424
rect 114770 5456 114928 5456
rect 114770 5424 114773 5456
rect 114805 5424 114813 5456
rect 114845 5424 114853 5456
rect 114885 5424 114893 5456
rect 114925 5424 114928 5456
rect 114770 5423 114928 5424
rect 19522 5184 19680 5184
rect 19522 5152 19525 5184
rect 19557 5152 19565 5184
rect 19597 5152 19605 5184
rect 19637 5152 19645 5184
rect 19677 5152 19680 5184
rect 19522 5151 19680 5152
rect 57621 5184 57779 5184
rect 57621 5152 57624 5184
rect 57656 5152 57664 5184
rect 57696 5152 57704 5184
rect 57736 5152 57744 5184
rect 57776 5152 57779 5184
rect 57621 5151 57779 5152
rect 95720 5184 95878 5184
rect 95720 5152 95723 5184
rect 95755 5152 95763 5184
rect 95795 5152 95803 5184
rect 95835 5152 95843 5184
rect 95875 5152 95878 5184
rect 95720 5151 95878 5152
rect 133819 5184 133977 5184
rect 133819 5152 133822 5184
rect 133854 5152 133862 5184
rect 133894 5152 133902 5184
rect 133934 5152 133942 5184
rect 133974 5152 133977 5184
rect 133819 5151 133977 5152
rect 152220 5013 152253 5014
rect 153100 5013 153500 5028
rect 152220 5012 153500 5013
rect 152220 4984 152223 5012
rect 152251 4984 153500 5012
rect 152220 4983 153500 4984
rect 152220 4981 152253 4983
rect 153100 4968 153500 4983
rect 38572 4912 38730 4912
rect 38572 4880 38575 4912
rect 38607 4880 38615 4912
rect 38647 4880 38655 4912
rect 38687 4880 38695 4912
rect 38727 4880 38730 4912
rect 38572 4879 38730 4880
rect 76671 4912 76829 4912
rect 76671 4880 76674 4912
rect 76706 4880 76714 4912
rect 76746 4880 76754 4912
rect 76786 4880 76794 4912
rect 76826 4880 76829 4912
rect 76671 4879 76829 4880
rect 114770 4912 114928 4912
rect 114770 4880 114773 4912
rect 114805 4880 114813 4912
rect 114845 4880 114853 4912
rect 114885 4880 114893 4912
rect 114925 4880 114928 4912
rect 114770 4879 114928 4880
rect 19522 4640 19680 4640
rect 19522 4608 19525 4640
rect 19557 4608 19565 4640
rect 19597 4608 19605 4640
rect 19637 4608 19645 4640
rect 19677 4608 19680 4640
rect 19522 4607 19680 4608
rect 57621 4640 57779 4640
rect 57621 4608 57624 4640
rect 57656 4608 57664 4640
rect 57696 4608 57704 4640
rect 57736 4608 57744 4640
rect 57776 4608 57779 4640
rect 57621 4607 57779 4608
rect 95720 4640 95878 4640
rect 95720 4608 95723 4640
rect 95755 4608 95763 4640
rect 95795 4608 95803 4640
rect 95835 4608 95843 4640
rect 95875 4608 95878 4640
rect 95720 4607 95878 4608
rect 133819 4640 133977 4640
rect 133819 4608 133822 4640
rect 133854 4608 133862 4640
rect 133894 4608 133902 4640
rect 133934 4608 133942 4640
rect 133974 4608 133977 4640
rect 133819 4607 133977 4608
rect 38572 4368 38730 4368
rect 38572 4336 38575 4368
rect 38607 4336 38615 4368
rect 38647 4336 38655 4368
rect 38687 4336 38695 4368
rect 38727 4336 38730 4368
rect 38572 4335 38730 4336
rect 76671 4368 76829 4368
rect 76671 4336 76674 4368
rect 76706 4336 76714 4368
rect 76746 4336 76754 4368
rect 76786 4336 76794 4368
rect 76826 4336 76829 4368
rect 76671 4335 76829 4336
rect 114770 4368 114928 4368
rect 114770 4336 114773 4368
rect 114805 4336 114813 4368
rect 114845 4336 114853 4368
rect 114885 4336 114893 4368
rect 114925 4336 114928 4368
rect 114770 4335 114928 4336
rect 19522 4096 19680 4096
rect 0 4061 400 4076
rect 19522 4064 19525 4096
rect 19557 4064 19565 4096
rect 19597 4064 19605 4096
rect 19637 4064 19645 4096
rect 19677 4064 19680 4096
rect 19522 4063 19680 4064
rect 57621 4096 57779 4096
rect 57621 4064 57624 4096
rect 57656 4064 57664 4096
rect 57696 4064 57704 4096
rect 57736 4064 57744 4096
rect 57776 4064 57779 4096
rect 57621 4063 57779 4064
rect 95720 4096 95878 4096
rect 95720 4064 95723 4096
rect 95755 4064 95763 4096
rect 95795 4064 95803 4096
rect 95835 4064 95843 4096
rect 95875 4064 95878 4096
rect 95720 4063 95878 4064
rect 133819 4096 133977 4096
rect 133819 4064 133822 4096
rect 133854 4064 133862 4096
rect 133894 4064 133902 4096
rect 133934 4064 133942 4096
rect 133974 4064 133977 4096
rect 133819 4063 133977 4064
rect 696 4061 729 4062
rect 0 4060 729 4061
rect 0 4032 699 4060
rect 727 4032 729 4060
rect 0 4031 729 4032
rect 0 4016 400 4031
rect 696 4029 729 4031
rect 38572 3824 38730 3824
rect 38572 3792 38575 3824
rect 38607 3792 38615 3824
rect 38647 3792 38655 3824
rect 38687 3792 38695 3824
rect 38727 3792 38730 3824
rect 38572 3791 38730 3792
rect 76671 3824 76829 3824
rect 76671 3792 76674 3824
rect 76706 3792 76714 3824
rect 76746 3792 76754 3824
rect 76786 3792 76794 3824
rect 76826 3792 76829 3824
rect 76671 3791 76829 3792
rect 114770 3824 114928 3824
rect 114770 3792 114773 3824
rect 114805 3792 114813 3824
rect 114845 3792 114853 3824
rect 114885 3792 114893 3824
rect 114925 3792 114928 3824
rect 114770 3791 114928 3792
rect 19522 3552 19680 3552
rect 19522 3520 19525 3552
rect 19557 3520 19565 3552
rect 19597 3520 19605 3552
rect 19637 3520 19645 3552
rect 19677 3520 19680 3552
rect 19522 3519 19680 3520
rect 57621 3552 57779 3552
rect 57621 3520 57624 3552
rect 57656 3520 57664 3552
rect 57696 3520 57704 3552
rect 57736 3520 57744 3552
rect 57776 3520 57779 3552
rect 57621 3519 57779 3520
rect 95720 3552 95878 3552
rect 95720 3520 95723 3552
rect 95755 3520 95763 3552
rect 95795 3520 95803 3552
rect 95835 3520 95843 3552
rect 95875 3520 95878 3552
rect 95720 3519 95878 3520
rect 133819 3552 133977 3552
rect 133819 3520 133822 3552
rect 133854 3520 133862 3552
rect 133894 3520 133902 3552
rect 133934 3520 133942 3552
rect 133974 3520 133977 3552
rect 133819 3519 133977 3520
rect 38572 3280 38730 3280
rect 38572 3248 38575 3280
rect 38607 3248 38615 3280
rect 38647 3248 38655 3280
rect 38687 3248 38695 3280
rect 38727 3248 38730 3280
rect 38572 3247 38730 3248
rect 76671 3280 76829 3280
rect 76671 3248 76674 3280
rect 76706 3248 76714 3280
rect 76746 3248 76754 3280
rect 76786 3248 76794 3280
rect 76826 3248 76829 3280
rect 76671 3247 76829 3248
rect 114770 3280 114928 3280
rect 114770 3248 114773 3280
rect 114805 3248 114813 3280
rect 114845 3248 114853 3280
rect 114885 3248 114893 3280
rect 114925 3248 114928 3280
rect 114770 3247 114928 3248
rect 19522 3008 19680 3008
rect 19522 2976 19525 3008
rect 19557 2976 19565 3008
rect 19597 2976 19605 3008
rect 19637 2976 19645 3008
rect 19677 2976 19680 3008
rect 19522 2975 19680 2976
rect 57621 3008 57779 3008
rect 57621 2976 57624 3008
rect 57656 2976 57664 3008
rect 57696 2976 57704 3008
rect 57736 2976 57744 3008
rect 57776 2976 57779 3008
rect 57621 2975 57779 2976
rect 95720 3008 95878 3008
rect 95720 2976 95723 3008
rect 95755 2976 95763 3008
rect 95795 2976 95803 3008
rect 95835 2976 95843 3008
rect 95875 2976 95878 3008
rect 95720 2975 95878 2976
rect 133819 3008 133977 3008
rect 133819 2976 133822 3008
rect 133854 2976 133862 3008
rect 133894 2976 133902 3008
rect 133934 2976 133942 3008
rect 133974 2976 133977 3008
rect 133819 2975 133977 2976
rect 151990 2973 152023 2974
rect 153100 2973 153500 2988
rect 151990 2972 153500 2973
rect 151990 2944 151993 2972
rect 152021 2944 153500 2972
rect 151990 2943 153500 2944
rect 151990 2941 152023 2943
rect 153100 2928 153500 2943
rect 38572 2736 38730 2736
rect 38572 2704 38575 2736
rect 38607 2704 38615 2736
rect 38647 2704 38655 2736
rect 38687 2704 38695 2736
rect 38727 2704 38730 2736
rect 38572 2703 38730 2704
rect 76671 2736 76829 2736
rect 76671 2704 76674 2736
rect 76706 2704 76714 2736
rect 76746 2704 76754 2736
rect 76786 2704 76794 2736
rect 76826 2704 76829 2736
rect 76671 2703 76829 2704
rect 114770 2736 114928 2736
rect 114770 2704 114773 2736
rect 114805 2704 114813 2736
rect 114845 2704 114853 2736
rect 114885 2704 114893 2736
rect 114925 2704 114928 2736
rect 114770 2703 114928 2704
rect 19522 2464 19680 2464
rect 19522 2432 19525 2464
rect 19557 2432 19565 2464
rect 19597 2432 19605 2464
rect 19637 2432 19645 2464
rect 19677 2432 19680 2464
rect 19522 2431 19680 2432
rect 57621 2464 57779 2464
rect 57621 2432 57624 2464
rect 57656 2432 57664 2464
rect 57696 2432 57704 2464
rect 57736 2432 57744 2464
rect 57776 2432 57779 2464
rect 57621 2431 57779 2432
rect 95720 2464 95878 2464
rect 95720 2432 95723 2464
rect 95755 2432 95763 2464
rect 95795 2432 95803 2464
rect 95835 2432 95843 2464
rect 95875 2432 95878 2464
rect 95720 2431 95878 2432
rect 133819 2464 133977 2464
rect 133819 2432 133822 2464
rect 133854 2432 133862 2464
rect 133894 2432 133902 2464
rect 133934 2432 133942 2464
rect 133974 2432 133977 2464
rect 133819 2431 133977 2432
rect 38572 2192 38730 2192
rect 38572 2160 38575 2192
rect 38607 2160 38615 2192
rect 38647 2160 38655 2192
rect 38687 2160 38695 2192
rect 38727 2160 38730 2192
rect 38572 2159 38730 2160
rect 76671 2192 76829 2192
rect 76671 2160 76674 2192
rect 76706 2160 76714 2192
rect 76746 2160 76754 2192
rect 76786 2160 76794 2192
rect 76826 2160 76829 2192
rect 76671 2159 76829 2160
rect 114770 2192 114928 2192
rect 114770 2160 114773 2192
rect 114805 2160 114813 2192
rect 114845 2160 114853 2192
rect 114885 2160 114893 2192
rect 114925 2160 114928 2192
rect 114770 2159 114928 2160
rect 19522 1920 19680 1920
rect 19522 1888 19525 1920
rect 19557 1888 19565 1920
rect 19597 1888 19605 1920
rect 19637 1888 19645 1920
rect 19677 1888 19680 1920
rect 19522 1887 19680 1888
rect 57621 1920 57779 1920
rect 57621 1888 57624 1920
rect 57656 1888 57664 1920
rect 57696 1888 57704 1920
rect 57736 1888 57744 1920
rect 57776 1888 57779 1920
rect 57621 1887 57779 1888
rect 95720 1920 95878 1920
rect 95720 1888 95723 1920
rect 95755 1888 95763 1920
rect 95795 1888 95803 1920
rect 95835 1888 95843 1920
rect 95875 1888 95878 1920
rect 95720 1887 95878 1888
rect 133819 1920 133977 1920
rect 133819 1888 133822 1920
rect 133854 1888 133862 1920
rect 133894 1888 133902 1920
rect 133934 1888 133942 1920
rect 133974 1888 133977 1920
rect 133819 1887 133977 1888
rect 38572 1648 38730 1648
rect 38572 1616 38575 1648
rect 38607 1616 38615 1648
rect 38647 1616 38655 1648
rect 38687 1616 38695 1648
rect 38727 1616 38730 1648
rect 38572 1615 38730 1616
rect 76671 1648 76829 1648
rect 76671 1616 76674 1648
rect 76706 1616 76714 1648
rect 76746 1616 76754 1648
rect 76786 1616 76794 1648
rect 76826 1616 76829 1648
rect 76671 1615 76829 1616
rect 114770 1648 114928 1648
rect 114770 1616 114773 1648
rect 114805 1616 114813 1648
rect 114845 1616 114853 1648
rect 114885 1616 114893 1648
rect 114925 1616 114928 1648
rect 114770 1615 114928 1616
rect 19522 1376 19680 1376
rect 19522 1344 19525 1376
rect 19557 1344 19565 1376
rect 19597 1344 19605 1376
rect 19637 1344 19645 1376
rect 19677 1344 19680 1376
rect 19522 1343 19680 1344
rect 57621 1376 57779 1376
rect 57621 1344 57624 1376
rect 57656 1344 57664 1376
rect 57696 1344 57704 1376
rect 57736 1344 57744 1376
rect 57776 1344 57779 1376
rect 57621 1343 57779 1344
rect 95720 1376 95878 1376
rect 95720 1344 95723 1376
rect 95755 1344 95763 1376
rect 95795 1344 95803 1376
rect 95835 1344 95843 1376
rect 95875 1344 95878 1376
rect 95720 1343 95878 1344
rect 133819 1376 133977 1376
rect 133819 1344 133822 1376
rect 133854 1344 133862 1376
rect 133894 1344 133902 1376
rect 133934 1344 133942 1376
rect 133974 1344 133977 1376
rect 133819 1343 133977 1344
rect 38572 1104 38730 1104
rect 38572 1072 38575 1104
rect 38607 1072 38615 1104
rect 38647 1072 38655 1104
rect 38687 1072 38695 1104
rect 38727 1072 38730 1104
rect 38572 1071 38730 1072
rect 76671 1104 76829 1104
rect 76671 1072 76674 1104
rect 76706 1072 76714 1104
rect 76746 1072 76754 1104
rect 76786 1072 76794 1104
rect 76826 1072 76829 1104
rect 76671 1071 76829 1072
rect 114770 1104 114928 1104
rect 114770 1072 114773 1104
rect 114805 1072 114813 1104
rect 114845 1072 114853 1104
rect 114885 1072 114893 1104
rect 114925 1072 114928 1104
rect 114770 1071 114928 1072
rect 151116 1001 151149 1002
rect 153100 1001 153500 1016
rect 151116 1000 153500 1001
rect 151116 972 151119 1000
rect 151147 972 153500 1000
rect 151116 971 153500 972
rect 151116 969 151149 971
rect 153100 956 153500 971
<< via3 >>
rect 19525 6814 19557 6816
rect 19525 6786 19527 6814
rect 19527 6786 19555 6814
rect 19555 6786 19557 6814
rect 19525 6784 19557 6786
rect 19565 6814 19597 6816
rect 19565 6786 19567 6814
rect 19567 6786 19595 6814
rect 19595 6786 19597 6814
rect 19565 6784 19597 6786
rect 19605 6814 19637 6816
rect 19605 6786 19607 6814
rect 19607 6786 19635 6814
rect 19635 6786 19637 6814
rect 19605 6784 19637 6786
rect 19645 6814 19677 6816
rect 19645 6786 19647 6814
rect 19647 6786 19675 6814
rect 19675 6786 19677 6814
rect 19645 6784 19677 6786
rect 57624 6814 57656 6816
rect 57624 6786 57626 6814
rect 57626 6786 57654 6814
rect 57654 6786 57656 6814
rect 57624 6784 57656 6786
rect 57664 6814 57696 6816
rect 57664 6786 57666 6814
rect 57666 6786 57694 6814
rect 57694 6786 57696 6814
rect 57664 6784 57696 6786
rect 57704 6814 57736 6816
rect 57704 6786 57706 6814
rect 57706 6786 57734 6814
rect 57734 6786 57736 6814
rect 57704 6784 57736 6786
rect 57744 6814 57776 6816
rect 57744 6786 57746 6814
rect 57746 6786 57774 6814
rect 57774 6786 57776 6814
rect 57744 6784 57776 6786
rect 95723 6814 95755 6816
rect 95723 6786 95725 6814
rect 95725 6786 95753 6814
rect 95753 6786 95755 6814
rect 95723 6784 95755 6786
rect 95763 6814 95795 6816
rect 95763 6786 95765 6814
rect 95765 6786 95793 6814
rect 95793 6786 95795 6814
rect 95763 6784 95795 6786
rect 95803 6814 95835 6816
rect 95803 6786 95805 6814
rect 95805 6786 95833 6814
rect 95833 6786 95835 6814
rect 95803 6784 95835 6786
rect 95843 6814 95875 6816
rect 95843 6786 95845 6814
rect 95845 6786 95873 6814
rect 95873 6786 95875 6814
rect 95843 6784 95875 6786
rect 133822 6814 133854 6816
rect 133822 6786 133824 6814
rect 133824 6786 133852 6814
rect 133852 6786 133854 6814
rect 133822 6784 133854 6786
rect 133862 6814 133894 6816
rect 133862 6786 133864 6814
rect 133864 6786 133892 6814
rect 133892 6786 133894 6814
rect 133862 6784 133894 6786
rect 133902 6814 133934 6816
rect 133902 6786 133904 6814
rect 133904 6786 133932 6814
rect 133932 6786 133934 6814
rect 133902 6784 133934 6786
rect 133942 6814 133974 6816
rect 133942 6786 133944 6814
rect 133944 6786 133972 6814
rect 133972 6786 133974 6814
rect 133942 6784 133974 6786
rect 38575 6542 38607 6544
rect 38575 6514 38577 6542
rect 38577 6514 38605 6542
rect 38605 6514 38607 6542
rect 38575 6512 38607 6514
rect 38615 6542 38647 6544
rect 38615 6514 38617 6542
rect 38617 6514 38645 6542
rect 38645 6514 38647 6542
rect 38615 6512 38647 6514
rect 38655 6542 38687 6544
rect 38655 6514 38657 6542
rect 38657 6514 38685 6542
rect 38685 6514 38687 6542
rect 38655 6512 38687 6514
rect 38695 6542 38727 6544
rect 38695 6514 38697 6542
rect 38697 6514 38725 6542
rect 38725 6514 38727 6542
rect 38695 6512 38727 6514
rect 76674 6542 76706 6544
rect 76674 6514 76676 6542
rect 76676 6514 76704 6542
rect 76704 6514 76706 6542
rect 76674 6512 76706 6514
rect 76714 6542 76746 6544
rect 76714 6514 76716 6542
rect 76716 6514 76744 6542
rect 76744 6514 76746 6542
rect 76714 6512 76746 6514
rect 76754 6542 76786 6544
rect 76754 6514 76756 6542
rect 76756 6514 76784 6542
rect 76784 6514 76786 6542
rect 76754 6512 76786 6514
rect 76794 6542 76826 6544
rect 76794 6514 76796 6542
rect 76796 6514 76824 6542
rect 76824 6514 76826 6542
rect 76794 6512 76826 6514
rect 114773 6542 114805 6544
rect 114773 6514 114775 6542
rect 114775 6514 114803 6542
rect 114803 6514 114805 6542
rect 114773 6512 114805 6514
rect 114813 6542 114845 6544
rect 114813 6514 114815 6542
rect 114815 6514 114843 6542
rect 114843 6514 114845 6542
rect 114813 6512 114845 6514
rect 114853 6542 114885 6544
rect 114853 6514 114855 6542
rect 114855 6514 114883 6542
rect 114883 6514 114885 6542
rect 114853 6512 114885 6514
rect 114893 6542 114925 6544
rect 114893 6514 114895 6542
rect 114895 6514 114923 6542
rect 114923 6514 114925 6542
rect 114893 6512 114925 6514
rect 19525 6270 19557 6272
rect 19525 6242 19527 6270
rect 19527 6242 19555 6270
rect 19555 6242 19557 6270
rect 19525 6240 19557 6242
rect 19565 6270 19597 6272
rect 19565 6242 19567 6270
rect 19567 6242 19595 6270
rect 19595 6242 19597 6270
rect 19565 6240 19597 6242
rect 19605 6270 19637 6272
rect 19605 6242 19607 6270
rect 19607 6242 19635 6270
rect 19635 6242 19637 6270
rect 19605 6240 19637 6242
rect 19645 6270 19677 6272
rect 19645 6242 19647 6270
rect 19647 6242 19675 6270
rect 19675 6242 19677 6270
rect 19645 6240 19677 6242
rect 57624 6270 57656 6272
rect 57624 6242 57626 6270
rect 57626 6242 57654 6270
rect 57654 6242 57656 6270
rect 57624 6240 57656 6242
rect 57664 6270 57696 6272
rect 57664 6242 57666 6270
rect 57666 6242 57694 6270
rect 57694 6242 57696 6270
rect 57664 6240 57696 6242
rect 57704 6270 57736 6272
rect 57704 6242 57706 6270
rect 57706 6242 57734 6270
rect 57734 6242 57736 6270
rect 57704 6240 57736 6242
rect 57744 6270 57776 6272
rect 57744 6242 57746 6270
rect 57746 6242 57774 6270
rect 57774 6242 57776 6270
rect 57744 6240 57776 6242
rect 95723 6270 95755 6272
rect 95723 6242 95725 6270
rect 95725 6242 95753 6270
rect 95753 6242 95755 6270
rect 95723 6240 95755 6242
rect 95763 6270 95795 6272
rect 95763 6242 95765 6270
rect 95765 6242 95793 6270
rect 95793 6242 95795 6270
rect 95763 6240 95795 6242
rect 95803 6270 95835 6272
rect 95803 6242 95805 6270
rect 95805 6242 95833 6270
rect 95833 6242 95835 6270
rect 95803 6240 95835 6242
rect 95843 6270 95875 6272
rect 95843 6242 95845 6270
rect 95845 6242 95873 6270
rect 95873 6242 95875 6270
rect 95843 6240 95875 6242
rect 133822 6270 133854 6272
rect 133822 6242 133824 6270
rect 133824 6242 133852 6270
rect 133852 6242 133854 6270
rect 133822 6240 133854 6242
rect 133862 6270 133894 6272
rect 133862 6242 133864 6270
rect 133864 6242 133892 6270
rect 133892 6242 133894 6270
rect 133862 6240 133894 6242
rect 133902 6270 133934 6272
rect 133902 6242 133904 6270
rect 133904 6242 133932 6270
rect 133932 6242 133934 6270
rect 133902 6240 133934 6242
rect 133942 6270 133974 6272
rect 133942 6242 133944 6270
rect 133944 6242 133972 6270
rect 133972 6242 133974 6270
rect 133942 6240 133974 6242
rect 38575 5998 38607 6000
rect 38575 5970 38577 5998
rect 38577 5970 38605 5998
rect 38605 5970 38607 5998
rect 38575 5968 38607 5970
rect 38615 5998 38647 6000
rect 38615 5970 38617 5998
rect 38617 5970 38645 5998
rect 38645 5970 38647 5998
rect 38615 5968 38647 5970
rect 38655 5998 38687 6000
rect 38655 5970 38657 5998
rect 38657 5970 38685 5998
rect 38685 5970 38687 5998
rect 38655 5968 38687 5970
rect 38695 5998 38727 6000
rect 38695 5970 38697 5998
rect 38697 5970 38725 5998
rect 38725 5970 38727 5998
rect 38695 5968 38727 5970
rect 76674 5998 76706 6000
rect 76674 5970 76676 5998
rect 76676 5970 76704 5998
rect 76704 5970 76706 5998
rect 76674 5968 76706 5970
rect 76714 5998 76746 6000
rect 76714 5970 76716 5998
rect 76716 5970 76744 5998
rect 76744 5970 76746 5998
rect 76714 5968 76746 5970
rect 76754 5998 76786 6000
rect 76754 5970 76756 5998
rect 76756 5970 76784 5998
rect 76784 5970 76786 5998
rect 76754 5968 76786 5970
rect 76794 5998 76826 6000
rect 76794 5970 76796 5998
rect 76796 5970 76824 5998
rect 76824 5970 76826 5998
rect 76794 5968 76826 5970
rect 114773 5998 114805 6000
rect 114773 5970 114775 5998
rect 114775 5970 114803 5998
rect 114803 5970 114805 5998
rect 114773 5968 114805 5970
rect 114813 5998 114845 6000
rect 114813 5970 114815 5998
rect 114815 5970 114843 5998
rect 114843 5970 114845 5998
rect 114813 5968 114845 5970
rect 114853 5998 114885 6000
rect 114853 5970 114855 5998
rect 114855 5970 114883 5998
rect 114883 5970 114885 5998
rect 114853 5968 114885 5970
rect 114893 5998 114925 6000
rect 114893 5970 114895 5998
rect 114895 5970 114923 5998
rect 114923 5970 114925 5998
rect 114893 5968 114925 5970
rect 19525 5726 19557 5728
rect 19525 5698 19527 5726
rect 19527 5698 19555 5726
rect 19555 5698 19557 5726
rect 19525 5696 19557 5698
rect 19565 5726 19597 5728
rect 19565 5698 19567 5726
rect 19567 5698 19595 5726
rect 19595 5698 19597 5726
rect 19565 5696 19597 5698
rect 19605 5726 19637 5728
rect 19605 5698 19607 5726
rect 19607 5698 19635 5726
rect 19635 5698 19637 5726
rect 19605 5696 19637 5698
rect 19645 5726 19677 5728
rect 19645 5698 19647 5726
rect 19647 5698 19675 5726
rect 19675 5698 19677 5726
rect 19645 5696 19677 5698
rect 57624 5726 57656 5728
rect 57624 5698 57626 5726
rect 57626 5698 57654 5726
rect 57654 5698 57656 5726
rect 57624 5696 57656 5698
rect 57664 5726 57696 5728
rect 57664 5698 57666 5726
rect 57666 5698 57694 5726
rect 57694 5698 57696 5726
rect 57664 5696 57696 5698
rect 57704 5726 57736 5728
rect 57704 5698 57706 5726
rect 57706 5698 57734 5726
rect 57734 5698 57736 5726
rect 57704 5696 57736 5698
rect 57744 5726 57776 5728
rect 57744 5698 57746 5726
rect 57746 5698 57774 5726
rect 57774 5698 57776 5726
rect 57744 5696 57776 5698
rect 95723 5726 95755 5728
rect 95723 5698 95725 5726
rect 95725 5698 95753 5726
rect 95753 5698 95755 5726
rect 95723 5696 95755 5698
rect 95763 5726 95795 5728
rect 95763 5698 95765 5726
rect 95765 5698 95793 5726
rect 95793 5698 95795 5726
rect 95763 5696 95795 5698
rect 95803 5726 95835 5728
rect 95803 5698 95805 5726
rect 95805 5698 95833 5726
rect 95833 5698 95835 5726
rect 95803 5696 95835 5698
rect 95843 5726 95875 5728
rect 95843 5698 95845 5726
rect 95845 5698 95873 5726
rect 95873 5698 95875 5726
rect 95843 5696 95875 5698
rect 133822 5726 133854 5728
rect 133822 5698 133824 5726
rect 133824 5698 133852 5726
rect 133852 5698 133854 5726
rect 133822 5696 133854 5698
rect 133862 5726 133894 5728
rect 133862 5698 133864 5726
rect 133864 5698 133892 5726
rect 133892 5698 133894 5726
rect 133862 5696 133894 5698
rect 133902 5726 133934 5728
rect 133902 5698 133904 5726
rect 133904 5698 133932 5726
rect 133932 5698 133934 5726
rect 133902 5696 133934 5698
rect 133942 5726 133974 5728
rect 133942 5698 133944 5726
rect 133944 5698 133972 5726
rect 133972 5698 133974 5726
rect 133942 5696 133974 5698
rect 38575 5454 38607 5456
rect 38575 5426 38577 5454
rect 38577 5426 38605 5454
rect 38605 5426 38607 5454
rect 38575 5424 38607 5426
rect 38615 5454 38647 5456
rect 38615 5426 38617 5454
rect 38617 5426 38645 5454
rect 38645 5426 38647 5454
rect 38615 5424 38647 5426
rect 38655 5454 38687 5456
rect 38655 5426 38657 5454
rect 38657 5426 38685 5454
rect 38685 5426 38687 5454
rect 38655 5424 38687 5426
rect 38695 5454 38727 5456
rect 38695 5426 38697 5454
rect 38697 5426 38725 5454
rect 38725 5426 38727 5454
rect 38695 5424 38727 5426
rect 76674 5454 76706 5456
rect 76674 5426 76676 5454
rect 76676 5426 76704 5454
rect 76704 5426 76706 5454
rect 76674 5424 76706 5426
rect 76714 5454 76746 5456
rect 76714 5426 76716 5454
rect 76716 5426 76744 5454
rect 76744 5426 76746 5454
rect 76714 5424 76746 5426
rect 76754 5454 76786 5456
rect 76754 5426 76756 5454
rect 76756 5426 76784 5454
rect 76784 5426 76786 5454
rect 76754 5424 76786 5426
rect 76794 5454 76826 5456
rect 76794 5426 76796 5454
rect 76796 5426 76824 5454
rect 76824 5426 76826 5454
rect 76794 5424 76826 5426
rect 114773 5454 114805 5456
rect 114773 5426 114775 5454
rect 114775 5426 114803 5454
rect 114803 5426 114805 5454
rect 114773 5424 114805 5426
rect 114813 5454 114845 5456
rect 114813 5426 114815 5454
rect 114815 5426 114843 5454
rect 114843 5426 114845 5454
rect 114813 5424 114845 5426
rect 114853 5454 114885 5456
rect 114853 5426 114855 5454
rect 114855 5426 114883 5454
rect 114883 5426 114885 5454
rect 114853 5424 114885 5426
rect 114893 5454 114925 5456
rect 114893 5426 114895 5454
rect 114895 5426 114923 5454
rect 114923 5426 114925 5454
rect 114893 5424 114925 5426
rect 19525 5182 19557 5184
rect 19525 5154 19527 5182
rect 19527 5154 19555 5182
rect 19555 5154 19557 5182
rect 19525 5152 19557 5154
rect 19565 5182 19597 5184
rect 19565 5154 19567 5182
rect 19567 5154 19595 5182
rect 19595 5154 19597 5182
rect 19565 5152 19597 5154
rect 19605 5182 19637 5184
rect 19605 5154 19607 5182
rect 19607 5154 19635 5182
rect 19635 5154 19637 5182
rect 19605 5152 19637 5154
rect 19645 5182 19677 5184
rect 19645 5154 19647 5182
rect 19647 5154 19675 5182
rect 19675 5154 19677 5182
rect 19645 5152 19677 5154
rect 57624 5182 57656 5184
rect 57624 5154 57626 5182
rect 57626 5154 57654 5182
rect 57654 5154 57656 5182
rect 57624 5152 57656 5154
rect 57664 5182 57696 5184
rect 57664 5154 57666 5182
rect 57666 5154 57694 5182
rect 57694 5154 57696 5182
rect 57664 5152 57696 5154
rect 57704 5182 57736 5184
rect 57704 5154 57706 5182
rect 57706 5154 57734 5182
rect 57734 5154 57736 5182
rect 57704 5152 57736 5154
rect 57744 5182 57776 5184
rect 57744 5154 57746 5182
rect 57746 5154 57774 5182
rect 57774 5154 57776 5182
rect 57744 5152 57776 5154
rect 95723 5182 95755 5184
rect 95723 5154 95725 5182
rect 95725 5154 95753 5182
rect 95753 5154 95755 5182
rect 95723 5152 95755 5154
rect 95763 5182 95795 5184
rect 95763 5154 95765 5182
rect 95765 5154 95793 5182
rect 95793 5154 95795 5182
rect 95763 5152 95795 5154
rect 95803 5182 95835 5184
rect 95803 5154 95805 5182
rect 95805 5154 95833 5182
rect 95833 5154 95835 5182
rect 95803 5152 95835 5154
rect 95843 5182 95875 5184
rect 95843 5154 95845 5182
rect 95845 5154 95873 5182
rect 95873 5154 95875 5182
rect 95843 5152 95875 5154
rect 133822 5182 133854 5184
rect 133822 5154 133824 5182
rect 133824 5154 133852 5182
rect 133852 5154 133854 5182
rect 133822 5152 133854 5154
rect 133862 5182 133894 5184
rect 133862 5154 133864 5182
rect 133864 5154 133892 5182
rect 133892 5154 133894 5182
rect 133862 5152 133894 5154
rect 133902 5182 133934 5184
rect 133902 5154 133904 5182
rect 133904 5154 133932 5182
rect 133932 5154 133934 5182
rect 133902 5152 133934 5154
rect 133942 5182 133974 5184
rect 133942 5154 133944 5182
rect 133944 5154 133972 5182
rect 133972 5154 133974 5182
rect 133942 5152 133974 5154
rect 38575 4910 38607 4912
rect 38575 4882 38577 4910
rect 38577 4882 38605 4910
rect 38605 4882 38607 4910
rect 38575 4880 38607 4882
rect 38615 4910 38647 4912
rect 38615 4882 38617 4910
rect 38617 4882 38645 4910
rect 38645 4882 38647 4910
rect 38615 4880 38647 4882
rect 38655 4910 38687 4912
rect 38655 4882 38657 4910
rect 38657 4882 38685 4910
rect 38685 4882 38687 4910
rect 38655 4880 38687 4882
rect 38695 4910 38727 4912
rect 38695 4882 38697 4910
rect 38697 4882 38725 4910
rect 38725 4882 38727 4910
rect 38695 4880 38727 4882
rect 76674 4910 76706 4912
rect 76674 4882 76676 4910
rect 76676 4882 76704 4910
rect 76704 4882 76706 4910
rect 76674 4880 76706 4882
rect 76714 4910 76746 4912
rect 76714 4882 76716 4910
rect 76716 4882 76744 4910
rect 76744 4882 76746 4910
rect 76714 4880 76746 4882
rect 76754 4910 76786 4912
rect 76754 4882 76756 4910
rect 76756 4882 76784 4910
rect 76784 4882 76786 4910
rect 76754 4880 76786 4882
rect 76794 4910 76826 4912
rect 76794 4882 76796 4910
rect 76796 4882 76824 4910
rect 76824 4882 76826 4910
rect 76794 4880 76826 4882
rect 114773 4910 114805 4912
rect 114773 4882 114775 4910
rect 114775 4882 114803 4910
rect 114803 4882 114805 4910
rect 114773 4880 114805 4882
rect 114813 4910 114845 4912
rect 114813 4882 114815 4910
rect 114815 4882 114843 4910
rect 114843 4882 114845 4910
rect 114813 4880 114845 4882
rect 114853 4910 114885 4912
rect 114853 4882 114855 4910
rect 114855 4882 114883 4910
rect 114883 4882 114885 4910
rect 114853 4880 114885 4882
rect 114893 4910 114925 4912
rect 114893 4882 114895 4910
rect 114895 4882 114923 4910
rect 114923 4882 114925 4910
rect 114893 4880 114925 4882
rect 19525 4638 19557 4640
rect 19525 4610 19527 4638
rect 19527 4610 19555 4638
rect 19555 4610 19557 4638
rect 19525 4608 19557 4610
rect 19565 4638 19597 4640
rect 19565 4610 19567 4638
rect 19567 4610 19595 4638
rect 19595 4610 19597 4638
rect 19565 4608 19597 4610
rect 19605 4638 19637 4640
rect 19605 4610 19607 4638
rect 19607 4610 19635 4638
rect 19635 4610 19637 4638
rect 19605 4608 19637 4610
rect 19645 4638 19677 4640
rect 19645 4610 19647 4638
rect 19647 4610 19675 4638
rect 19675 4610 19677 4638
rect 19645 4608 19677 4610
rect 57624 4638 57656 4640
rect 57624 4610 57626 4638
rect 57626 4610 57654 4638
rect 57654 4610 57656 4638
rect 57624 4608 57656 4610
rect 57664 4638 57696 4640
rect 57664 4610 57666 4638
rect 57666 4610 57694 4638
rect 57694 4610 57696 4638
rect 57664 4608 57696 4610
rect 57704 4638 57736 4640
rect 57704 4610 57706 4638
rect 57706 4610 57734 4638
rect 57734 4610 57736 4638
rect 57704 4608 57736 4610
rect 57744 4638 57776 4640
rect 57744 4610 57746 4638
rect 57746 4610 57774 4638
rect 57774 4610 57776 4638
rect 57744 4608 57776 4610
rect 95723 4638 95755 4640
rect 95723 4610 95725 4638
rect 95725 4610 95753 4638
rect 95753 4610 95755 4638
rect 95723 4608 95755 4610
rect 95763 4638 95795 4640
rect 95763 4610 95765 4638
rect 95765 4610 95793 4638
rect 95793 4610 95795 4638
rect 95763 4608 95795 4610
rect 95803 4638 95835 4640
rect 95803 4610 95805 4638
rect 95805 4610 95833 4638
rect 95833 4610 95835 4638
rect 95803 4608 95835 4610
rect 95843 4638 95875 4640
rect 95843 4610 95845 4638
rect 95845 4610 95873 4638
rect 95873 4610 95875 4638
rect 95843 4608 95875 4610
rect 133822 4638 133854 4640
rect 133822 4610 133824 4638
rect 133824 4610 133852 4638
rect 133852 4610 133854 4638
rect 133822 4608 133854 4610
rect 133862 4638 133894 4640
rect 133862 4610 133864 4638
rect 133864 4610 133892 4638
rect 133892 4610 133894 4638
rect 133862 4608 133894 4610
rect 133902 4638 133934 4640
rect 133902 4610 133904 4638
rect 133904 4610 133932 4638
rect 133932 4610 133934 4638
rect 133902 4608 133934 4610
rect 133942 4638 133974 4640
rect 133942 4610 133944 4638
rect 133944 4610 133972 4638
rect 133972 4610 133974 4638
rect 133942 4608 133974 4610
rect 38575 4366 38607 4368
rect 38575 4338 38577 4366
rect 38577 4338 38605 4366
rect 38605 4338 38607 4366
rect 38575 4336 38607 4338
rect 38615 4366 38647 4368
rect 38615 4338 38617 4366
rect 38617 4338 38645 4366
rect 38645 4338 38647 4366
rect 38615 4336 38647 4338
rect 38655 4366 38687 4368
rect 38655 4338 38657 4366
rect 38657 4338 38685 4366
rect 38685 4338 38687 4366
rect 38655 4336 38687 4338
rect 38695 4366 38727 4368
rect 38695 4338 38697 4366
rect 38697 4338 38725 4366
rect 38725 4338 38727 4366
rect 38695 4336 38727 4338
rect 76674 4366 76706 4368
rect 76674 4338 76676 4366
rect 76676 4338 76704 4366
rect 76704 4338 76706 4366
rect 76674 4336 76706 4338
rect 76714 4366 76746 4368
rect 76714 4338 76716 4366
rect 76716 4338 76744 4366
rect 76744 4338 76746 4366
rect 76714 4336 76746 4338
rect 76754 4366 76786 4368
rect 76754 4338 76756 4366
rect 76756 4338 76784 4366
rect 76784 4338 76786 4366
rect 76754 4336 76786 4338
rect 76794 4366 76826 4368
rect 76794 4338 76796 4366
rect 76796 4338 76824 4366
rect 76824 4338 76826 4366
rect 76794 4336 76826 4338
rect 114773 4366 114805 4368
rect 114773 4338 114775 4366
rect 114775 4338 114803 4366
rect 114803 4338 114805 4366
rect 114773 4336 114805 4338
rect 114813 4366 114845 4368
rect 114813 4338 114815 4366
rect 114815 4338 114843 4366
rect 114843 4338 114845 4366
rect 114813 4336 114845 4338
rect 114853 4366 114885 4368
rect 114853 4338 114855 4366
rect 114855 4338 114883 4366
rect 114883 4338 114885 4366
rect 114853 4336 114885 4338
rect 114893 4366 114925 4368
rect 114893 4338 114895 4366
rect 114895 4338 114923 4366
rect 114923 4338 114925 4366
rect 114893 4336 114925 4338
rect 19525 4094 19557 4096
rect 19525 4066 19527 4094
rect 19527 4066 19555 4094
rect 19555 4066 19557 4094
rect 19525 4064 19557 4066
rect 19565 4094 19597 4096
rect 19565 4066 19567 4094
rect 19567 4066 19595 4094
rect 19595 4066 19597 4094
rect 19565 4064 19597 4066
rect 19605 4094 19637 4096
rect 19605 4066 19607 4094
rect 19607 4066 19635 4094
rect 19635 4066 19637 4094
rect 19605 4064 19637 4066
rect 19645 4094 19677 4096
rect 19645 4066 19647 4094
rect 19647 4066 19675 4094
rect 19675 4066 19677 4094
rect 19645 4064 19677 4066
rect 57624 4094 57656 4096
rect 57624 4066 57626 4094
rect 57626 4066 57654 4094
rect 57654 4066 57656 4094
rect 57624 4064 57656 4066
rect 57664 4094 57696 4096
rect 57664 4066 57666 4094
rect 57666 4066 57694 4094
rect 57694 4066 57696 4094
rect 57664 4064 57696 4066
rect 57704 4094 57736 4096
rect 57704 4066 57706 4094
rect 57706 4066 57734 4094
rect 57734 4066 57736 4094
rect 57704 4064 57736 4066
rect 57744 4094 57776 4096
rect 57744 4066 57746 4094
rect 57746 4066 57774 4094
rect 57774 4066 57776 4094
rect 57744 4064 57776 4066
rect 95723 4094 95755 4096
rect 95723 4066 95725 4094
rect 95725 4066 95753 4094
rect 95753 4066 95755 4094
rect 95723 4064 95755 4066
rect 95763 4094 95795 4096
rect 95763 4066 95765 4094
rect 95765 4066 95793 4094
rect 95793 4066 95795 4094
rect 95763 4064 95795 4066
rect 95803 4094 95835 4096
rect 95803 4066 95805 4094
rect 95805 4066 95833 4094
rect 95833 4066 95835 4094
rect 95803 4064 95835 4066
rect 95843 4094 95875 4096
rect 95843 4066 95845 4094
rect 95845 4066 95873 4094
rect 95873 4066 95875 4094
rect 95843 4064 95875 4066
rect 133822 4094 133854 4096
rect 133822 4066 133824 4094
rect 133824 4066 133852 4094
rect 133852 4066 133854 4094
rect 133822 4064 133854 4066
rect 133862 4094 133894 4096
rect 133862 4066 133864 4094
rect 133864 4066 133892 4094
rect 133892 4066 133894 4094
rect 133862 4064 133894 4066
rect 133902 4094 133934 4096
rect 133902 4066 133904 4094
rect 133904 4066 133932 4094
rect 133932 4066 133934 4094
rect 133902 4064 133934 4066
rect 133942 4094 133974 4096
rect 133942 4066 133944 4094
rect 133944 4066 133972 4094
rect 133972 4066 133974 4094
rect 133942 4064 133974 4066
rect 38575 3822 38607 3824
rect 38575 3794 38577 3822
rect 38577 3794 38605 3822
rect 38605 3794 38607 3822
rect 38575 3792 38607 3794
rect 38615 3822 38647 3824
rect 38615 3794 38617 3822
rect 38617 3794 38645 3822
rect 38645 3794 38647 3822
rect 38615 3792 38647 3794
rect 38655 3822 38687 3824
rect 38655 3794 38657 3822
rect 38657 3794 38685 3822
rect 38685 3794 38687 3822
rect 38655 3792 38687 3794
rect 38695 3822 38727 3824
rect 38695 3794 38697 3822
rect 38697 3794 38725 3822
rect 38725 3794 38727 3822
rect 38695 3792 38727 3794
rect 76674 3822 76706 3824
rect 76674 3794 76676 3822
rect 76676 3794 76704 3822
rect 76704 3794 76706 3822
rect 76674 3792 76706 3794
rect 76714 3822 76746 3824
rect 76714 3794 76716 3822
rect 76716 3794 76744 3822
rect 76744 3794 76746 3822
rect 76714 3792 76746 3794
rect 76754 3822 76786 3824
rect 76754 3794 76756 3822
rect 76756 3794 76784 3822
rect 76784 3794 76786 3822
rect 76754 3792 76786 3794
rect 76794 3822 76826 3824
rect 76794 3794 76796 3822
rect 76796 3794 76824 3822
rect 76824 3794 76826 3822
rect 76794 3792 76826 3794
rect 114773 3822 114805 3824
rect 114773 3794 114775 3822
rect 114775 3794 114803 3822
rect 114803 3794 114805 3822
rect 114773 3792 114805 3794
rect 114813 3822 114845 3824
rect 114813 3794 114815 3822
rect 114815 3794 114843 3822
rect 114843 3794 114845 3822
rect 114813 3792 114845 3794
rect 114853 3822 114885 3824
rect 114853 3794 114855 3822
rect 114855 3794 114883 3822
rect 114883 3794 114885 3822
rect 114853 3792 114885 3794
rect 114893 3822 114925 3824
rect 114893 3794 114895 3822
rect 114895 3794 114923 3822
rect 114923 3794 114925 3822
rect 114893 3792 114925 3794
rect 19525 3550 19557 3552
rect 19525 3522 19527 3550
rect 19527 3522 19555 3550
rect 19555 3522 19557 3550
rect 19525 3520 19557 3522
rect 19565 3550 19597 3552
rect 19565 3522 19567 3550
rect 19567 3522 19595 3550
rect 19595 3522 19597 3550
rect 19565 3520 19597 3522
rect 19605 3550 19637 3552
rect 19605 3522 19607 3550
rect 19607 3522 19635 3550
rect 19635 3522 19637 3550
rect 19605 3520 19637 3522
rect 19645 3550 19677 3552
rect 19645 3522 19647 3550
rect 19647 3522 19675 3550
rect 19675 3522 19677 3550
rect 19645 3520 19677 3522
rect 57624 3550 57656 3552
rect 57624 3522 57626 3550
rect 57626 3522 57654 3550
rect 57654 3522 57656 3550
rect 57624 3520 57656 3522
rect 57664 3550 57696 3552
rect 57664 3522 57666 3550
rect 57666 3522 57694 3550
rect 57694 3522 57696 3550
rect 57664 3520 57696 3522
rect 57704 3550 57736 3552
rect 57704 3522 57706 3550
rect 57706 3522 57734 3550
rect 57734 3522 57736 3550
rect 57704 3520 57736 3522
rect 57744 3550 57776 3552
rect 57744 3522 57746 3550
rect 57746 3522 57774 3550
rect 57774 3522 57776 3550
rect 57744 3520 57776 3522
rect 95723 3550 95755 3552
rect 95723 3522 95725 3550
rect 95725 3522 95753 3550
rect 95753 3522 95755 3550
rect 95723 3520 95755 3522
rect 95763 3550 95795 3552
rect 95763 3522 95765 3550
rect 95765 3522 95793 3550
rect 95793 3522 95795 3550
rect 95763 3520 95795 3522
rect 95803 3550 95835 3552
rect 95803 3522 95805 3550
rect 95805 3522 95833 3550
rect 95833 3522 95835 3550
rect 95803 3520 95835 3522
rect 95843 3550 95875 3552
rect 95843 3522 95845 3550
rect 95845 3522 95873 3550
rect 95873 3522 95875 3550
rect 95843 3520 95875 3522
rect 133822 3550 133854 3552
rect 133822 3522 133824 3550
rect 133824 3522 133852 3550
rect 133852 3522 133854 3550
rect 133822 3520 133854 3522
rect 133862 3550 133894 3552
rect 133862 3522 133864 3550
rect 133864 3522 133892 3550
rect 133892 3522 133894 3550
rect 133862 3520 133894 3522
rect 133902 3550 133934 3552
rect 133902 3522 133904 3550
rect 133904 3522 133932 3550
rect 133932 3522 133934 3550
rect 133902 3520 133934 3522
rect 133942 3550 133974 3552
rect 133942 3522 133944 3550
rect 133944 3522 133972 3550
rect 133972 3522 133974 3550
rect 133942 3520 133974 3522
rect 38575 3278 38607 3280
rect 38575 3250 38577 3278
rect 38577 3250 38605 3278
rect 38605 3250 38607 3278
rect 38575 3248 38607 3250
rect 38615 3278 38647 3280
rect 38615 3250 38617 3278
rect 38617 3250 38645 3278
rect 38645 3250 38647 3278
rect 38615 3248 38647 3250
rect 38655 3278 38687 3280
rect 38655 3250 38657 3278
rect 38657 3250 38685 3278
rect 38685 3250 38687 3278
rect 38655 3248 38687 3250
rect 38695 3278 38727 3280
rect 38695 3250 38697 3278
rect 38697 3250 38725 3278
rect 38725 3250 38727 3278
rect 38695 3248 38727 3250
rect 76674 3278 76706 3280
rect 76674 3250 76676 3278
rect 76676 3250 76704 3278
rect 76704 3250 76706 3278
rect 76674 3248 76706 3250
rect 76714 3278 76746 3280
rect 76714 3250 76716 3278
rect 76716 3250 76744 3278
rect 76744 3250 76746 3278
rect 76714 3248 76746 3250
rect 76754 3278 76786 3280
rect 76754 3250 76756 3278
rect 76756 3250 76784 3278
rect 76784 3250 76786 3278
rect 76754 3248 76786 3250
rect 76794 3278 76826 3280
rect 76794 3250 76796 3278
rect 76796 3250 76824 3278
rect 76824 3250 76826 3278
rect 76794 3248 76826 3250
rect 114773 3278 114805 3280
rect 114773 3250 114775 3278
rect 114775 3250 114803 3278
rect 114803 3250 114805 3278
rect 114773 3248 114805 3250
rect 114813 3278 114845 3280
rect 114813 3250 114815 3278
rect 114815 3250 114843 3278
rect 114843 3250 114845 3278
rect 114813 3248 114845 3250
rect 114853 3278 114885 3280
rect 114853 3250 114855 3278
rect 114855 3250 114883 3278
rect 114883 3250 114885 3278
rect 114853 3248 114885 3250
rect 114893 3278 114925 3280
rect 114893 3250 114895 3278
rect 114895 3250 114923 3278
rect 114923 3250 114925 3278
rect 114893 3248 114925 3250
rect 19525 3006 19557 3008
rect 19525 2978 19527 3006
rect 19527 2978 19555 3006
rect 19555 2978 19557 3006
rect 19525 2976 19557 2978
rect 19565 3006 19597 3008
rect 19565 2978 19567 3006
rect 19567 2978 19595 3006
rect 19595 2978 19597 3006
rect 19565 2976 19597 2978
rect 19605 3006 19637 3008
rect 19605 2978 19607 3006
rect 19607 2978 19635 3006
rect 19635 2978 19637 3006
rect 19605 2976 19637 2978
rect 19645 3006 19677 3008
rect 19645 2978 19647 3006
rect 19647 2978 19675 3006
rect 19675 2978 19677 3006
rect 19645 2976 19677 2978
rect 57624 3006 57656 3008
rect 57624 2978 57626 3006
rect 57626 2978 57654 3006
rect 57654 2978 57656 3006
rect 57624 2976 57656 2978
rect 57664 3006 57696 3008
rect 57664 2978 57666 3006
rect 57666 2978 57694 3006
rect 57694 2978 57696 3006
rect 57664 2976 57696 2978
rect 57704 3006 57736 3008
rect 57704 2978 57706 3006
rect 57706 2978 57734 3006
rect 57734 2978 57736 3006
rect 57704 2976 57736 2978
rect 57744 3006 57776 3008
rect 57744 2978 57746 3006
rect 57746 2978 57774 3006
rect 57774 2978 57776 3006
rect 57744 2976 57776 2978
rect 95723 3006 95755 3008
rect 95723 2978 95725 3006
rect 95725 2978 95753 3006
rect 95753 2978 95755 3006
rect 95723 2976 95755 2978
rect 95763 3006 95795 3008
rect 95763 2978 95765 3006
rect 95765 2978 95793 3006
rect 95793 2978 95795 3006
rect 95763 2976 95795 2978
rect 95803 3006 95835 3008
rect 95803 2978 95805 3006
rect 95805 2978 95833 3006
rect 95833 2978 95835 3006
rect 95803 2976 95835 2978
rect 95843 3006 95875 3008
rect 95843 2978 95845 3006
rect 95845 2978 95873 3006
rect 95873 2978 95875 3006
rect 95843 2976 95875 2978
rect 133822 3006 133854 3008
rect 133822 2978 133824 3006
rect 133824 2978 133852 3006
rect 133852 2978 133854 3006
rect 133822 2976 133854 2978
rect 133862 3006 133894 3008
rect 133862 2978 133864 3006
rect 133864 2978 133892 3006
rect 133892 2978 133894 3006
rect 133862 2976 133894 2978
rect 133902 3006 133934 3008
rect 133902 2978 133904 3006
rect 133904 2978 133932 3006
rect 133932 2978 133934 3006
rect 133902 2976 133934 2978
rect 133942 3006 133974 3008
rect 133942 2978 133944 3006
rect 133944 2978 133972 3006
rect 133972 2978 133974 3006
rect 133942 2976 133974 2978
rect 38575 2734 38607 2736
rect 38575 2706 38577 2734
rect 38577 2706 38605 2734
rect 38605 2706 38607 2734
rect 38575 2704 38607 2706
rect 38615 2734 38647 2736
rect 38615 2706 38617 2734
rect 38617 2706 38645 2734
rect 38645 2706 38647 2734
rect 38615 2704 38647 2706
rect 38655 2734 38687 2736
rect 38655 2706 38657 2734
rect 38657 2706 38685 2734
rect 38685 2706 38687 2734
rect 38655 2704 38687 2706
rect 38695 2734 38727 2736
rect 38695 2706 38697 2734
rect 38697 2706 38725 2734
rect 38725 2706 38727 2734
rect 38695 2704 38727 2706
rect 76674 2734 76706 2736
rect 76674 2706 76676 2734
rect 76676 2706 76704 2734
rect 76704 2706 76706 2734
rect 76674 2704 76706 2706
rect 76714 2734 76746 2736
rect 76714 2706 76716 2734
rect 76716 2706 76744 2734
rect 76744 2706 76746 2734
rect 76714 2704 76746 2706
rect 76754 2734 76786 2736
rect 76754 2706 76756 2734
rect 76756 2706 76784 2734
rect 76784 2706 76786 2734
rect 76754 2704 76786 2706
rect 76794 2734 76826 2736
rect 76794 2706 76796 2734
rect 76796 2706 76824 2734
rect 76824 2706 76826 2734
rect 76794 2704 76826 2706
rect 114773 2734 114805 2736
rect 114773 2706 114775 2734
rect 114775 2706 114803 2734
rect 114803 2706 114805 2734
rect 114773 2704 114805 2706
rect 114813 2734 114845 2736
rect 114813 2706 114815 2734
rect 114815 2706 114843 2734
rect 114843 2706 114845 2734
rect 114813 2704 114845 2706
rect 114853 2734 114885 2736
rect 114853 2706 114855 2734
rect 114855 2706 114883 2734
rect 114883 2706 114885 2734
rect 114853 2704 114885 2706
rect 114893 2734 114925 2736
rect 114893 2706 114895 2734
rect 114895 2706 114923 2734
rect 114923 2706 114925 2734
rect 114893 2704 114925 2706
rect 19525 2462 19557 2464
rect 19525 2434 19527 2462
rect 19527 2434 19555 2462
rect 19555 2434 19557 2462
rect 19525 2432 19557 2434
rect 19565 2462 19597 2464
rect 19565 2434 19567 2462
rect 19567 2434 19595 2462
rect 19595 2434 19597 2462
rect 19565 2432 19597 2434
rect 19605 2462 19637 2464
rect 19605 2434 19607 2462
rect 19607 2434 19635 2462
rect 19635 2434 19637 2462
rect 19605 2432 19637 2434
rect 19645 2462 19677 2464
rect 19645 2434 19647 2462
rect 19647 2434 19675 2462
rect 19675 2434 19677 2462
rect 19645 2432 19677 2434
rect 57624 2462 57656 2464
rect 57624 2434 57626 2462
rect 57626 2434 57654 2462
rect 57654 2434 57656 2462
rect 57624 2432 57656 2434
rect 57664 2462 57696 2464
rect 57664 2434 57666 2462
rect 57666 2434 57694 2462
rect 57694 2434 57696 2462
rect 57664 2432 57696 2434
rect 57704 2462 57736 2464
rect 57704 2434 57706 2462
rect 57706 2434 57734 2462
rect 57734 2434 57736 2462
rect 57704 2432 57736 2434
rect 57744 2462 57776 2464
rect 57744 2434 57746 2462
rect 57746 2434 57774 2462
rect 57774 2434 57776 2462
rect 57744 2432 57776 2434
rect 95723 2462 95755 2464
rect 95723 2434 95725 2462
rect 95725 2434 95753 2462
rect 95753 2434 95755 2462
rect 95723 2432 95755 2434
rect 95763 2462 95795 2464
rect 95763 2434 95765 2462
rect 95765 2434 95793 2462
rect 95793 2434 95795 2462
rect 95763 2432 95795 2434
rect 95803 2462 95835 2464
rect 95803 2434 95805 2462
rect 95805 2434 95833 2462
rect 95833 2434 95835 2462
rect 95803 2432 95835 2434
rect 95843 2462 95875 2464
rect 95843 2434 95845 2462
rect 95845 2434 95873 2462
rect 95873 2434 95875 2462
rect 95843 2432 95875 2434
rect 133822 2462 133854 2464
rect 133822 2434 133824 2462
rect 133824 2434 133852 2462
rect 133852 2434 133854 2462
rect 133822 2432 133854 2434
rect 133862 2462 133894 2464
rect 133862 2434 133864 2462
rect 133864 2434 133892 2462
rect 133892 2434 133894 2462
rect 133862 2432 133894 2434
rect 133902 2462 133934 2464
rect 133902 2434 133904 2462
rect 133904 2434 133932 2462
rect 133932 2434 133934 2462
rect 133902 2432 133934 2434
rect 133942 2462 133974 2464
rect 133942 2434 133944 2462
rect 133944 2434 133972 2462
rect 133972 2434 133974 2462
rect 133942 2432 133974 2434
rect 38575 2190 38607 2192
rect 38575 2162 38577 2190
rect 38577 2162 38605 2190
rect 38605 2162 38607 2190
rect 38575 2160 38607 2162
rect 38615 2190 38647 2192
rect 38615 2162 38617 2190
rect 38617 2162 38645 2190
rect 38645 2162 38647 2190
rect 38615 2160 38647 2162
rect 38655 2190 38687 2192
rect 38655 2162 38657 2190
rect 38657 2162 38685 2190
rect 38685 2162 38687 2190
rect 38655 2160 38687 2162
rect 38695 2190 38727 2192
rect 38695 2162 38697 2190
rect 38697 2162 38725 2190
rect 38725 2162 38727 2190
rect 38695 2160 38727 2162
rect 76674 2190 76706 2192
rect 76674 2162 76676 2190
rect 76676 2162 76704 2190
rect 76704 2162 76706 2190
rect 76674 2160 76706 2162
rect 76714 2190 76746 2192
rect 76714 2162 76716 2190
rect 76716 2162 76744 2190
rect 76744 2162 76746 2190
rect 76714 2160 76746 2162
rect 76754 2190 76786 2192
rect 76754 2162 76756 2190
rect 76756 2162 76784 2190
rect 76784 2162 76786 2190
rect 76754 2160 76786 2162
rect 76794 2190 76826 2192
rect 76794 2162 76796 2190
rect 76796 2162 76824 2190
rect 76824 2162 76826 2190
rect 76794 2160 76826 2162
rect 114773 2190 114805 2192
rect 114773 2162 114775 2190
rect 114775 2162 114803 2190
rect 114803 2162 114805 2190
rect 114773 2160 114805 2162
rect 114813 2190 114845 2192
rect 114813 2162 114815 2190
rect 114815 2162 114843 2190
rect 114843 2162 114845 2190
rect 114813 2160 114845 2162
rect 114853 2190 114885 2192
rect 114853 2162 114855 2190
rect 114855 2162 114883 2190
rect 114883 2162 114885 2190
rect 114853 2160 114885 2162
rect 114893 2190 114925 2192
rect 114893 2162 114895 2190
rect 114895 2162 114923 2190
rect 114923 2162 114925 2190
rect 114893 2160 114925 2162
rect 19525 1918 19557 1920
rect 19525 1890 19527 1918
rect 19527 1890 19555 1918
rect 19555 1890 19557 1918
rect 19525 1888 19557 1890
rect 19565 1918 19597 1920
rect 19565 1890 19567 1918
rect 19567 1890 19595 1918
rect 19595 1890 19597 1918
rect 19565 1888 19597 1890
rect 19605 1918 19637 1920
rect 19605 1890 19607 1918
rect 19607 1890 19635 1918
rect 19635 1890 19637 1918
rect 19605 1888 19637 1890
rect 19645 1918 19677 1920
rect 19645 1890 19647 1918
rect 19647 1890 19675 1918
rect 19675 1890 19677 1918
rect 19645 1888 19677 1890
rect 57624 1918 57656 1920
rect 57624 1890 57626 1918
rect 57626 1890 57654 1918
rect 57654 1890 57656 1918
rect 57624 1888 57656 1890
rect 57664 1918 57696 1920
rect 57664 1890 57666 1918
rect 57666 1890 57694 1918
rect 57694 1890 57696 1918
rect 57664 1888 57696 1890
rect 57704 1918 57736 1920
rect 57704 1890 57706 1918
rect 57706 1890 57734 1918
rect 57734 1890 57736 1918
rect 57704 1888 57736 1890
rect 57744 1918 57776 1920
rect 57744 1890 57746 1918
rect 57746 1890 57774 1918
rect 57774 1890 57776 1918
rect 57744 1888 57776 1890
rect 95723 1918 95755 1920
rect 95723 1890 95725 1918
rect 95725 1890 95753 1918
rect 95753 1890 95755 1918
rect 95723 1888 95755 1890
rect 95763 1918 95795 1920
rect 95763 1890 95765 1918
rect 95765 1890 95793 1918
rect 95793 1890 95795 1918
rect 95763 1888 95795 1890
rect 95803 1918 95835 1920
rect 95803 1890 95805 1918
rect 95805 1890 95833 1918
rect 95833 1890 95835 1918
rect 95803 1888 95835 1890
rect 95843 1918 95875 1920
rect 95843 1890 95845 1918
rect 95845 1890 95873 1918
rect 95873 1890 95875 1918
rect 95843 1888 95875 1890
rect 133822 1918 133854 1920
rect 133822 1890 133824 1918
rect 133824 1890 133852 1918
rect 133852 1890 133854 1918
rect 133822 1888 133854 1890
rect 133862 1918 133894 1920
rect 133862 1890 133864 1918
rect 133864 1890 133892 1918
rect 133892 1890 133894 1918
rect 133862 1888 133894 1890
rect 133902 1918 133934 1920
rect 133902 1890 133904 1918
rect 133904 1890 133932 1918
rect 133932 1890 133934 1918
rect 133902 1888 133934 1890
rect 133942 1918 133974 1920
rect 133942 1890 133944 1918
rect 133944 1890 133972 1918
rect 133972 1890 133974 1918
rect 133942 1888 133974 1890
rect 38575 1646 38607 1648
rect 38575 1618 38577 1646
rect 38577 1618 38605 1646
rect 38605 1618 38607 1646
rect 38575 1616 38607 1618
rect 38615 1646 38647 1648
rect 38615 1618 38617 1646
rect 38617 1618 38645 1646
rect 38645 1618 38647 1646
rect 38615 1616 38647 1618
rect 38655 1646 38687 1648
rect 38655 1618 38657 1646
rect 38657 1618 38685 1646
rect 38685 1618 38687 1646
rect 38655 1616 38687 1618
rect 38695 1646 38727 1648
rect 38695 1618 38697 1646
rect 38697 1618 38725 1646
rect 38725 1618 38727 1646
rect 38695 1616 38727 1618
rect 76674 1646 76706 1648
rect 76674 1618 76676 1646
rect 76676 1618 76704 1646
rect 76704 1618 76706 1646
rect 76674 1616 76706 1618
rect 76714 1646 76746 1648
rect 76714 1618 76716 1646
rect 76716 1618 76744 1646
rect 76744 1618 76746 1646
rect 76714 1616 76746 1618
rect 76754 1646 76786 1648
rect 76754 1618 76756 1646
rect 76756 1618 76784 1646
rect 76784 1618 76786 1646
rect 76754 1616 76786 1618
rect 76794 1646 76826 1648
rect 76794 1618 76796 1646
rect 76796 1618 76824 1646
rect 76824 1618 76826 1646
rect 76794 1616 76826 1618
rect 114773 1646 114805 1648
rect 114773 1618 114775 1646
rect 114775 1618 114803 1646
rect 114803 1618 114805 1646
rect 114773 1616 114805 1618
rect 114813 1646 114845 1648
rect 114813 1618 114815 1646
rect 114815 1618 114843 1646
rect 114843 1618 114845 1646
rect 114813 1616 114845 1618
rect 114853 1646 114885 1648
rect 114853 1618 114855 1646
rect 114855 1618 114883 1646
rect 114883 1618 114885 1646
rect 114853 1616 114885 1618
rect 114893 1646 114925 1648
rect 114893 1618 114895 1646
rect 114895 1618 114923 1646
rect 114923 1618 114925 1646
rect 114893 1616 114925 1618
rect 19525 1374 19557 1376
rect 19525 1346 19527 1374
rect 19527 1346 19555 1374
rect 19555 1346 19557 1374
rect 19525 1344 19557 1346
rect 19565 1374 19597 1376
rect 19565 1346 19567 1374
rect 19567 1346 19595 1374
rect 19595 1346 19597 1374
rect 19565 1344 19597 1346
rect 19605 1374 19637 1376
rect 19605 1346 19607 1374
rect 19607 1346 19635 1374
rect 19635 1346 19637 1374
rect 19605 1344 19637 1346
rect 19645 1374 19677 1376
rect 19645 1346 19647 1374
rect 19647 1346 19675 1374
rect 19675 1346 19677 1374
rect 19645 1344 19677 1346
rect 57624 1374 57656 1376
rect 57624 1346 57626 1374
rect 57626 1346 57654 1374
rect 57654 1346 57656 1374
rect 57624 1344 57656 1346
rect 57664 1374 57696 1376
rect 57664 1346 57666 1374
rect 57666 1346 57694 1374
rect 57694 1346 57696 1374
rect 57664 1344 57696 1346
rect 57704 1374 57736 1376
rect 57704 1346 57706 1374
rect 57706 1346 57734 1374
rect 57734 1346 57736 1374
rect 57704 1344 57736 1346
rect 57744 1374 57776 1376
rect 57744 1346 57746 1374
rect 57746 1346 57774 1374
rect 57774 1346 57776 1374
rect 57744 1344 57776 1346
rect 95723 1374 95755 1376
rect 95723 1346 95725 1374
rect 95725 1346 95753 1374
rect 95753 1346 95755 1374
rect 95723 1344 95755 1346
rect 95763 1374 95795 1376
rect 95763 1346 95765 1374
rect 95765 1346 95793 1374
rect 95793 1346 95795 1374
rect 95763 1344 95795 1346
rect 95803 1374 95835 1376
rect 95803 1346 95805 1374
rect 95805 1346 95833 1374
rect 95833 1346 95835 1374
rect 95803 1344 95835 1346
rect 95843 1374 95875 1376
rect 95843 1346 95845 1374
rect 95845 1346 95873 1374
rect 95873 1346 95875 1374
rect 95843 1344 95875 1346
rect 133822 1374 133854 1376
rect 133822 1346 133824 1374
rect 133824 1346 133852 1374
rect 133852 1346 133854 1374
rect 133822 1344 133854 1346
rect 133862 1374 133894 1376
rect 133862 1346 133864 1374
rect 133864 1346 133892 1374
rect 133892 1346 133894 1374
rect 133862 1344 133894 1346
rect 133902 1374 133934 1376
rect 133902 1346 133904 1374
rect 133904 1346 133932 1374
rect 133932 1346 133934 1374
rect 133902 1344 133934 1346
rect 133942 1374 133974 1376
rect 133942 1346 133944 1374
rect 133944 1346 133972 1374
rect 133972 1346 133974 1374
rect 133942 1344 133974 1346
rect 38575 1102 38607 1104
rect 38575 1074 38577 1102
rect 38577 1074 38605 1102
rect 38605 1074 38607 1102
rect 38575 1072 38607 1074
rect 38615 1102 38647 1104
rect 38615 1074 38617 1102
rect 38617 1074 38645 1102
rect 38645 1074 38647 1102
rect 38615 1072 38647 1074
rect 38655 1102 38687 1104
rect 38655 1074 38657 1102
rect 38657 1074 38685 1102
rect 38685 1074 38687 1102
rect 38655 1072 38687 1074
rect 38695 1102 38727 1104
rect 38695 1074 38697 1102
rect 38697 1074 38725 1102
rect 38725 1074 38727 1102
rect 38695 1072 38727 1074
rect 76674 1102 76706 1104
rect 76674 1074 76676 1102
rect 76676 1074 76704 1102
rect 76704 1074 76706 1102
rect 76674 1072 76706 1074
rect 76714 1102 76746 1104
rect 76714 1074 76716 1102
rect 76716 1074 76744 1102
rect 76744 1074 76746 1102
rect 76714 1072 76746 1074
rect 76754 1102 76786 1104
rect 76754 1074 76756 1102
rect 76756 1074 76784 1102
rect 76784 1074 76786 1102
rect 76754 1072 76786 1074
rect 76794 1102 76826 1104
rect 76794 1074 76796 1102
rect 76796 1074 76824 1102
rect 76824 1074 76826 1102
rect 76794 1072 76826 1074
rect 114773 1102 114805 1104
rect 114773 1074 114775 1102
rect 114775 1074 114803 1102
rect 114803 1074 114805 1102
rect 114773 1072 114805 1074
rect 114813 1102 114845 1104
rect 114813 1074 114815 1102
rect 114815 1074 114843 1102
rect 114843 1074 114845 1102
rect 114813 1072 114845 1074
rect 114853 1102 114885 1104
rect 114853 1074 114855 1102
rect 114855 1074 114883 1102
rect 114883 1074 114885 1102
rect 114853 1072 114885 1074
rect 114893 1102 114925 1104
rect 114893 1074 114895 1102
rect 114895 1074 114923 1102
rect 114923 1074 114925 1102
rect 114893 1072 114925 1074
<< metal4 >>
rect -538 7869 -378 7890
rect -538 7751 -517 7869
rect -399 7751 -378 7869
rect -538 5515 -378 7751
rect -538 5397 -517 5515
rect -399 5397 -378 5515
rect -538 4059 -378 5397
rect -538 3941 -517 4059
rect -399 3941 -378 4059
rect -538 2603 -378 3941
rect -538 2485 -517 2603
rect -399 2485 -378 2603
rect -538 137 -378 2485
rect -208 7539 -48 7560
rect -208 7421 -187 7539
rect -69 7421 -48 7539
rect -208 6243 -48 7421
rect -208 6125 -187 6243
rect -69 6125 -48 6243
rect -208 4787 -48 6125
rect -208 4669 -187 4787
rect -69 4669 -48 4787
rect -208 3331 -48 4669
rect -208 3213 -187 3331
rect -69 3213 -48 3331
rect -208 1875 -48 3213
rect -208 1757 -187 1875
rect -69 1757 -48 1875
rect -208 467 -48 1757
rect -208 349 -187 467
rect -69 349 -48 467
rect -208 328 -48 349
rect 19521 7539 19681 7890
rect 19521 7421 19542 7539
rect 19660 7421 19681 7539
rect 19521 6816 19681 7421
rect 19521 6784 19525 6816
rect 19557 6784 19565 6816
rect 19597 6784 19605 6816
rect 19637 6784 19645 6816
rect 19677 6784 19681 6816
rect 19521 6272 19681 6784
rect 19521 6240 19525 6272
rect 19557 6243 19565 6272
rect 19597 6243 19605 6272
rect 19637 6243 19645 6272
rect 19677 6240 19681 6272
rect 19521 6125 19542 6240
rect 19660 6125 19681 6240
rect 19521 5728 19681 6125
rect 19521 5696 19525 5728
rect 19557 5696 19565 5728
rect 19597 5696 19605 5728
rect 19637 5696 19645 5728
rect 19677 5696 19681 5728
rect 19521 5184 19681 5696
rect 19521 5152 19525 5184
rect 19557 5152 19565 5184
rect 19597 5152 19605 5184
rect 19637 5152 19645 5184
rect 19677 5152 19681 5184
rect 19521 4787 19681 5152
rect 19521 4669 19542 4787
rect 19660 4669 19681 4787
rect 19521 4640 19681 4669
rect 19521 4608 19525 4640
rect 19557 4608 19565 4640
rect 19597 4608 19605 4640
rect 19637 4608 19645 4640
rect 19677 4608 19681 4640
rect 19521 4096 19681 4608
rect 19521 4064 19525 4096
rect 19557 4064 19565 4096
rect 19597 4064 19605 4096
rect 19637 4064 19645 4096
rect 19677 4064 19681 4096
rect 19521 3552 19681 4064
rect 19521 3520 19525 3552
rect 19557 3520 19565 3552
rect 19597 3520 19605 3552
rect 19637 3520 19645 3552
rect 19677 3520 19681 3552
rect 19521 3331 19681 3520
rect 19521 3213 19542 3331
rect 19660 3213 19681 3331
rect 19521 3008 19681 3213
rect 19521 2976 19525 3008
rect 19557 2976 19565 3008
rect 19597 2976 19605 3008
rect 19637 2976 19645 3008
rect 19677 2976 19681 3008
rect 19521 2464 19681 2976
rect 19521 2432 19525 2464
rect 19557 2432 19565 2464
rect 19597 2432 19605 2464
rect 19637 2432 19645 2464
rect 19677 2432 19681 2464
rect 19521 1920 19681 2432
rect 19521 1888 19525 1920
rect 19557 1888 19565 1920
rect 19597 1888 19605 1920
rect 19637 1888 19645 1920
rect 19677 1888 19681 1920
rect 19521 1875 19681 1888
rect 19521 1757 19542 1875
rect 19660 1757 19681 1875
rect 19521 1376 19681 1757
rect 19521 1344 19525 1376
rect 19557 1344 19565 1376
rect 19597 1344 19605 1376
rect 19637 1344 19645 1376
rect 19677 1344 19681 1376
rect 19521 467 19681 1344
rect 19521 349 19542 467
rect 19660 349 19681 467
rect -538 19 -517 137
rect -399 19 -378 137
rect -538 -2 -378 19
rect 19521 -2 19681 349
rect 38571 7869 38731 7890
rect 38571 7751 38592 7869
rect 38710 7751 38731 7869
rect 38571 6544 38731 7751
rect 38571 6512 38575 6544
rect 38607 6512 38615 6544
rect 38647 6512 38655 6544
rect 38687 6512 38695 6544
rect 38727 6512 38731 6544
rect 38571 6000 38731 6512
rect 38571 5968 38575 6000
rect 38607 5968 38615 6000
rect 38647 5968 38655 6000
rect 38687 5968 38695 6000
rect 38727 5968 38731 6000
rect 38571 5515 38731 5968
rect 38571 5456 38592 5515
rect 38710 5456 38731 5515
rect 38571 5424 38575 5456
rect 38727 5424 38731 5456
rect 38571 5397 38592 5424
rect 38710 5397 38731 5424
rect 38571 4912 38731 5397
rect 38571 4880 38575 4912
rect 38607 4880 38615 4912
rect 38647 4880 38655 4912
rect 38687 4880 38695 4912
rect 38727 4880 38731 4912
rect 38571 4368 38731 4880
rect 38571 4336 38575 4368
rect 38607 4336 38615 4368
rect 38647 4336 38655 4368
rect 38687 4336 38695 4368
rect 38727 4336 38731 4368
rect 38571 4059 38731 4336
rect 38571 3941 38592 4059
rect 38710 3941 38731 4059
rect 38571 3824 38731 3941
rect 38571 3792 38575 3824
rect 38607 3792 38615 3824
rect 38647 3792 38655 3824
rect 38687 3792 38695 3824
rect 38727 3792 38731 3824
rect 38571 3280 38731 3792
rect 38571 3248 38575 3280
rect 38607 3248 38615 3280
rect 38647 3248 38655 3280
rect 38687 3248 38695 3280
rect 38727 3248 38731 3280
rect 38571 2736 38731 3248
rect 38571 2704 38575 2736
rect 38607 2704 38615 2736
rect 38647 2704 38655 2736
rect 38687 2704 38695 2736
rect 38727 2704 38731 2736
rect 38571 2603 38731 2704
rect 38571 2485 38592 2603
rect 38710 2485 38731 2603
rect 38571 2192 38731 2485
rect 38571 2160 38575 2192
rect 38607 2160 38615 2192
rect 38647 2160 38655 2192
rect 38687 2160 38695 2192
rect 38727 2160 38731 2192
rect 38571 1648 38731 2160
rect 38571 1616 38575 1648
rect 38607 1616 38615 1648
rect 38647 1616 38655 1648
rect 38687 1616 38695 1648
rect 38727 1616 38731 1648
rect 38571 1104 38731 1616
rect 38571 1072 38575 1104
rect 38607 1072 38615 1104
rect 38647 1072 38655 1104
rect 38687 1072 38695 1104
rect 38727 1072 38731 1104
rect 38571 137 38731 1072
rect 38571 19 38592 137
rect 38710 19 38731 137
rect 38571 -2 38731 19
rect 57620 7539 57780 7890
rect 57620 7421 57641 7539
rect 57759 7421 57780 7539
rect 57620 6816 57780 7421
rect 57620 6784 57624 6816
rect 57656 6784 57664 6816
rect 57696 6784 57704 6816
rect 57736 6784 57744 6816
rect 57776 6784 57780 6816
rect 57620 6272 57780 6784
rect 57620 6240 57624 6272
rect 57656 6243 57664 6272
rect 57696 6243 57704 6272
rect 57736 6243 57744 6272
rect 57776 6240 57780 6272
rect 57620 6125 57641 6240
rect 57759 6125 57780 6240
rect 57620 5728 57780 6125
rect 57620 5696 57624 5728
rect 57656 5696 57664 5728
rect 57696 5696 57704 5728
rect 57736 5696 57744 5728
rect 57776 5696 57780 5728
rect 57620 5184 57780 5696
rect 57620 5152 57624 5184
rect 57656 5152 57664 5184
rect 57696 5152 57704 5184
rect 57736 5152 57744 5184
rect 57776 5152 57780 5184
rect 57620 4787 57780 5152
rect 57620 4669 57641 4787
rect 57759 4669 57780 4787
rect 57620 4640 57780 4669
rect 57620 4608 57624 4640
rect 57656 4608 57664 4640
rect 57696 4608 57704 4640
rect 57736 4608 57744 4640
rect 57776 4608 57780 4640
rect 57620 4096 57780 4608
rect 57620 4064 57624 4096
rect 57656 4064 57664 4096
rect 57696 4064 57704 4096
rect 57736 4064 57744 4096
rect 57776 4064 57780 4096
rect 57620 3552 57780 4064
rect 57620 3520 57624 3552
rect 57656 3520 57664 3552
rect 57696 3520 57704 3552
rect 57736 3520 57744 3552
rect 57776 3520 57780 3552
rect 57620 3331 57780 3520
rect 57620 3213 57641 3331
rect 57759 3213 57780 3331
rect 57620 3008 57780 3213
rect 57620 2976 57624 3008
rect 57656 2976 57664 3008
rect 57696 2976 57704 3008
rect 57736 2976 57744 3008
rect 57776 2976 57780 3008
rect 57620 2464 57780 2976
rect 57620 2432 57624 2464
rect 57656 2432 57664 2464
rect 57696 2432 57704 2464
rect 57736 2432 57744 2464
rect 57776 2432 57780 2464
rect 57620 1920 57780 2432
rect 57620 1888 57624 1920
rect 57656 1888 57664 1920
rect 57696 1888 57704 1920
rect 57736 1888 57744 1920
rect 57776 1888 57780 1920
rect 57620 1875 57780 1888
rect 57620 1757 57641 1875
rect 57759 1757 57780 1875
rect 57620 1376 57780 1757
rect 57620 1344 57624 1376
rect 57656 1344 57664 1376
rect 57696 1344 57704 1376
rect 57736 1344 57744 1376
rect 57776 1344 57780 1376
rect 57620 467 57780 1344
rect 57620 349 57641 467
rect 57759 349 57780 467
rect 57620 -2 57780 349
rect 76670 7869 76830 7890
rect 76670 7751 76691 7869
rect 76809 7751 76830 7869
rect 76670 6544 76830 7751
rect 76670 6512 76674 6544
rect 76706 6512 76714 6544
rect 76746 6512 76754 6544
rect 76786 6512 76794 6544
rect 76826 6512 76830 6544
rect 76670 6000 76830 6512
rect 76670 5968 76674 6000
rect 76706 5968 76714 6000
rect 76746 5968 76754 6000
rect 76786 5968 76794 6000
rect 76826 5968 76830 6000
rect 76670 5515 76830 5968
rect 76670 5456 76691 5515
rect 76809 5456 76830 5515
rect 76670 5424 76674 5456
rect 76826 5424 76830 5456
rect 76670 5397 76691 5424
rect 76809 5397 76830 5424
rect 76670 4912 76830 5397
rect 76670 4880 76674 4912
rect 76706 4880 76714 4912
rect 76746 4880 76754 4912
rect 76786 4880 76794 4912
rect 76826 4880 76830 4912
rect 76670 4368 76830 4880
rect 76670 4336 76674 4368
rect 76706 4336 76714 4368
rect 76746 4336 76754 4368
rect 76786 4336 76794 4368
rect 76826 4336 76830 4368
rect 76670 4059 76830 4336
rect 76670 3941 76691 4059
rect 76809 3941 76830 4059
rect 76670 3824 76830 3941
rect 76670 3792 76674 3824
rect 76706 3792 76714 3824
rect 76746 3792 76754 3824
rect 76786 3792 76794 3824
rect 76826 3792 76830 3824
rect 76670 3280 76830 3792
rect 76670 3248 76674 3280
rect 76706 3248 76714 3280
rect 76746 3248 76754 3280
rect 76786 3248 76794 3280
rect 76826 3248 76830 3280
rect 76670 2736 76830 3248
rect 76670 2704 76674 2736
rect 76706 2704 76714 2736
rect 76746 2704 76754 2736
rect 76786 2704 76794 2736
rect 76826 2704 76830 2736
rect 76670 2603 76830 2704
rect 76670 2485 76691 2603
rect 76809 2485 76830 2603
rect 76670 2192 76830 2485
rect 76670 2160 76674 2192
rect 76706 2160 76714 2192
rect 76746 2160 76754 2192
rect 76786 2160 76794 2192
rect 76826 2160 76830 2192
rect 76670 1648 76830 2160
rect 76670 1616 76674 1648
rect 76706 1616 76714 1648
rect 76746 1616 76754 1648
rect 76786 1616 76794 1648
rect 76826 1616 76830 1648
rect 76670 1104 76830 1616
rect 76670 1072 76674 1104
rect 76706 1072 76714 1104
rect 76746 1072 76754 1104
rect 76786 1072 76794 1104
rect 76826 1072 76830 1104
rect 76670 137 76830 1072
rect 76670 19 76691 137
rect 76809 19 76830 137
rect 76670 -2 76830 19
rect 95719 7539 95879 7890
rect 95719 7421 95740 7539
rect 95858 7421 95879 7539
rect 95719 6816 95879 7421
rect 95719 6784 95723 6816
rect 95755 6784 95763 6816
rect 95795 6784 95803 6816
rect 95835 6784 95843 6816
rect 95875 6784 95879 6816
rect 95719 6272 95879 6784
rect 95719 6240 95723 6272
rect 95755 6243 95763 6272
rect 95795 6243 95803 6272
rect 95835 6243 95843 6272
rect 95875 6240 95879 6272
rect 95719 6125 95740 6240
rect 95858 6125 95879 6240
rect 95719 5728 95879 6125
rect 95719 5696 95723 5728
rect 95755 5696 95763 5728
rect 95795 5696 95803 5728
rect 95835 5696 95843 5728
rect 95875 5696 95879 5728
rect 95719 5184 95879 5696
rect 95719 5152 95723 5184
rect 95755 5152 95763 5184
rect 95795 5152 95803 5184
rect 95835 5152 95843 5184
rect 95875 5152 95879 5184
rect 95719 4787 95879 5152
rect 95719 4669 95740 4787
rect 95858 4669 95879 4787
rect 95719 4640 95879 4669
rect 95719 4608 95723 4640
rect 95755 4608 95763 4640
rect 95795 4608 95803 4640
rect 95835 4608 95843 4640
rect 95875 4608 95879 4640
rect 95719 4096 95879 4608
rect 95719 4064 95723 4096
rect 95755 4064 95763 4096
rect 95795 4064 95803 4096
rect 95835 4064 95843 4096
rect 95875 4064 95879 4096
rect 95719 3552 95879 4064
rect 95719 3520 95723 3552
rect 95755 3520 95763 3552
rect 95795 3520 95803 3552
rect 95835 3520 95843 3552
rect 95875 3520 95879 3552
rect 95719 3331 95879 3520
rect 95719 3213 95740 3331
rect 95858 3213 95879 3331
rect 95719 3008 95879 3213
rect 95719 2976 95723 3008
rect 95755 2976 95763 3008
rect 95795 2976 95803 3008
rect 95835 2976 95843 3008
rect 95875 2976 95879 3008
rect 95719 2464 95879 2976
rect 95719 2432 95723 2464
rect 95755 2432 95763 2464
rect 95795 2432 95803 2464
rect 95835 2432 95843 2464
rect 95875 2432 95879 2464
rect 95719 1920 95879 2432
rect 95719 1888 95723 1920
rect 95755 1888 95763 1920
rect 95795 1888 95803 1920
rect 95835 1888 95843 1920
rect 95875 1888 95879 1920
rect 95719 1875 95879 1888
rect 95719 1757 95740 1875
rect 95858 1757 95879 1875
rect 95719 1376 95879 1757
rect 95719 1344 95723 1376
rect 95755 1344 95763 1376
rect 95795 1344 95803 1376
rect 95835 1344 95843 1376
rect 95875 1344 95879 1376
rect 95719 467 95879 1344
rect 95719 349 95740 467
rect 95858 349 95879 467
rect 95719 -2 95879 349
rect 114769 7869 114929 7890
rect 114769 7751 114790 7869
rect 114908 7751 114929 7869
rect 114769 6544 114929 7751
rect 114769 6512 114773 6544
rect 114805 6512 114813 6544
rect 114845 6512 114853 6544
rect 114885 6512 114893 6544
rect 114925 6512 114929 6544
rect 114769 6000 114929 6512
rect 114769 5968 114773 6000
rect 114805 5968 114813 6000
rect 114845 5968 114853 6000
rect 114885 5968 114893 6000
rect 114925 5968 114929 6000
rect 114769 5515 114929 5968
rect 114769 5456 114790 5515
rect 114908 5456 114929 5515
rect 114769 5424 114773 5456
rect 114925 5424 114929 5456
rect 114769 5397 114790 5424
rect 114908 5397 114929 5424
rect 114769 4912 114929 5397
rect 114769 4880 114773 4912
rect 114805 4880 114813 4912
rect 114845 4880 114853 4912
rect 114885 4880 114893 4912
rect 114925 4880 114929 4912
rect 114769 4368 114929 4880
rect 114769 4336 114773 4368
rect 114805 4336 114813 4368
rect 114845 4336 114853 4368
rect 114885 4336 114893 4368
rect 114925 4336 114929 4368
rect 114769 4059 114929 4336
rect 114769 3941 114790 4059
rect 114908 3941 114929 4059
rect 114769 3824 114929 3941
rect 114769 3792 114773 3824
rect 114805 3792 114813 3824
rect 114845 3792 114853 3824
rect 114885 3792 114893 3824
rect 114925 3792 114929 3824
rect 114769 3280 114929 3792
rect 114769 3248 114773 3280
rect 114805 3248 114813 3280
rect 114845 3248 114853 3280
rect 114885 3248 114893 3280
rect 114925 3248 114929 3280
rect 114769 2736 114929 3248
rect 114769 2704 114773 2736
rect 114805 2704 114813 2736
rect 114845 2704 114853 2736
rect 114885 2704 114893 2736
rect 114925 2704 114929 2736
rect 114769 2603 114929 2704
rect 114769 2485 114790 2603
rect 114908 2485 114929 2603
rect 114769 2192 114929 2485
rect 114769 2160 114773 2192
rect 114805 2160 114813 2192
rect 114845 2160 114853 2192
rect 114885 2160 114893 2192
rect 114925 2160 114929 2192
rect 114769 1648 114929 2160
rect 114769 1616 114773 1648
rect 114805 1616 114813 1648
rect 114845 1616 114853 1648
rect 114885 1616 114893 1648
rect 114925 1616 114929 1648
rect 114769 1104 114929 1616
rect 114769 1072 114773 1104
rect 114805 1072 114813 1104
rect 114845 1072 114853 1104
rect 114885 1072 114893 1104
rect 114925 1072 114929 1104
rect 114769 137 114929 1072
rect 114769 19 114790 137
rect 114908 19 114929 137
rect 114769 -2 114929 19
rect 133818 7539 133978 7890
rect 153834 7869 153994 7890
rect 153834 7751 153855 7869
rect 153973 7751 153994 7869
rect 133818 7421 133839 7539
rect 133957 7421 133978 7539
rect 133818 6816 133978 7421
rect 133818 6784 133822 6816
rect 133854 6784 133862 6816
rect 133894 6784 133902 6816
rect 133934 6784 133942 6816
rect 133974 6784 133978 6816
rect 133818 6272 133978 6784
rect 133818 6240 133822 6272
rect 133854 6243 133862 6272
rect 133894 6243 133902 6272
rect 133934 6243 133942 6272
rect 133974 6240 133978 6272
rect 133818 6125 133839 6240
rect 133957 6125 133978 6240
rect 133818 5728 133978 6125
rect 133818 5696 133822 5728
rect 133854 5696 133862 5728
rect 133894 5696 133902 5728
rect 133934 5696 133942 5728
rect 133974 5696 133978 5728
rect 133818 5184 133978 5696
rect 133818 5152 133822 5184
rect 133854 5152 133862 5184
rect 133894 5152 133902 5184
rect 133934 5152 133942 5184
rect 133974 5152 133978 5184
rect 133818 4787 133978 5152
rect 133818 4669 133839 4787
rect 133957 4669 133978 4787
rect 133818 4640 133978 4669
rect 133818 4608 133822 4640
rect 133854 4608 133862 4640
rect 133894 4608 133902 4640
rect 133934 4608 133942 4640
rect 133974 4608 133978 4640
rect 133818 4096 133978 4608
rect 133818 4064 133822 4096
rect 133854 4064 133862 4096
rect 133894 4064 133902 4096
rect 133934 4064 133942 4096
rect 133974 4064 133978 4096
rect 133818 3552 133978 4064
rect 133818 3520 133822 3552
rect 133854 3520 133862 3552
rect 133894 3520 133902 3552
rect 133934 3520 133942 3552
rect 133974 3520 133978 3552
rect 133818 3331 133978 3520
rect 133818 3213 133839 3331
rect 133957 3213 133978 3331
rect 133818 3008 133978 3213
rect 133818 2976 133822 3008
rect 133854 2976 133862 3008
rect 133894 2976 133902 3008
rect 133934 2976 133942 3008
rect 133974 2976 133978 3008
rect 133818 2464 133978 2976
rect 133818 2432 133822 2464
rect 133854 2432 133862 2464
rect 133894 2432 133902 2464
rect 133934 2432 133942 2464
rect 133974 2432 133978 2464
rect 133818 1920 133978 2432
rect 133818 1888 133822 1920
rect 133854 1888 133862 1920
rect 133894 1888 133902 1920
rect 133934 1888 133942 1920
rect 133974 1888 133978 1920
rect 133818 1875 133978 1888
rect 133818 1757 133839 1875
rect 133957 1757 133978 1875
rect 133818 1376 133978 1757
rect 133818 1344 133822 1376
rect 133854 1344 133862 1376
rect 133894 1344 133902 1376
rect 133934 1344 133942 1376
rect 133974 1344 133978 1376
rect 133818 467 133978 1344
rect 133818 349 133839 467
rect 133957 349 133978 467
rect 133818 -2 133978 349
rect 153504 7539 153664 7560
rect 153504 7421 153525 7539
rect 153643 7421 153664 7539
rect 153504 6243 153664 7421
rect 153504 6125 153525 6243
rect 153643 6125 153664 6243
rect 153504 4787 153664 6125
rect 153504 4669 153525 4787
rect 153643 4669 153664 4787
rect 153504 3331 153664 4669
rect 153504 3213 153525 3331
rect 153643 3213 153664 3331
rect 153504 1875 153664 3213
rect 153504 1757 153525 1875
rect 153643 1757 153664 1875
rect 153504 467 153664 1757
rect 153504 349 153525 467
rect 153643 349 153664 467
rect 153504 328 153664 349
rect 153834 5515 153994 7751
rect 153834 5397 153855 5515
rect 153973 5397 153994 5515
rect 153834 4059 153994 5397
rect 153834 3941 153855 4059
rect 153973 3941 153994 4059
rect 153834 2603 153994 3941
rect 153834 2485 153855 2603
rect 153973 2485 153994 2603
rect 153834 137 153994 2485
rect 153834 19 153855 137
rect 153973 19 153994 137
rect 153834 -2 153994 19
<< via4 >>
rect -517 7751 -399 7869
rect -517 5397 -399 5515
rect -517 3941 -399 4059
rect -517 2485 -399 2603
rect -187 7421 -69 7539
rect -187 6125 -69 6243
rect -187 4669 -69 4787
rect -187 3213 -69 3331
rect -187 1757 -69 1875
rect -187 349 -69 467
rect 19542 7421 19660 7539
rect 19542 6240 19557 6243
rect 19557 6240 19565 6243
rect 19565 6240 19597 6243
rect 19597 6240 19605 6243
rect 19605 6240 19637 6243
rect 19637 6240 19645 6243
rect 19645 6240 19660 6243
rect 19542 6125 19660 6240
rect 19542 4669 19660 4787
rect 19542 3213 19660 3331
rect 19542 1757 19660 1875
rect 19542 349 19660 467
rect -517 19 -399 137
rect 38592 7751 38710 7869
rect 38592 5456 38710 5515
rect 38592 5424 38607 5456
rect 38607 5424 38615 5456
rect 38615 5424 38647 5456
rect 38647 5424 38655 5456
rect 38655 5424 38687 5456
rect 38687 5424 38695 5456
rect 38695 5424 38710 5456
rect 38592 5397 38710 5424
rect 38592 3941 38710 4059
rect 38592 2485 38710 2603
rect 38592 19 38710 137
rect 57641 7421 57759 7539
rect 57641 6240 57656 6243
rect 57656 6240 57664 6243
rect 57664 6240 57696 6243
rect 57696 6240 57704 6243
rect 57704 6240 57736 6243
rect 57736 6240 57744 6243
rect 57744 6240 57759 6243
rect 57641 6125 57759 6240
rect 57641 4669 57759 4787
rect 57641 3213 57759 3331
rect 57641 1757 57759 1875
rect 57641 349 57759 467
rect 76691 7751 76809 7869
rect 76691 5456 76809 5515
rect 76691 5424 76706 5456
rect 76706 5424 76714 5456
rect 76714 5424 76746 5456
rect 76746 5424 76754 5456
rect 76754 5424 76786 5456
rect 76786 5424 76794 5456
rect 76794 5424 76809 5456
rect 76691 5397 76809 5424
rect 76691 3941 76809 4059
rect 76691 2485 76809 2603
rect 76691 19 76809 137
rect 95740 7421 95858 7539
rect 95740 6240 95755 6243
rect 95755 6240 95763 6243
rect 95763 6240 95795 6243
rect 95795 6240 95803 6243
rect 95803 6240 95835 6243
rect 95835 6240 95843 6243
rect 95843 6240 95858 6243
rect 95740 6125 95858 6240
rect 95740 4669 95858 4787
rect 95740 3213 95858 3331
rect 95740 1757 95858 1875
rect 95740 349 95858 467
rect 114790 7751 114908 7869
rect 114790 5456 114908 5515
rect 114790 5424 114805 5456
rect 114805 5424 114813 5456
rect 114813 5424 114845 5456
rect 114845 5424 114853 5456
rect 114853 5424 114885 5456
rect 114885 5424 114893 5456
rect 114893 5424 114908 5456
rect 114790 5397 114908 5424
rect 114790 3941 114908 4059
rect 114790 2485 114908 2603
rect 114790 19 114908 137
rect 153855 7751 153973 7869
rect 133839 7421 133957 7539
rect 133839 6240 133854 6243
rect 133854 6240 133862 6243
rect 133862 6240 133894 6243
rect 133894 6240 133902 6243
rect 133902 6240 133934 6243
rect 133934 6240 133942 6243
rect 133942 6240 133957 6243
rect 133839 6125 133957 6240
rect 133839 4669 133957 4787
rect 133839 3213 133957 3331
rect 133839 1757 133957 1875
rect 133839 349 133957 467
rect 153525 7421 153643 7539
rect 153525 6125 153643 6243
rect 153525 4669 153643 4787
rect 153525 3213 153643 3331
rect 153525 1757 153643 1875
rect 153525 349 153643 467
rect 153855 5397 153973 5515
rect 153855 3941 153973 4059
rect 153855 2485 153973 2603
rect 153855 19 153973 137
<< metal5 >>
rect -538 7869 153994 7890
rect -538 7751 -517 7869
rect -399 7751 38592 7869
rect 38710 7751 76691 7869
rect 76809 7751 114790 7869
rect 114908 7751 153855 7869
rect 153973 7751 153994 7869
rect -538 7730 153994 7751
rect -208 7539 153664 7560
rect -208 7421 -187 7539
rect -69 7421 19542 7539
rect 19660 7421 57641 7539
rect 57759 7421 95740 7539
rect 95858 7421 133839 7539
rect 133957 7421 153525 7539
rect 153643 7421 153664 7539
rect -208 7400 153664 7421
rect -538 6243 153994 6264
rect -538 6125 -187 6243
rect -69 6125 19542 6243
rect 19660 6125 57641 6243
rect 57759 6125 95740 6243
rect 95858 6125 133839 6243
rect 133957 6125 153525 6243
rect 153643 6125 153994 6243
rect -538 6104 153994 6125
rect -538 5515 153994 5536
rect -538 5397 -517 5515
rect -399 5397 38592 5515
rect 38710 5397 76691 5515
rect 76809 5397 114790 5515
rect 114908 5397 153855 5515
rect 153973 5397 153994 5515
rect -538 5376 153994 5397
rect -538 4787 153994 4808
rect -538 4669 -187 4787
rect -69 4669 19542 4787
rect 19660 4669 57641 4787
rect 57759 4669 95740 4787
rect 95858 4669 133839 4787
rect 133957 4669 153525 4787
rect 153643 4669 153994 4787
rect -538 4648 153994 4669
rect -538 4059 153994 4080
rect -538 3941 -517 4059
rect -399 3941 38592 4059
rect 38710 3941 76691 4059
rect 76809 3941 114790 4059
rect 114908 3941 153855 4059
rect 153973 3941 153994 4059
rect -538 3920 153994 3941
rect -538 3331 153994 3352
rect -538 3213 -187 3331
rect -69 3213 19542 3331
rect 19660 3213 57641 3331
rect 57759 3213 95740 3331
rect 95858 3213 133839 3331
rect 133957 3213 153525 3331
rect 153643 3213 153994 3331
rect -538 3192 153994 3213
rect -538 2603 153994 2624
rect -538 2485 -517 2603
rect -399 2485 38592 2603
rect 38710 2485 76691 2603
rect 76809 2485 114790 2603
rect 114908 2485 153855 2603
rect 153973 2485 153994 2603
rect -538 2464 153994 2485
rect -538 1875 153994 1896
rect -538 1757 -187 1875
rect -69 1757 19542 1875
rect 19660 1757 57641 1875
rect 57759 1757 95740 1875
rect 95858 1757 133839 1875
rect 133957 1757 153525 1875
rect 153643 1757 153994 1875
rect -538 1736 153994 1757
rect -208 467 153664 488
rect -208 349 -187 467
rect -69 349 19542 467
rect 19660 349 57641 467
rect 57759 349 95740 467
rect 95858 349 133839 467
rect 133957 349 153525 467
rect 153643 349 153664 467
rect -208 328 153664 349
rect -538 137 153994 158
rect -538 19 -517 137
rect -399 19 38592 137
rect 38710 19 76691 137
rect 76809 19 114790 137
rect 114908 19 153855 137
rect 153973 19 153994 137
rect -538 -2 153994 19
use sky130_fd_sc_hd__buf_4  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 68862 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__clkbuf_2  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 28474 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 29072 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 28106 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1712078602
transform 1 0 28060 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1712078602
transform 1 0 28980 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1712078602
transform 1 0 27462 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1712078602
transform 1 0 27646 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1712078602
transform 1 0 26772 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp 1712078602
transform 1 0 25990 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1712078602
transform 1 0 25484 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1712078602
transform 1 0 26404 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _360_
timestamp 1712078602
transform 1 0 21804 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1712078602
transform 1 0 21528 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1712078602
transform 1 0 20838 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1712078602
transform 1 0 22494 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1712078602
transform 1 0 20792 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1712078602
transform 1 0 20102 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1712078602
transform 1 0 20148 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1712078602
transform 1 0 19826 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1712078602
transform 1 0 19504 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1712078602
transform 1 0 18998 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1712078602
transform 1 0 19228 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1712078602
transform 1 0 18492 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1712078602
transform 1 0 17158 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1712078602
transform 1 0 16974 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1712078602
transform 1 0 16054 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1712078602
transform 1 0 16376 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1712078602
transform 1 0 15916 0 1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1712078602
transform 1 0 16698 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1712078602
transform 1 0 14306 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1712078602
transform 1 0 17480 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1712078602
transform 1 0 15134 0 -1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1712078602
transform 1 0 16054 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _382_
timestamp 1712078602
transform 1 0 18124 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1712078602
transform 1 0 14122 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1712078602
transform 1 0 15456 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1712078602
transform 1 0 14214 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1712078602
transform 1 0 14812 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1712078602
transform 1 0 12834 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1712078602
transform 1 0 14398 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1712078602
transform 1 0 13524 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _390_
timestamp 1712078602
transform 1 0 15134 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1712078602
transform 1 0 13708 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _392_
timestamp 1712078602
transform 1 0 15548 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_4  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 72864 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1712078602
transform 1 0 77234 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp 1712078602
transform 1 0 75394 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1712078602
transform 1 0 97750 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _397_
timestamp 1712078602
transform 1 0 94254 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1712078602
transform 1 0 97198 0 1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1712078602
transform 1 0 96554 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1712078602
transform 1 0 98486 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1712078602
transform 1 0 96140 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1712078602
transform 1 0 99084 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1712078602
transform 1 0 98118 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _404_
timestamp 1712078602
transform 1 0 124476 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__clkbuf_2  _405_
timestamp 1712078602
transform 1 0 131192 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1712078602
transform 1 0 134412 0 1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1712078602
transform 1 0 133860 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1712078602
transform 1 0 136252 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1712078602
transform 1 0 134182 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1712078602
transform 1 0 135838 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1712078602
transform 1 0 133538 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1712078602
transform 1 0 135010 0 1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1712078602
transform 1 0 133860 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1712078602
transform 1 0 135654 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1712078602
transform 1 0 133998 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _416_
timestamp 1712078602
transform 1 0 130870 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1712078602
transform 1 0 133906 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 1712078602
transform 1 0 132894 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1712078602
transform 1 0 133400 0 1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1712078602
transform 1 0 132480 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1712078602
transform 1 0 133722 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1712078602
transform 1 0 131974 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1712078602
transform 1 0 132618 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1712078602
transform 1 0 132296 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1712078602
transform 1 0 131330 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1712078602
transform 1 0 132296 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _427_
timestamp 1712078602
transform 1 0 125902 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1712078602
transform 1 0 127926 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1712078602
transform 1 0 126822 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _430_
timestamp 1712078602
transform 1 0 127374 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _431_
timestamp 1712078602
transform 1 0 126868 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1712078602
transform 1 0 126822 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1712078602
transform 1 0 126546 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1712078602
transform 1 0 125994 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1712078602
transform 1 0 125902 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1712078602
transform 1 0 124752 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1712078602
transform 1 0 125534 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _438_
timestamp 1712078602
transform 1 0 121854 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1712078602
transform 1 0 121164 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1712078602
transform 1 0 121762 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _441_
timestamp 1712078602
transform 1 0 120428 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1712078602
transform 1 0 120704 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1712078602
transform 1 0 119922 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1712078602
transform 1 0 120520 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 1712078602
transform 1 0 119370 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _446_
timestamp 1712078602
transform 1 0 119968 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1712078602
transform 1 0 118358 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1712078602
transform 1 0 118404 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _449_
timestamp 1712078602
transform 1 0 119278 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _450_
timestamp 1712078602
transform 1 0 115460 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _451_
timestamp 1712078602
transform 1 0 115782 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1712078602
transform 1 0 114540 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _453_
timestamp 1712078602
transform 1 0 114586 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1712078602
transform 1 0 113942 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _455_
timestamp 1712078602
transform 1 0 115046 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1712078602
transform 1 0 113298 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _457_
timestamp 1712078602
transform 1 0 113574 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1712078602
transform 1 0 111826 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _459_
timestamp 1712078602
transform 1 0 113252 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _460_
timestamp 1712078602
transform 1 0 82892 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__clkbuf_2  _461_
timestamp 1712078602
transform 1 0 96692 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1712078602
transform 1 0 103638 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _463_
timestamp 1712078602
transform 1 0 101062 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _464_
timestamp 1712078602
transform 1 0 102396 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _465_
timestamp 1712078602
transform 1 0 101430 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1712078602
transform 1 0 101798 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _467_
timestamp 1712078602
transform 1 0 99912 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1712078602
transform 1 0 101430 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp 1712078602
transform 1 0 101430 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 1712078602
transform 1 0 100234 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _471_
timestamp 1712078602
transform 1 0 100832 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _472_
timestamp 1712078602
transform 1 0 94622 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1712078602
transform 1 0 98486 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _474_
timestamp 1712078602
transform 1 0 96232 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1712078602
transform 1 0 96508 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _476_
timestamp 1712078602
transform 1 0 94714 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 1712078602
transform 1 0 95266 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _478_
timestamp 1712078602
transform 1 0 95542 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _479_
timestamp 1712078602
transform 1 0 95910 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp 1712078602
transform 1 0 95910 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1712078602
transform 1 0 93978 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp 1712078602
transform 1 0 95082 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _483_
timestamp 1712078602
transform 1 0 87768 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _484_
timestamp 1712078602
transform 1 0 90758 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp 1712078602
transform 1 0 89470 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _486_
timestamp 1712078602
transform 1 0 89378 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _487_
timestamp 1712078602
transform 1 0 90390 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _488_
timestamp 1712078602
transform 1 0 88780 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _489_
timestamp 1712078602
transform 1 0 87492 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _490_
timestamp 1712078602
transform 1 0 88274 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _491_
timestamp 1712078602
transform 1 0 88228 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 1712078602
transform 1 0 86894 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _493_
timestamp 1712078602
transform 1 0 87814 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _494_
timestamp 1712078602
transform 1 0 83628 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _495_
timestamp 1712078602
transform 1 0 83030 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp 1712078602
transform 1 0 81328 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _497_
timestamp 1712078602
transform 1 0 82018 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp 1712078602
transform 1 0 81742 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _499_
timestamp 1712078602
transform 1 0 81006 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _500_
timestamp 1712078602
transform 1 0 81006 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _501_
timestamp 1712078602
transform 1 0 80408 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _502_
timestamp 1712078602
transform 1 0 80454 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _503_
timestamp 1712078602
transform 1 0 79396 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1712078602
transform 1 0 79994 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _505_
timestamp 1712078602
transform 1 0 80546 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _506_
timestamp 1712078602
transform 1 0 76636 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _507_
timestamp 1712078602
transform 1 0 77050 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _508_
timestamp 1712078602
transform 1 0 75532 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _509_
timestamp 1712078602
transform 1 0 75532 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _510_
timestamp 1712078602
transform 1 0 75808 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _511_
timestamp 1712078602
transform 1 0 74428 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _512_
timestamp 1712078602
transform 1 0 74014 0 1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _513_
timestamp 1712078602
transform 1 0 73646 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _514_
timestamp 1712078602
transform 1 0 72726 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _515_
timestamp 1712078602
transform 1 0 73784 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__buf_2  _516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 65826 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__clkbuf_2  _517_
timestamp 1712078602
transform 1 0 62698 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _518_
timestamp 1712078602
transform 1 0 66562 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1712078602
transform 1 0 65872 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _520_
timestamp 1712078602
transform 1 0 65642 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1712078602
transform 1 0 66194 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 1712078602
transform 1 0 65228 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1712078602
transform 1 0 64032 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _524_
timestamp 1712078602
transform 1 0 64354 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1712078602
transform 1 0 64216 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _526_
timestamp 1712078602
transform 1 0 63066 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1712078602
transform 1 0 63848 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _528_
timestamp 1712078602
transform 1 0 56856 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _529_
timestamp 1712078602
transform 1 0 59846 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp 1712078602
transform 1 0 58558 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _531_
timestamp 1712078602
transform 1 0 58558 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1712078602
transform 1 0 58098 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _533_
timestamp 1712078602
transform 1 0 57638 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp 1712078602
transform 1 0 58006 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _535_
timestamp 1712078602
transform 1 0 57316 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _536_
timestamp 1712078602
transform 1 0 56902 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _537_
timestamp 1712078602
transform 1 0 55936 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _538_
timestamp 1712078602
transform 1 0 56534 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _539_
timestamp 1712078602
transform 1 0 51014 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1712078602
transform 1 0 52118 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1712078602
transform 1 0 51474 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _542_
timestamp 1712078602
transform 1 0 51290 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1712078602
transform 1 0 51750 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _544_
timestamp 1712078602
transform 1 0 50738 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1712078602
transform 1 0 50830 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _546_
timestamp 1712078602
transform 1 0 50186 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1712078602
transform 1 0 50094 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _548_
timestamp 1712078602
transform 1 0 48760 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1712078602
transform 1 0 49542 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _550_
timestamp 1712078602
transform 1 0 45172 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1712078602
transform 1 0 44574 0 -1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1712078602
transform 1 0 44114 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1712078602
transform 1 0 43792 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1712078602
transform 1 0 43792 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1712078602
transform 1 0 43194 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1712078602
transform 1 0 41446 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1712078602
transform 1 0 42826 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1712078602
transform 1 0 43102 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1712078602
transform 1 0 41998 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1712078602
transform 1 0 42504 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _561_
timestamp 1712078602
transform 1 0 43838 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__mux2_1  _562_
timestamp 1712078602
transform 1 0 40526 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1712078602
transform 1 0 39560 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _564_
timestamp 1712078602
transform 1 0 38732 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1712078602
transform 1 0 39100 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _566_
timestamp 1712078602
transform 1 0 38134 0 1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1712078602
transform 1 0 38456 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _568_
timestamp 1712078602
transform 1 0 37766 0 -1 5984
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1712078602
transform 1 0 37444 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__mux2_1  _570_
timestamp 1712078602
transform 1 0 36018 0 1 6528
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1712078602
transform 1 0 38226 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__buf_2  _572_
timestamp 1712078602
transform 1 0 67666 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__buf_2  _573_
timestamp 1712078602
transform 1 0 43470 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 38870 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1712078602
transform 1 0 38870 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1712078602
transform 1 0 39238 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1712078602
transform 1 0 39606 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1712078602
transform 1 0 40066 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _579_
timestamp 1712078602
transform 1 0 45862 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1712078602
transform 1 0 43424 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1712078602
transform 1 0 42734 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1712078602
transform 1 0 45034 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1712078602
transform 1 0 44390 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1712078602
transform 1 0 44390 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _585_
timestamp 1712078602
transform 1 0 50922 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1712078602
transform 1 0 49864 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1712078602
transform 1 0 50416 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1712078602
transform 1 0 52532 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _589_
timestamp 1712078602
transform 1 0 52210 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _590_
timestamp 1712078602
transform 1 0 51888 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _591_
timestamp 1712078602
transform 1 0 57270 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _592_
timestamp 1712078602
transform 1 0 57638 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1712078602
transform 1 0 56534 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _594_
timestamp 1712078602
transform 1 0 59156 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _595_
timestamp 1712078602
transform 1 0 58420 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _596_
timestamp 1712078602
transform 1 0 58742 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _597_
timestamp 1712078602
transform 1 0 63664 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _598_
timestamp 1712078602
transform 1 0 64630 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1712078602
transform 1 0 65182 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _600_
timestamp 1712078602
transform 1 0 65550 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _601_
timestamp 1712078602
transform 1 0 66286 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _602_
timestamp 1712078602
transform 1 0 65090 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _603_
timestamp 1712078602
transform 1 0 82616 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__buf_2  _604_
timestamp 1712078602
transform 1 0 79994 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _605_
timestamp 1712078602
transform 1 0 74152 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _606_
timestamp 1712078602
transform 1 0 75302 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1712078602
transform 1 0 74934 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1712078602
transform 1 0 76222 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _609_
timestamp 1712078602
transform 1 0 76314 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _610_
timestamp 1712078602
transform 1 0 83214 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _611_
timestamp 1712078602
transform 1 0 81098 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _612_
timestamp 1712078602
transform 1 0 81420 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _613_
timestamp 1712078602
transform 1 0 81742 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1712078602
transform 1 0 82386 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _615_
timestamp 1712078602
transform 1 0 82064 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _616_
timestamp 1712078602
transform 1 0 88918 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _617_
timestamp 1712078602
transform 1 0 88734 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1712078602
transform 1 0 89056 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _619_
timestamp 1712078602
transform 1 0 89976 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _620_
timestamp 1712078602
transform 1 0 90758 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _621_
timestamp 1712078602
transform 1 0 91080 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _622_
timestamp 1712078602
transform 1 0 94254 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _623_
timestamp 1712078602
transform 1 0 93656 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _624_
timestamp 1712078602
transform 1 0 95082 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1712078602
transform 1 0 97060 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1712078602
transform 1 0 96462 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _627_
timestamp 1712078602
transform 1 0 98348 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__buf_2  _628_
timestamp 1712078602
transform 1 0 96324 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _629_
timestamp 1712078602
transform 1 0 101108 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1712078602
transform 1 0 101384 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1712078602
transform 1 0 101706 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1712078602
transform 1 0 100510 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1712078602
transform 1 0 100234 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _634_
timestamp 1712078602
transform 1 0 126316 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__buf_2  _635_
timestamp 1712078602
transform 1 0 119002 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _636_
timestamp 1712078602
transform 1 0 116518 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1712078602
transform 1 0 115138 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1712078602
transform 1 0 115460 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1712078602
transform 1 0 116058 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1712078602
transform 1 0 116518 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _641_
timestamp 1712078602
transform 1 0 122222 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1712078602
transform 1 0 119922 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _643_
timestamp 1712078602
transform 1 0 120382 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _644_
timestamp 1712078602
transform 1 0 120842 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _645_
timestamp 1712078602
transform 1 0 121026 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _646_
timestamp 1712078602
transform 1 0 122590 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _647_
timestamp 1712078602
transform 1 0 125626 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _648_
timestamp 1712078602
transform 1 0 126224 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _649_
timestamp 1712078602
transform 1 0 127420 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _650_
timestamp 1712078602
transform 1 0 127742 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1712078602
transform 1 0 128524 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1712078602
transform 1 0 128110 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _653_
timestamp 1712078602
transform 1 0 130824 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _654_
timestamp 1712078602
transform 1 0 131974 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _655_
timestamp 1712078602
transform 1 0 133216 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _656_
timestamp 1712078602
transform 1 0 132158 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _657_
timestamp 1712078602
transform 1 0 132434 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1712078602
transform 1 0 133538 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _659_
timestamp 1712078602
transform 1 0 131560 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _660_
timestamp 1712078602
transform 1 0 135470 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _661_
timestamp 1712078602
transform 1 0 134182 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _662_
timestamp 1712078602
transform 1 0 134550 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _663_
timestamp 1712078602
transform 1 0 133906 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1712078602
transform 1 0 135654 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__buf_4  _665_
timestamp 1712078602
transform 1 0 71484 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__clkbuf_4  _666_
timestamp 1712078602
transform 1 0 74750 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__inv_2  _667_
timestamp 1712078602
transform 1 0 94760 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _668_
timestamp 1712078602
transform 1 0 95404 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _669_
timestamp 1712078602
transform 1 0 95036 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _670_
timestamp 1712078602
transform 1 0 95358 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _671_
timestamp 1712078602
transform 1 0 78200 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _672_
timestamp 1712078602
transform 1 0 18216 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _673_
timestamp 1712078602
transform 1 0 15778 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _674_
timestamp 1712078602
transform 1 0 16054 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _675_
timestamp 1712078602
transform 1 0 16744 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _676_
timestamp 1712078602
transform 1 0 16376 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _677_
timestamp 1712078602
transform 1 0 16100 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _678_
timestamp 1712078602
transform 1 0 18630 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _679_
timestamp 1712078602
transform 1 0 16744 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _680_
timestamp 1712078602
transform 1 0 17664 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _681_
timestamp 1712078602
transform 1 0 17158 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _682_
timestamp 1712078602
transform 1 0 16836 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1712078602
transform 1 0 17342 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _684_
timestamp 1712078602
transform 1 0 21390 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _685_
timestamp 1712078602
transform 1 0 19550 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _686_
timestamp 1712078602
transform 1 0 20470 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _687_
timestamp 1712078602
transform 1 0 20516 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _688_
timestamp 1712078602
transform 1 0 20838 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _689_
timestamp 1712078602
transform 1 0 21206 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_2  _690_
timestamp 1712078602
transform 1 0 27692 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  _691_
timestamp 1712078602
transform 1 0 26450 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _692_
timestamp 1712078602
transform 1 0 27140 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _693_
timestamp 1712078602
transform 1 0 27278 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _694_
timestamp 1712078602
transform 1 0 28198 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  _695_
timestamp 1712078602
transform 1 0 28520 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__dfrtp_1  _696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 36800 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _697_
timestamp 1712078602
transform 1 0 37766 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _698_
timestamp 1712078602
transform 1 0 38088 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _699_
timestamp 1712078602
transform 1 0 39238 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _700_
timestamp 1712078602
transform 1 0 39882 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _701_
timestamp 1712078602
transform 1 0 41998 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _702_
timestamp 1712078602
transform 1 0 41952 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _703_
timestamp 1712078602
transform 1 0 43102 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _704_
timestamp 1712078602
transform 1 0 43240 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _705_
timestamp 1712078602
transform 1 0 44390 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _706_
timestamp 1712078602
transform 1 0 49588 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _707_
timestamp 1712078602
transform 1 0 49680 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _708_
timestamp 1712078602
transform 1 0 50692 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _709_
timestamp 1712078602
transform 1 0 50968 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _710_
timestamp 1712078602
transform 1 0 52118 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _711_
timestamp 1712078602
transform 1 0 56120 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _712_
timestamp 1712078602
transform 1 0 57178 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _713_
timestamp 1712078602
transform 1 0 57408 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _714_
timestamp 1712078602
transform 1 0 58236 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _715_
timestamp 1712078602
transform 1 0 58696 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _716_
timestamp 1712078602
transform 1 0 63756 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _717_
timestamp 1712078602
transform 1 0 64538 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _718_
timestamp 1712078602
transform 1 0 65136 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _719_
timestamp 1712078602
transform 1 0 65412 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _720_
timestamp 1712078602
transform 1 0 66286 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _721_
timestamp 1712078602
transform 1 0 72864 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _722_
timestamp 1712078602
transform 1 0 73738 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _723_
timestamp 1712078602
transform 1 0 74152 0 -1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _724_
timestamp 1712078602
transform 1 0 75440 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _725_
timestamp 1712078602
transform 1 0 76728 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _726_
timestamp 1712078602
transform 1 0 79304 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _727_
timestamp 1712078602
transform 1 0 80454 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _728_
timestamp 1712078602
transform 1 0 80914 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _729_
timestamp 1712078602
transform 1 0 81742 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _730_
timestamp 1712078602
transform 1 0 81788 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _731_
timestamp 1712078602
transform 1 0 88182 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _732_
timestamp 1712078602
transform 1 0 88182 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _733_
timestamp 1712078602
transform 1 0 89470 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _734_
timestamp 1712078602
transform 1 0 89286 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _735_
timestamp 1712078602
transform 1 0 89562 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _736_
timestamp 1712078602
transform 1 0 94760 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _737_
timestamp 1712078602
transform 1 0 95404 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _738_
timestamp 1712078602
transform 1 0 95910 0 -1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _739_
timestamp 1712078602
transform 1 0 96002 0 1 5440
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _740_
timestamp 1712078602
transform 1 0 97014 0 -1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _741_
timestamp 1712078602
transform 1 0 101062 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _742_
timestamp 1712078602
transform 1 0 101292 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _743_
timestamp 1712078602
transform 1 0 102350 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _744_
timestamp 1712078602
transform 1 0 102396 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _745_
timestamp 1712078602
transform 1 0 102350 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _746_
timestamp 1712078602
transform 1 0 113942 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _747_
timestamp 1712078602
transform 1 0 113942 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _748_
timestamp 1712078602
transform 1 0 113758 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _749_
timestamp 1712078602
transform 1 0 115230 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _750_
timestamp 1712078602
transform 1 0 115368 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _751_
timestamp 1712078602
transform 1 0 119094 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _752_
timestamp 1712078602
transform 1 0 119232 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _753_
timestamp 1712078602
transform 1 0 120382 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _754_
timestamp 1712078602
transform 1 0 120336 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _755_
timestamp 1712078602
transform 1 0 121670 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _756_
timestamp 1712078602
transform 1 0 125534 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _757_
timestamp 1712078602
transform 1 0 126822 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _758_
timestamp 1712078602
transform 1 0 126270 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _759_
timestamp 1712078602
transform 1 0 126822 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _760_
timestamp 1712078602
transform 1 0 128110 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _761_
timestamp 1712078602
transform 1 0 132112 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _762_
timestamp 1712078602
transform 1 0 132618 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _763_
timestamp 1712078602
transform 1 0 132802 0 -1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _764_
timestamp 1712078602
transform 1 0 133262 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _765_
timestamp 1712078602
transform 1 0 134550 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _766_
timestamp 1712078602
transform 1 0 134550 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _767_
timestamp 1712078602
transform 1 0 134366 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _768_
timestamp 1712078602
transform 1 0 135838 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _769_
timestamp 1712078602
transform 1 0 134550 0 -1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_4  _770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 133262 0 1 6528
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrtp_4  _771_
timestamp 1712078602
transform 1 0 97198 0 1 5984
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrtp_4  _772_
timestamp 1712078602
transform 1 0 97198 0 1 6528
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrtp_4  _773_
timestamp 1712078602
transform 1 0 95910 0 1 6528
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrtp_4  _774_
timestamp 1712078602
transform 1 0 96508 0 -1 6528
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrtp_4  _775_
timestamp 1712078602
transform 1 0 74014 0 1 6528
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrtp_1  _776_
timestamp 1712078602
transform 1 0 14812 0 1 5440
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _777_
timestamp 1712078602
transform 1 0 13616 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _778_
timestamp 1712078602
transform 1 0 14812 0 -1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _779_
timestamp 1712078602
transform 1 0 14766 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _780_
timestamp 1712078602
transform 1 0 14904 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _781_
timestamp 1712078602
transform 1 0 14904 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _782_
timestamp 1712078602
transform 1 0 15870 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _783_
timestamp 1712078602
transform 1 0 16054 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _784_
timestamp 1712078602
transform 1 0 16192 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _785_
timestamp 1712078602
transform 1 0 17342 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _786_
timestamp 1712078602
transform 1 0 18768 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _787_
timestamp 1712078602
transform 1 0 19734 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _788_
timestamp 1712078602
transform 1 0 20056 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _789_
timestamp 1712078602
transform 1 0 20700 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _790_
timestamp 1712078602
transform 1 0 21252 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _791_
timestamp 1712078602
transform 1 0 26174 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _792_
timestamp 1712078602
transform 1 0 26496 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _793_
timestamp 1712078602
transform 1 0 27370 0 -1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _794_
timestamp 1712078602
transform 1 0 27784 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__dfrtp_1  _795_
timestamp 1712078602
transform 1 0 28934 0 1 6528
box -19 -24 939 296
use sky130_fd_sc_hd__buf_6  _796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 93564 0 -1 5440
box -19 -24 433 296
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform -1 0 21758 0 -1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1712078602
transform 1 0 27968 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1712078602
transform 1 0 77050 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1712078602
transform 1 0 76866 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1712078602
transform 1 0 77970 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1712078602
transform 1 0 76682 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1712078602
transform 1 0 78154 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1712078602
transform 1 0 76498 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1712078602
transform 1 0 78338 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1712078602
transform 1 0 76314 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1712078602
transform 1 0 78522 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1712078602
transform 1 0 76130 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1712078602
transform -1 0 151754 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1712078602
transform -1 0 151570 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1712078602
transform -1 0 151156 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1712078602
transform -1 0 150972 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1712078602
transform -1 0 150788 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1712078602
transform 1 0 152674 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1712078602
transform 1 0 152444 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1712078602
transform 1 0 152674 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1712078602
transform 1 0 152444 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1712078602
transform 1 0 152674 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1712078602
transform 1 0 920 0 -1 4352
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1712078602
transform 1 0 1104 0 -1 4352
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1712078602
transform 1 0 1288 0 -1 4352
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1712078602
transform 1 0 1472 0 -1 4352
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1712078602
transform 1 0 134228 0 1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1712078602
transform 1 0 126132 0 -1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1712078602
transform 1 0 98992 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1712078602
transform 1 0 98900 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1712078602
transform 1 0 147936 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 74704 0 1 5984
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1712078602
transform 1 0 70334 0 -1 5440
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1712078602
transform 1 0 70196 0 1 4896
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1712078602
transform 1 0 70196 0 1 5440
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1712078602
transform 1 0 70334 0 -1 4896
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1712078602
transform 1 0 78062 0 -1 5440
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1712078602
transform 1 0 78016 0 1 4896
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1712078602
transform 1 0 78016 0 1 5440
box -19 -24 939 296
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1712078602
transform 1 0 78062 0 -1 4896
box -19 -24 939 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 690 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1712078602
transform 1 0 1242 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 1794 0 1 1088
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1712078602
transform 1 0 1886 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1712078602
transform 1 0 2438 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 2990 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1712078602
transform 1 0 3174 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1712078602
transform 1 0 3726 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1712078602
transform 1 0 4278 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1712078602
transform 1 0 4462 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1712078602
transform 1 0 5014 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1712078602
transform 1 0 5566 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1712078602
transform 1 0 5750 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1712078602
transform 1 0 6302 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1712078602
transform 1 0 6854 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1712078602
transform 1 0 7038 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1712078602
transform 1 0 7590 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1712078602
transform 1 0 8142 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1712078602
transform 1 0 8326 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1712078602
transform 1 0 8878 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1712078602
transform 1 0 9430 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1712078602
transform 1 0 9614 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1712078602
transform 1 0 10166 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1712078602
transform 1 0 10718 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1712078602
transform 1 0 10902 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1712078602
transform 1 0 11454 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1712078602
transform 1 0 12006 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1712078602
transform 1 0 12190 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1712078602
transform 1 0 12742 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1712078602
transform 1 0 13294 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1712078602
transform 1 0 13478 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1712078602
transform 1 0 14030 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1712078602
transform 1 0 14582 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1712078602
transform 1 0 14766 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1712078602
transform 1 0 15318 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1712078602
transform 1 0 15870 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1712078602
transform 1 0 16054 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1712078602
transform 1 0 16606 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1712078602
transform 1 0 17158 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1712078602
transform 1 0 17342 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1712078602
transform 1 0 17894 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1712078602
transform 1 0 18446 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1712078602
transform 1 0 18630 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1712078602
transform 1 0 19182 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1712078602
transform 1 0 19734 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1712078602
transform 1 0 19918 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1712078602
transform 1 0 20470 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1712078602
transform 1 0 21022 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1712078602
transform 1 0 21206 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1712078602
transform 1 0 21758 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1712078602
transform 1 0 22310 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1712078602
transform 1 0 22494 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1712078602
transform 1 0 23046 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1712078602
transform 1 0 23598 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1712078602
transform 1 0 23782 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1712078602
transform 1 0 24334 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1712078602
transform 1 0 24886 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1712078602
transform 1 0 25070 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1712078602
transform 1 0 25622 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1712078602
transform 1 0 26174 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1712078602
transform 1 0 26358 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1712078602
transform 1 0 26910 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1712078602
transform 1 0 27462 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1712078602
transform 1 0 27646 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1712078602
transform 1 0 28198 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1712078602
transform 1 0 28750 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1712078602
transform 1 0 28934 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1712078602
transform 1 0 29486 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1712078602
transform 1 0 30038 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1712078602
transform 1 0 30222 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1712078602
transform 1 0 30774 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1712078602
transform 1 0 31326 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1712078602
transform 1 0 31510 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1712078602
transform 1 0 32062 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1712078602
transform 1 0 32614 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1712078602
transform 1 0 32798 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1712078602
transform 1 0 33350 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1712078602
transform 1 0 33902 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1712078602
transform 1 0 34086 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1712078602
transform 1 0 34638 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1712078602
transform 1 0 35190 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1712078602
transform 1 0 35374 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1712078602
transform 1 0 35926 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1712078602
transform 1 0 36478 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1712078602
transform 1 0 36662 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1712078602
transform 1 0 37214 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1712078602
transform 1 0 37766 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1712078602
transform 1 0 37950 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1712078602
transform 1 0 38502 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1712078602
transform 1 0 39054 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1712078602
transform 1 0 39238 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1712078602
transform 1 0 39790 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1712078602
transform 1 0 40342 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1712078602
transform 1 0 40526 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1712078602
transform 1 0 41078 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1712078602
transform 1 0 41630 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1712078602
transform 1 0 41814 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1712078602
transform 1 0 42366 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1712078602
transform 1 0 42918 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1712078602
transform 1 0 43102 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1712078602
transform 1 0 43654 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1712078602
transform 1 0 44206 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1712078602
transform 1 0 44390 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1712078602
transform 1 0 44942 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1712078602
transform 1 0 45494 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1712078602
transform 1 0 45678 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1712078602
transform 1 0 46230 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1712078602
transform 1 0 46782 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1712078602
transform 1 0 46966 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1712078602
transform 1 0 47518 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1712078602
transform 1 0 48070 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1712078602
transform 1 0 48254 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1712078602
transform 1 0 48806 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1712078602
transform 1 0 49358 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1712078602
transform 1 0 49542 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1712078602
transform 1 0 50094 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1712078602
transform 1 0 50646 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1712078602
transform 1 0 50830 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1712078602
transform 1 0 51382 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1712078602
transform 1 0 51934 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1712078602
transform 1 0 52118 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1712078602
transform 1 0 52670 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1712078602
transform 1 0 53222 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1712078602
transform 1 0 53406 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1161
timestamp 1712078602
transform 1 0 53958 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1712078602
transform 1 0 54510 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1177
timestamp 1712078602
transform 1 0 54694 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1189
timestamp 1712078602
transform 1 0 55246 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1712078602
transform 1 0 55798 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1205
timestamp 1712078602
transform 1 0 55982 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1217
timestamp 1712078602
transform 1 0 56534 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1229
timestamp 1712078602
transform 1 0 57086 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1233
timestamp 1712078602
transform 1 0 57270 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1245
timestamp 1712078602
transform 1 0 57822 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1257
timestamp 1712078602
transform 1 0 58374 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1261
timestamp 1712078602
transform 1 0 58558 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1273
timestamp 1712078602
transform 1 0 59110 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1285
timestamp 1712078602
transform 1 0 59662 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1289
timestamp 1712078602
transform 1 0 59846 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1301
timestamp 1712078602
transform 1 0 60398 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1313
timestamp 1712078602
transform 1 0 60950 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1317
timestamp 1712078602
transform 1 0 61134 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1329
timestamp 1712078602
transform 1 0 61686 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1341
timestamp 1712078602
transform 1 0 62238 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1345
timestamp 1712078602
transform 1 0 62422 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1357
timestamp 1712078602
transform 1 0 62974 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1369
timestamp 1712078602
transform 1 0 63526 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1373
timestamp 1712078602
transform 1 0 63710 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1385
timestamp 1712078602
transform 1 0 64262 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1397
timestamp 1712078602
transform 1 0 64814 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1401
timestamp 1712078602
transform 1 0 64998 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1413
timestamp 1712078602
transform 1 0 65550 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1425
timestamp 1712078602
transform 1 0 66102 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1429
timestamp 1712078602
transform 1 0 66286 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1441
timestamp 1712078602
transform 1 0 66838 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1453
timestamp 1712078602
transform 1 0 67390 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1457
timestamp 1712078602
transform 1 0 67574 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1469
timestamp 1712078602
transform 1 0 68126 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1481
timestamp 1712078602
transform 1 0 68678 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1485
timestamp 1712078602
transform 1 0 68862 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1497
timestamp 1712078602
transform 1 0 69414 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1509
timestamp 1712078602
transform 1 0 69966 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1513
timestamp 1712078602
transform 1 0 70150 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1525
timestamp 1712078602
transform 1 0 70702 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1537
timestamp 1712078602
transform 1 0 71254 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1541
timestamp 1712078602
transform 1 0 71438 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1553
timestamp 1712078602
transform 1 0 71990 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1565
timestamp 1712078602
transform 1 0 72542 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1569
timestamp 1712078602
transform 1 0 72726 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1581
timestamp 1712078602
transform 1 0 73278 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1593
timestamp 1712078602
transform 1 0 73830 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1597
timestamp 1712078602
transform 1 0 74014 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1609
timestamp 1712078602
transform 1 0 74566 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1621
timestamp 1712078602
transform 1 0 75118 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1625
timestamp 1712078602
transform 1 0 75302 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1637
timestamp 1712078602
transform 1 0 75854 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1649
timestamp 1712078602
transform 1 0 76406 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1653
timestamp 1712078602
transform 1 0 76590 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1665
timestamp 1712078602
transform 1 0 77142 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1677
timestamp 1712078602
transform 1 0 77694 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1681
timestamp 1712078602
transform 1 0 77878 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1693
timestamp 1712078602
transform 1 0 78430 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1705
timestamp 1712078602
transform 1 0 78982 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1709
timestamp 1712078602
transform 1 0 79166 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1721
timestamp 1712078602
transform 1 0 79718 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1733
timestamp 1712078602
transform 1 0 80270 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1737
timestamp 1712078602
transform 1 0 80454 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1749
timestamp 1712078602
transform 1 0 81006 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1761
timestamp 1712078602
transform 1 0 81558 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1765
timestamp 1712078602
transform 1 0 81742 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1777
timestamp 1712078602
transform 1 0 82294 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1789
timestamp 1712078602
transform 1 0 82846 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1793
timestamp 1712078602
transform 1 0 83030 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1805
timestamp 1712078602
transform 1 0 83582 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1817
timestamp 1712078602
transform 1 0 84134 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1821
timestamp 1712078602
transform 1 0 84318 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1833
timestamp 1712078602
transform 1 0 84870 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1845
timestamp 1712078602
transform 1 0 85422 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1849
timestamp 1712078602
transform 1 0 85606 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1861
timestamp 1712078602
transform 1 0 86158 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1873
timestamp 1712078602
transform 1 0 86710 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1877
timestamp 1712078602
transform 1 0 86894 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1889
timestamp 1712078602
transform 1 0 87446 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1901
timestamp 1712078602
transform 1 0 87998 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1905
timestamp 1712078602
transform 1 0 88182 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1917
timestamp 1712078602
transform 1 0 88734 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1929
timestamp 1712078602
transform 1 0 89286 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1933
timestamp 1712078602
transform 1 0 89470 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1945
timestamp 1712078602
transform 1 0 90022 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1957
timestamp 1712078602
transform 1 0 90574 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1961
timestamp 1712078602
transform 1 0 90758 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1973
timestamp 1712078602
transform 1 0 91310 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_1985
timestamp 1712078602
transform 1 0 91862 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_1989
timestamp 1712078602
transform 1 0 92046 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2001
timestamp 1712078602
transform 1 0 92598 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2013
timestamp 1712078602
transform 1 0 93150 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2017
timestamp 1712078602
transform 1 0 93334 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2029
timestamp 1712078602
transform 1 0 93886 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2041
timestamp 1712078602
transform 1 0 94438 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2045
timestamp 1712078602
transform 1 0 94622 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2057
timestamp 1712078602
transform 1 0 95174 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2069
timestamp 1712078602
transform 1 0 95726 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2073
timestamp 1712078602
transform 1 0 95910 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2085
timestamp 1712078602
transform 1 0 96462 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2097
timestamp 1712078602
transform 1 0 97014 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2101
timestamp 1712078602
transform 1 0 97198 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2113
timestamp 1712078602
transform 1 0 97750 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2125
timestamp 1712078602
transform 1 0 98302 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2129
timestamp 1712078602
transform 1 0 98486 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2141
timestamp 1712078602
transform 1 0 99038 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2153
timestamp 1712078602
transform 1 0 99590 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2157
timestamp 1712078602
transform 1 0 99774 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2169
timestamp 1712078602
transform 1 0 100326 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2181
timestamp 1712078602
transform 1 0 100878 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2185
timestamp 1712078602
transform 1 0 101062 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2197
timestamp 1712078602
transform 1 0 101614 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2209
timestamp 1712078602
transform 1 0 102166 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2213
timestamp 1712078602
transform 1 0 102350 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2225
timestamp 1712078602
transform 1 0 102902 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2237
timestamp 1712078602
transform 1 0 103454 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2241
timestamp 1712078602
transform 1 0 103638 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2253
timestamp 1712078602
transform 1 0 104190 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2265
timestamp 1712078602
transform 1 0 104742 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2269
timestamp 1712078602
transform 1 0 104926 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2281
timestamp 1712078602
transform 1 0 105478 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2293
timestamp 1712078602
transform 1 0 106030 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2297
timestamp 1712078602
transform 1 0 106214 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2309
timestamp 1712078602
transform 1 0 106766 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2321
timestamp 1712078602
transform 1 0 107318 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2325
timestamp 1712078602
transform 1 0 107502 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2337
timestamp 1712078602
transform 1 0 108054 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2349
timestamp 1712078602
transform 1 0 108606 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2353
timestamp 1712078602
transform 1 0 108790 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2365
timestamp 1712078602
transform 1 0 109342 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2377
timestamp 1712078602
transform 1 0 109894 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2381
timestamp 1712078602
transform 1 0 110078 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2393
timestamp 1712078602
transform 1 0 110630 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2405
timestamp 1712078602
transform 1 0 111182 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2409
timestamp 1712078602
transform 1 0 111366 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2421
timestamp 1712078602
transform 1 0 111918 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2433
timestamp 1712078602
transform 1 0 112470 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2437
timestamp 1712078602
transform 1 0 112654 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2449
timestamp 1712078602
transform 1 0 113206 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2461
timestamp 1712078602
transform 1 0 113758 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2465
timestamp 1712078602
transform 1 0 113942 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2477
timestamp 1712078602
transform 1 0 114494 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2489
timestamp 1712078602
transform 1 0 115046 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2493
timestamp 1712078602
transform 1 0 115230 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2505
timestamp 1712078602
transform 1 0 115782 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2517
timestamp 1712078602
transform 1 0 116334 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2521
timestamp 1712078602
transform 1 0 116518 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2533
timestamp 1712078602
transform 1 0 117070 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2545
timestamp 1712078602
transform 1 0 117622 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2549
timestamp 1712078602
transform 1 0 117806 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2561
timestamp 1712078602
transform 1 0 118358 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2573
timestamp 1712078602
transform 1 0 118910 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2577
timestamp 1712078602
transform 1 0 119094 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2589
timestamp 1712078602
transform 1 0 119646 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2601
timestamp 1712078602
transform 1 0 120198 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2605
timestamp 1712078602
transform 1 0 120382 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2617
timestamp 1712078602
transform 1 0 120934 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2629
timestamp 1712078602
transform 1 0 121486 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2633
timestamp 1712078602
transform 1 0 121670 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2645
timestamp 1712078602
transform 1 0 122222 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2657
timestamp 1712078602
transform 1 0 122774 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2661
timestamp 1712078602
transform 1 0 122958 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2673
timestamp 1712078602
transform 1 0 123510 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2685
timestamp 1712078602
transform 1 0 124062 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2689
timestamp 1712078602
transform 1 0 124246 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2701
timestamp 1712078602
transform 1 0 124798 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2713
timestamp 1712078602
transform 1 0 125350 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2717
timestamp 1712078602
transform 1 0 125534 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2729
timestamp 1712078602
transform 1 0 126086 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2741
timestamp 1712078602
transform 1 0 126638 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2745
timestamp 1712078602
transform 1 0 126822 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2757
timestamp 1712078602
transform 1 0 127374 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2769
timestamp 1712078602
transform 1 0 127926 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2773
timestamp 1712078602
transform 1 0 128110 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2785
timestamp 1712078602
transform 1 0 128662 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2797
timestamp 1712078602
transform 1 0 129214 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2801
timestamp 1712078602
transform 1 0 129398 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2813
timestamp 1712078602
transform 1 0 129950 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2825
timestamp 1712078602
transform 1 0 130502 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2829
timestamp 1712078602
transform 1 0 130686 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2841
timestamp 1712078602
transform 1 0 131238 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2853
timestamp 1712078602
transform 1 0 131790 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2857
timestamp 1712078602
transform 1 0 131974 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2869
timestamp 1712078602
transform 1 0 132526 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2881
timestamp 1712078602
transform 1 0 133078 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2885
timestamp 1712078602
transform 1 0 133262 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2897
timestamp 1712078602
transform 1 0 133814 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2909
timestamp 1712078602
transform 1 0 134366 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2913
timestamp 1712078602
transform 1 0 134550 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2925
timestamp 1712078602
transform 1 0 135102 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2937
timestamp 1712078602
transform 1 0 135654 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2941
timestamp 1712078602
transform 1 0 135838 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2953
timestamp 1712078602
transform 1 0 136390 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2965
timestamp 1712078602
transform 1 0 136942 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2969
timestamp 1712078602
transform 1 0 137126 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2981
timestamp 1712078602
transform 1 0 137678 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_2993
timestamp 1712078602
transform 1 0 138230 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_2997
timestamp 1712078602
transform 1 0 138414 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3009
timestamp 1712078602
transform 1 0 138966 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3021
timestamp 1712078602
transform 1 0 139518 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3025
timestamp 1712078602
transform 1 0 139702 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3037
timestamp 1712078602
transform 1 0 140254 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3049
timestamp 1712078602
transform 1 0 140806 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3053
timestamp 1712078602
transform 1 0 140990 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3065
timestamp 1712078602
transform 1 0 141542 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3077
timestamp 1712078602
transform 1 0 142094 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3081
timestamp 1712078602
transform 1 0 142278 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3093
timestamp 1712078602
transform 1 0 142830 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3105
timestamp 1712078602
transform 1 0 143382 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3109
timestamp 1712078602
transform 1 0 143566 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3121
timestamp 1712078602
transform 1 0 144118 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3133
timestamp 1712078602
transform 1 0 144670 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3137
timestamp 1712078602
transform 1 0 144854 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3149
timestamp 1712078602
transform 1 0 145406 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3161
timestamp 1712078602
transform 1 0 145958 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3165
timestamp 1712078602
transform 1 0 146142 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3177
timestamp 1712078602
transform 1 0 146694 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3189
timestamp 1712078602
transform 1 0 147246 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3193
timestamp 1712078602
transform 1 0 147430 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3205
timestamp 1712078602
transform 1 0 147982 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3217
timestamp 1712078602
transform 1 0 148534 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3221
timestamp 1712078602
transform 1 0 148718 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3233
timestamp 1712078602
transform 1 0 149270 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3245
timestamp 1712078602
transform 1 0 149822 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3249
timestamp 1712078602
transform 1 0 150006 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3261
timestamp 1712078602
transform 1 0 150558 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3273
timestamp 1712078602
transform 1 0 151110 0 1 1088
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3277
timestamp 1712078602
transform 1 0 151294 0 1 1088
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_0_3289
timestamp 1712078602
transform 1 0 151846 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_3301
timestamp 1712078602
transform 1 0 152398 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_0_3305 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 152582 0 1 1088
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1712078602
transform 1 0 690 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1712078602
transform 1 0 1242 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1712078602
transform 1 0 1794 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1712078602
transform 1 0 2346 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1712078602
transform 1 0 2898 0 -1 1632
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1712078602
transform 1 0 3082 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1712078602
transform 1 0 3174 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1712078602
transform 1 0 3726 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1712078602
transform 1 0 4278 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1712078602
transform 1 0 4830 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 5382 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1712078602
transform 1 0 5658 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1712078602
transform 1 0 5750 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1712078602
transform 1 0 6302 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1712078602
transform 1 0 6854 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1712078602
transform 1 0 7406 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1712078602
transform 1 0 7958 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1712078602
transform 1 0 8234 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1712078602
transform 1 0 8326 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1712078602
transform 1 0 8878 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1712078602
transform 1 0 9430 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1712078602
transform 1 0 9982 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1712078602
transform 1 0 10534 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1712078602
transform 1 0 10810 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1712078602
transform 1 0 10902 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1712078602
transform 1 0 11454 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1712078602
transform 1 0 12006 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1712078602
transform 1 0 12558 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1712078602
transform 1 0 13110 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1712078602
transform 1 0 13386 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1712078602
transform 1 0 13478 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1712078602
transform 1 0 14030 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1712078602
transform 1 0 14582 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1712078602
transform 1 0 15134 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1712078602
transform 1 0 15686 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1712078602
transform 1 0 15962 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1712078602
transform 1 0 16054 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1712078602
transform 1 0 16606 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1712078602
transform 1 0 17158 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1712078602
transform 1 0 17710 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1712078602
transform 1 0 18262 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1712078602
transform 1 0 18538 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1712078602
transform 1 0 18630 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1712078602
transform 1 0 19182 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1712078602
transform 1 0 19734 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1712078602
transform 1 0 20286 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1712078602
transform 1 0 20838 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1712078602
transform 1 0 21114 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1712078602
transform 1 0 21206 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1712078602
transform 1 0 21758 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1712078602
transform 1 0 22310 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1712078602
transform 1 0 22862 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1712078602
transform 1 0 23414 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1712078602
transform 1 0 23690 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1712078602
transform 1 0 23782 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1712078602
transform 1 0 24334 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1712078602
transform 1 0 24886 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1712078602
transform 1 0 25438 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1712078602
transform 1 0 25990 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1712078602
transform 1 0 26266 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1712078602
transform 1 0 26358 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1712078602
transform 1 0 26910 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1712078602
transform 1 0 27462 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1712078602
transform 1 0 28014 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1712078602
transform 1 0 28566 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1712078602
transform 1 0 28842 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1712078602
transform 1 0 28934 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1712078602
transform 1 0 29486 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1712078602
transform 1 0 30038 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1712078602
transform 1 0 30590 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1712078602
transform 1 0 31142 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1712078602
transform 1 0 31418 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1712078602
transform 1 0 31510 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1712078602
transform 1 0 32062 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1712078602
transform 1 0 32614 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1712078602
transform 1 0 33166 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1712078602
transform 1 0 33718 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1712078602
transform 1 0 33994 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1712078602
transform 1 0 34086 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1712078602
transform 1 0 34638 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1712078602
transform 1 0 35190 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1712078602
transform 1 0 35742 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1712078602
transform 1 0 36294 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1712078602
transform 1 0 36570 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1712078602
transform 1 0 36662 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1712078602
transform 1 0 37214 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1712078602
transform 1 0 37766 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1712078602
transform 1 0 38318 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1712078602
transform 1 0 38870 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1712078602
transform 1 0 39146 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1712078602
transform 1 0 39238 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1712078602
transform 1 0 39790 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1712078602
transform 1 0 40342 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1712078602
transform 1 0 40894 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1712078602
transform 1 0 41446 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1712078602
transform 1 0 41722 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1712078602
transform 1 0 41814 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1712078602
transform 1 0 42366 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1712078602
transform 1 0 42918 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1712078602
transform 1 0 43470 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1712078602
transform 1 0 44022 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1712078602
transform 1 0 44298 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1712078602
transform 1 0 44390 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1712078602
transform 1 0 44942 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1712078602
transform 1 0 45494 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1712078602
transform 1 0 46046 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1712078602
transform 1 0 46598 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1712078602
transform 1 0 46874 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1712078602
transform 1 0 46966 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1712078602
transform 1 0 47518 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1712078602
transform 1 0 48070 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1712078602
transform 1 0 48622 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1712078602
transform 1 0 49174 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1712078602
transform 1 0 49450 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1712078602
transform 1 0 49542 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1712078602
transform 1 0 50094 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1712078602
transform 1 0 50646 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1712078602
transform 1 0 51198 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1712078602
transform 1 0 51750 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1712078602
transform 1 0 52026 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1712078602
transform 1 0 52118 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1712078602
transform 1 0 52670 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1712078602
transform 1 0 53222 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1712078602
transform 1 0 53774 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1712078602
transform 1 0 54326 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1712078602
transform 1 0 54602 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1712078602
transform 1 0 54694 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1189
timestamp 1712078602
transform 1 0 55246 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1201
timestamp 1712078602
transform 1 0 55798 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1213
timestamp 1712078602
transform 1 0 56350 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1225
timestamp 1712078602
transform 1 0 56902 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1712078602
transform 1 0 57178 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1712078602
transform 1 0 57270 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1245
timestamp 1712078602
transform 1 0 57822 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1257
timestamp 1712078602
transform 1 0 58374 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1269
timestamp 1712078602
transform 1 0 58926 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1281
timestamp 1712078602
transform 1 0 59478 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1287
timestamp 1712078602
transform 1 0 59754 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1289
timestamp 1712078602
transform 1 0 59846 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1301
timestamp 1712078602
transform 1 0 60398 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1313
timestamp 1712078602
transform 1 0 60950 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1325
timestamp 1712078602
transform 1 0 61502 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1337
timestamp 1712078602
transform 1 0 62054 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1343
timestamp 1712078602
transform 1 0 62330 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1345
timestamp 1712078602
transform 1 0 62422 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1357
timestamp 1712078602
transform 1 0 62974 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1369
timestamp 1712078602
transform 1 0 63526 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1381
timestamp 1712078602
transform 1 0 64078 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1393
timestamp 1712078602
transform 1 0 64630 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1712078602
transform 1 0 64906 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1401
timestamp 1712078602
transform 1 0 64998 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1413
timestamp 1712078602
transform 1 0 65550 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1425
timestamp 1712078602
transform 1 0 66102 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1437
timestamp 1712078602
transform 1 0 66654 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1449
timestamp 1712078602
transform 1 0 67206 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1712078602
transform 1 0 67482 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1712078602
transform 1 0 67574 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1469
timestamp 1712078602
transform 1 0 68126 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1481
timestamp 1712078602
transform 1 0 68678 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1493
timestamp 1712078602
transform 1 0 69230 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1505
timestamp 1712078602
transform 1 0 69782 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1511
timestamp 1712078602
transform 1 0 70058 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1513
timestamp 1712078602
transform 1 0 70150 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1525
timestamp 1712078602
transform 1 0 70702 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1537
timestamp 1712078602
transform 1 0 71254 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1549
timestamp 1712078602
transform 1 0 71806 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1561
timestamp 1712078602
transform 1 0 72358 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1567
timestamp 1712078602
transform 1 0 72634 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1569
timestamp 1712078602
transform 1 0 72726 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1581
timestamp 1712078602
transform 1 0 73278 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1593
timestamp 1712078602
transform 1 0 73830 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1605
timestamp 1712078602
transform 1 0 74382 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1617
timestamp 1712078602
transform 1 0 74934 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1623
timestamp 1712078602
transform 1 0 75210 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1625
timestamp 1712078602
transform 1 0 75302 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1637
timestamp 1712078602
transform 1 0 75854 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1649
timestamp 1712078602
transform 1 0 76406 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1661
timestamp 1712078602
transform 1 0 76958 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1673
timestamp 1712078602
transform 1 0 77510 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1679
timestamp 1712078602
transform 1 0 77786 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1681
timestamp 1712078602
transform 1 0 77878 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1693
timestamp 1712078602
transform 1 0 78430 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1705
timestamp 1712078602
transform 1 0 78982 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1717
timestamp 1712078602
transform 1 0 79534 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1729
timestamp 1712078602
transform 1 0 80086 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1735
timestamp 1712078602
transform 1 0 80362 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1737
timestamp 1712078602
transform 1 0 80454 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1749
timestamp 1712078602
transform 1 0 81006 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1761
timestamp 1712078602
transform 1 0 81558 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1773
timestamp 1712078602
transform 1 0 82110 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1785
timestamp 1712078602
transform 1 0 82662 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1791
timestamp 1712078602
transform 1 0 82938 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1793
timestamp 1712078602
transform 1 0 83030 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1805
timestamp 1712078602
transform 1 0 83582 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1817
timestamp 1712078602
transform 1 0 84134 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1829
timestamp 1712078602
transform 1 0 84686 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1841
timestamp 1712078602
transform 1 0 85238 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1847
timestamp 1712078602
transform 1 0 85514 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1849
timestamp 1712078602
transform 1 0 85606 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1861
timestamp 1712078602
transform 1 0 86158 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1873
timestamp 1712078602
transform 1 0 86710 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1885
timestamp 1712078602
transform 1 0 87262 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1897
timestamp 1712078602
transform 1 0 87814 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1903
timestamp 1712078602
transform 1 0 88090 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1905
timestamp 1712078602
transform 1 0 88182 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1917
timestamp 1712078602
transform 1 0 88734 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1929
timestamp 1712078602
transform 1 0 89286 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1941
timestamp 1712078602
transform 1 0 89838 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_1953
timestamp 1712078602
transform 1 0 90390 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_1959
timestamp 1712078602
transform 1 0 90666 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1961
timestamp 1712078602
transform 1 0 90758 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1973
timestamp 1712078602
transform 1 0 91310 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1985
timestamp 1712078602
transform 1 0 91862 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_1997
timestamp 1712078602
transform 1 0 92414 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2009
timestamp 1712078602
transform 1 0 92966 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2015
timestamp 1712078602
transform 1 0 93242 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2017
timestamp 1712078602
transform 1 0 93334 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2029
timestamp 1712078602
transform 1 0 93886 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2041
timestamp 1712078602
transform 1 0 94438 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2053
timestamp 1712078602
transform 1 0 94990 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2065
timestamp 1712078602
transform 1 0 95542 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2071
timestamp 1712078602
transform 1 0 95818 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2073
timestamp 1712078602
transform 1 0 95910 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2085
timestamp 1712078602
transform 1 0 96462 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2097
timestamp 1712078602
transform 1 0 97014 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2109
timestamp 1712078602
transform 1 0 97566 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2121
timestamp 1712078602
transform 1 0 98118 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2127
timestamp 1712078602
transform 1 0 98394 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2129
timestamp 1712078602
transform 1 0 98486 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2141
timestamp 1712078602
transform 1 0 99038 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2153
timestamp 1712078602
transform 1 0 99590 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2165
timestamp 1712078602
transform 1 0 100142 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2177
timestamp 1712078602
transform 1 0 100694 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2183
timestamp 1712078602
transform 1 0 100970 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2185
timestamp 1712078602
transform 1 0 101062 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2197
timestamp 1712078602
transform 1 0 101614 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2209
timestamp 1712078602
transform 1 0 102166 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2221
timestamp 1712078602
transform 1 0 102718 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2233
timestamp 1712078602
transform 1 0 103270 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2239
timestamp 1712078602
transform 1 0 103546 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2241
timestamp 1712078602
transform 1 0 103638 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2253
timestamp 1712078602
transform 1 0 104190 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2265
timestamp 1712078602
transform 1 0 104742 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2277
timestamp 1712078602
transform 1 0 105294 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2289
timestamp 1712078602
transform 1 0 105846 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2295
timestamp 1712078602
transform 1 0 106122 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2297
timestamp 1712078602
transform 1 0 106214 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2309
timestamp 1712078602
transform 1 0 106766 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2321
timestamp 1712078602
transform 1 0 107318 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2333
timestamp 1712078602
transform 1 0 107870 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2345
timestamp 1712078602
transform 1 0 108422 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2351
timestamp 1712078602
transform 1 0 108698 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2353
timestamp 1712078602
transform 1 0 108790 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2365
timestamp 1712078602
transform 1 0 109342 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2377
timestamp 1712078602
transform 1 0 109894 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2389
timestamp 1712078602
transform 1 0 110446 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2401
timestamp 1712078602
transform 1 0 110998 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2407
timestamp 1712078602
transform 1 0 111274 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2409
timestamp 1712078602
transform 1 0 111366 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2421
timestamp 1712078602
transform 1 0 111918 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2433
timestamp 1712078602
transform 1 0 112470 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2445
timestamp 1712078602
transform 1 0 113022 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2457
timestamp 1712078602
transform 1 0 113574 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2463
timestamp 1712078602
transform 1 0 113850 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2465
timestamp 1712078602
transform 1 0 113942 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2477
timestamp 1712078602
transform 1 0 114494 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2489
timestamp 1712078602
transform 1 0 115046 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2501
timestamp 1712078602
transform 1 0 115598 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2513
timestamp 1712078602
transform 1 0 116150 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2519
timestamp 1712078602
transform 1 0 116426 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2521
timestamp 1712078602
transform 1 0 116518 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2533
timestamp 1712078602
transform 1 0 117070 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2545
timestamp 1712078602
transform 1 0 117622 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2557
timestamp 1712078602
transform 1 0 118174 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2569
timestamp 1712078602
transform 1 0 118726 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2575
timestamp 1712078602
transform 1 0 119002 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2577
timestamp 1712078602
transform 1 0 119094 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2589
timestamp 1712078602
transform 1 0 119646 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2601
timestamp 1712078602
transform 1 0 120198 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2613
timestamp 1712078602
transform 1 0 120750 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2625
timestamp 1712078602
transform 1 0 121302 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2631
timestamp 1712078602
transform 1 0 121578 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2633
timestamp 1712078602
transform 1 0 121670 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2645
timestamp 1712078602
transform 1 0 122222 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2657
timestamp 1712078602
transform 1 0 122774 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2669
timestamp 1712078602
transform 1 0 123326 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2681
timestamp 1712078602
transform 1 0 123878 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2687
timestamp 1712078602
transform 1 0 124154 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2689
timestamp 1712078602
transform 1 0 124246 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2701
timestamp 1712078602
transform 1 0 124798 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2713
timestamp 1712078602
transform 1 0 125350 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2725
timestamp 1712078602
transform 1 0 125902 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2737
timestamp 1712078602
transform 1 0 126454 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2743
timestamp 1712078602
transform 1 0 126730 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2745
timestamp 1712078602
transform 1 0 126822 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2757
timestamp 1712078602
transform 1 0 127374 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2769
timestamp 1712078602
transform 1 0 127926 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2781
timestamp 1712078602
transform 1 0 128478 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2793
timestamp 1712078602
transform 1 0 129030 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2799
timestamp 1712078602
transform 1 0 129306 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2801
timestamp 1712078602
transform 1 0 129398 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2813
timestamp 1712078602
transform 1 0 129950 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2825
timestamp 1712078602
transform 1 0 130502 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2837
timestamp 1712078602
transform 1 0 131054 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2849
timestamp 1712078602
transform 1 0 131606 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2855
timestamp 1712078602
transform 1 0 131882 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2857
timestamp 1712078602
transform 1 0 131974 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2869
timestamp 1712078602
transform 1 0 132526 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2881
timestamp 1712078602
transform 1 0 133078 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2893
timestamp 1712078602
transform 1 0 133630 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2905
timestamp 1712078602
transform 1 0 134182 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2911
timestamp 1712078602
transform 1 0 134458 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2913
timestamp 1712078602
transform 1 0 134550 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2925
timestamp 1712078602
transform 1 0 135102 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2937
timestamp 1712078602
transform 1 0 135654 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2949
timestamp 1712078602
transform 1 0 136206 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_2961
timestamp 1712078602
transform 1 0 136758 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_2967
timestamp 1712078602
transform 1 0 137034 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2969
timestamp 1712078602
transform 1 0 137126 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2981
timestamp 1712078602
transform 1 0 137678 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_2993
timestamp 1712078602
transform 1 0 138230 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3005
timestamp 1712078602
transform 1 0 138782 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_3017
timestamp 1712078602
transform 1 0 139334 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_3023
timestamp 1712078602
transform 1 0 139610 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3025
timestamp 1712078602
transform 1 0 139702 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3037
timestamp 1712078602
transform 1 0 140254 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3049
timestamp 1712078602
transform 1 0 140806 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3061
timestamp 1712078602
transform 1 0 141358 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_3073
timestamp 1712078602
transform 1 0 141910 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_3079
timestamp 1712078602
transform 1 0 142186 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3081
timestamp 1712078602
transform 1 0 142278 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3093
timestamp 1712078602
transform 1 0 142830 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3105
timestamp 1712078602
transform 1 0 143382 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3117
timestamp 1712078602
transform 1 0 143934 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_3129
timestamp 1712078602
transform 1 0 144486 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_3135
timestamp 1712078602
transform 1 0 144762 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3137
timestamp 1712078602
transform 1 0 144854 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3149
timestamp 1712078602
transform 1 0 145406 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3161
timestamp 1712078602
transform 1 0 145958 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3173
timestamp 1712078602
transform 1 0 146510 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_3185
timestamp 1712078602
transform 1 0 147062 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_3191
timestamp 1712078602
transform 1 0 147338 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3193
timestamp 1712078602
transform 1 0 147430 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3205
timestamp 1712078602
transform 1 0 147982 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3217
timestamp 1712078602
transform 1 0 148534 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3229
timestamp 1712078602
transform 1 0 149086 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_3241
timestamp 1712078602
transform 1 0 149638 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_3247
timestamp 1712078602
transform 1 0 149914 0 -1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3249
timestamp 1712078602
transform 1 0 150006 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3261
timestamp 1712078602
transform 1 0 150558 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3273
timestamp 1712078602
transform 1 0 151110 0 -1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_1_3285
timestamp 1712078602
transform 1 0 151662 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_3297
timestamp 1712078602
transform 1 0 152214 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_3303
timestamp 1712078602
transform 1 0 152490 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_1_3305
timestamp 1712078602
transform 1 0 152582 0 -1 1632
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1712078602
transform 1 0 690 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1712078602
transform 1 0 1242 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1712078602
transform 1 0 1794 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1712078602
transform 1 0 1886 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1712078602
transform 1 0 2438 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1712078602
transform 1 0 2990 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1712078602
transform 1 0 3542 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1712078602
transform 1 0 4094 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1712078602
transform 1 0 4370 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1712078602
transform 1 0 4462 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1712078602
transform 1 0 5014 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1712078602
transform 1 0 5566 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1712078602
transform 1 0 6118 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1712078602
transform 1 0 6670 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1712078602
transform 1 0 6946 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1712078602
transform 1 0 7038 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1712078602
transform 1 0 7590 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1712078602
transform 1 0 8142 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1712078602
transform 1 0 8694 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1712078602
transform 1 0 9246 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1712078602
transform 1 0 9522 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1712078602
transform 1 0 9614 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1712078602
transform 1 0 10166 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1712078602
transform 1 0 10718 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1712078602
transform 1 0 11270 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1712078602
transform 1 0 11822 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1712078602
transform 1 0 12098 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1712078602
transform 1 0 12190 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1712078602
transform 1 0 12742 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1712078602
transform 1 0 13294 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1712078602
transform 1 0 13846 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1712078602
transform 1 0 14398 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1712078602
transform 1 0 14674 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1712078602
transform 1 0 14766 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1712078602
transform 1 0 15318 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1712078602
transform 1 0 15870 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1712078602
transform 1 0 16422 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1712078602
transform 1 0 16974 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1712078602
transform 1 0 17250 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1712078602
transform 1 0 17342 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1712078602
transform 1 0 17894 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1712078602
transform 1 0 18446 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1712078602
transform 1 0 18998 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1712078602
transform 1 0 19550 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1712078602
transform 1 0 19826 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1712078602
transform 1 0 19918 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1712078602
transform 1 0 20470 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1712078602
transform 1 0 21022 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1712078602
transform 1 0 21574 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1712078602
transform 1 0 22126 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1712078602
transform 1 0 22402 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1712078602
transform 1 0 22494 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1712078602
transform 1 0 23046 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1712078602
transform 1 0 23598 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1712078602
transform 1 0 24150 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1712078602
transform 1 0 24702 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1712078602
transform 1 0 24978 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1712078602
transform 1 0 25070 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1712078602
transform 1 0 25622 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1712078602
transform 1 0 26174 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1712078602
transform 1 0 26726 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1712078602
transform 1 0 27278 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1712078602
transform 1 0 27554 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1712078602
transform 1 0 27646 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1712078602
transform 1 0 28198 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1712078602
transform 1 0 28750 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1712078602
transform 1 0 29302 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1712078602
transform 1 0 29854 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1712078602
transform 1 0 30130 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1712078602
transform 1 0 30222 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1712078602
transform 1 0 30774 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1712078602
transform 1 0 31326 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1712078602
transform 1 0 31878 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1712078602
transform 1 0 32430 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1712078602
transform 1 0 32706 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1712078602
transform 1 0 32798 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1712078602
transform 1 0 33350 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1712078602
transform 1 0 33902 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1712078602
transform 1 0 34454 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1712078602
transform 1 0 35006 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1712078602
transform 1 0 35282 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1712078602
transform 1 0 35374 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1712078602
transform 1 0 35926 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1712078602
transform 1 0 36478 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1712078602
transform 1 0 37030 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1712078602
transform 1 0 37582 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1712078602
transform 1 0 37858 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1712078602
transform 1 0 37950 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1712078602
transform 1 0 38502 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1712078602
transform 1 0 39054 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1712078602
transform 1 0 39606 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1712078602
transform 1 0 40158 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1712078602
transform 1 0 40434 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1712078602
transform 1 0 40526 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1712078602
transform 1 0 41078 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1712078602
transform 1 0 41630 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1712078602
transform 1 0 42182 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1712078602
transform 1 0 42734 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1712078602
transform 1 0 43010 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1712078602
transform 1 0 43102 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1712078602
transform 1 0 43654 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1712078602
transform 1 0 44206 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1712078602
transform 1 0 44758 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1712078602
transform 1 0 45310 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1712078602
transform 1 0 45586 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1712078602
transform 1 0 45678 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1712078602
transform 1 0 46230 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1712078602
transform 1 0 46782 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1712078602
transform 1 0 47334 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1712078602
transform 1 0 47886 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1712078602
transform 1 0 48162 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1712078602
transform 1 0 48254 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1712078602
transform 1 0 48806 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1712078602
transform 1 0 49358 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1712078602
transform 1 0 49910 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1712078602
transform 1 0 50462 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1712078602
transform 1 0 50738 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1712078602
transform 1 0 50830 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1712078602
transform 1 0 51382 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1712078602
transform 1 0 51934 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1712078602
transform 1 0 52486 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1712078602
transform 1 0 53038 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1712078602
transform 1 0 53314 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1712078602
transform 1 0 53406 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1712078602
transform 1 0 53958 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1712078602
transform 1 0 54510 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1712078602
transform 1 0 55062 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1712078602
transform 1 0 55614 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1712078602
transform 1 0 55890 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1712078602
transform 1 0 55982 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1712078602
transform 1 0 56534 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1712078602
transform 1 0 57086 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1712078602
transform 1 0 57638 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1253
timestamp 1712078602
transform 1 0 58190 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1712078602
transform 1 0 58466 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1261
timestamp 1712078602
transform 1 0 58558 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1273
timestamp 1712078602
transform 1 0 59110 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1285
timestamp 1712078602
transform 1 0 59662 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1297
timestamp 1712078602
transform 1 0 60214 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1309
timestamp 1712078602
transform 1 0 60766 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1315
timestamp 1712078602
transform 1 0 61042 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1317
timestamp 1712078602
transform 1 0 61134 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1329
timestamp 1712078602
transform 1 0 61686 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1341
timestamp 1712078602
transform 1 0 62238 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1353
timestamp 1712078602
transform 1 0 62790 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1365
timestamp 1712078602
transform 1 0 63342 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1712078602
transform 1 0 63618 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1373
timestamp 1712078602
transform 1 0 63710 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1385
timestamp 1712078602
transform 1 0 64262 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1397
timestamp 1712078602
transform 1 0 64814 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1409
timestamp 1712078602
transform 1 0 65366 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1421
timestamp 1712078602
transform 1 0 65918 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1712078602
transform 1 0 66194 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1429
timestamp 1712078602
transform 1 0 66286 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1441
timestamp 1712078602
transform 1 0 66838 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1453
timestamp 1712078602
transform 1 0 67390 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1465
timestamp 1712078602
transform 1 0 67942 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1477
timestamp 1712078602
transform 1 0 68494 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1483
timestamp 1712078602
transform 1 0 68770 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1712078602
transform 1 0 68862 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1712078602
transform 1 0 69414 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1712078602
transform 1 0 69966 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1712078602
transform 1 0 70518 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1712078602
transform 1 0 71070 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1712078602
transform 1 0 71346 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1712078602
transform 1 0 71438 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1712078602
transform 1 0 71990 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1712078602
transform 1 0 72542 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1712078602
transform 1 0 73094 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1712078602
transform 1 0 73646 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1712078602
transform 1 0 73922 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1597
timestamp 1712078602
transform 1 0 74014 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1609
timestamp 1712078602
transform 1 0 74566 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1621
timestamp 1712078602
transform 1 0 75118 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1633
timestamp 1712078602
transform 1 0 75670 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1645
timestamp 1712078602
transform 1 0 76222 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1651
timestamp 1712078602
transform 1 0 76498 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1653
timestamp 1712078602
transform 1 0 76590 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1665
timestamp 1712078602
transform 1 0 77142 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1677
timestamp 1712078602
transform 1 0 77694 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1689
timestamp 1712078602
transform 1 0 78246 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1701
timestamp 1712078602
transform 1 0 78798 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1707
timestamp 1712078602
transform 1 0 79074 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1709
timestamp 1712078602
transform 1 0 79166 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1721
timestamp 1712078602
transform 1 0 79718 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1733
timestamp 1712078602
transform 1 0 80270 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1745
timestamp 1712078602
transform 1 0 80822 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1757
timestamp 1712078602
transform 1 0 81374 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1763
timestamp 1712078602
transform 1 0 81650 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1765
timestamp 1712078602
transform 1 0 81742 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1777
timestamp 1712078602
transform 1 0 82294 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1789
timestamp 1712078602
transform 1 0 82846 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1801
timestamp 1712078602
transform 1 0 83398 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1813
timestamp 1712078602
transform 1 0 83950 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1819
timestamp 1712078602
transform 1 0 84226 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1821
timestamp 1712078602
transform 1 0 84318 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1833
timestamp 1712078602
transform 1 0 84870 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1845
timestamp 1712078602
transform 1 0 85422 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1857
timestamp 1712078602
transform 1 0 85974 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1869
timestamp 1712078602
transform 1 0 86526 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1875
timestamp 1712078602
transform 1 0 86802 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1877
timestamp 1712078602
transform 1 0 86894 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1889
timestamp 1712078602
transform 1 0 87446 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1901
timestamp 1712078602
transform 1 0 87998 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1913
timestamp 1712078602
transform 1 0 88550 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1925
timestamp 1712078602
transform 1 0 89102 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1931
timestamp 1712078602
transform 1 0 89378 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1933
timestamp 1712078602
transform 1 0 89470 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1945
timestamp 1712078602
transform 1 0 90022 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1957
timestamp 1712078602
transform 1 0 90574 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1969
timestamp 1712078602
transform 1 0 91126 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_1981
timestamp 1712078602
transform 1 0 91678 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_1987
timestamp 1712078602
transform 1 0 91954 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_1989
timestamp 1712078602
transform 1 0 92046 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2001
timestamp 1712078602
transform 1 0 92598 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2013
timestamp 1712078602
transform 1 0 93150 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2025
timestamp 1712078602
transform 1 0 93702 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2037
timestamp 1712078602
transform 1 0 94254 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2043
timestamp 1712078602
transform 1 0 94530 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2045
timestamp 1712078602
transform 1 0 94622 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2057
timestamp 1712078602
transform 1 0 95174 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2069
timestamp 1712078602
transform 1 0 95726 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2081
timestamp 1712078602
transform 1 0 96278 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2093
timestamp 1712078602
transform 1 0 96830 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2099
timestamp 1712078602
transform 1 0 97106 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2101
timestamp 1712078602
transform 1 0 97198 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2113
timestamp 1712078602
transform 1 0 97750 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2125
timestamp 1712078602
transform 1 0 98302 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2137
timestamp 1712078602
transform 1 0 98854 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2149
timestamp 1712078602
transform 1 0 99406 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2155
timestamp 1712078602
transform 1 0 99682 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2157
timestamp 1712078602
transform 1 0 99774 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2169
timestamp 1712078602
transform 1 0 100326 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2181
timestamp 1712078602
transform 1 0 100878 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2193
timestamp 1712078602
transform 1 0 101430 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2205
timestamp 1712078602
transform 1 0 101982 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2211
timestamp 1712078602
transform 1 0 102258 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2213
timestamp 1712078602
transform 1 0 102350 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2225
timestamp 1712078602
transform 1 0 102902 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2237
timestamp 1712078602
transform 1 0 103454 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2249
timestamp 1712078602
transform 1 0 104006 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2261
timestamp 1712078602
transform 1 0 104558 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2267
timestamp 1712078602
transform 1 0 104834 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2269
timestamp 1712078602
transform 1 0 104926 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2281
timestamp 1712078602
transform 1 0 105478 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2293
timestamp 1712078602
transform 1 0 106030 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2305
timestamp 1712078602
transform 1 0 106582 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2317
timestamp 1712078602
transform 1 0 107134 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2323
timestamp 1712078602
transform 1 0 107410 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2325
timestamp 1712078602
transform 1 0 107502 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2337
timestamp 1712078602
transform 1 0 108054 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2349
timestamp 1712078602
transform 1 0 108606 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2361
timestamp 1712078602
transform 1 0 109158 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2373
timestamp 1712078602
transform 1 0 109710 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2379
timestamp 1712078602
transform 1 0 109986 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2381
timestamp 1712078602
transform 1 0 110078 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2393
timestamp 1712078602
transform 1 0 110630 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2405
timestamp 1712078602
transform 1 0 111182 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2417
timestamp 1712078602
transform 1 0 111734 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2429
timestamp 1712078602
transform 1 0 112286 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2435
timestamp 1712078602
transform 1 0 112562 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2437
timestamp 1712078602
transform 1 0 112654 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2449
timestamp 1712078602
transform 1 0 113206 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2461
timestamp 1712078602
transform 1 0 113758 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2473
timestamp 1712078602
transform 1 0 114310 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2485
timestamp 1712078602
transform 1 0 114862 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2491
timestamp 1712078602
transform 1 0 115138 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2493
timestamp 1712078602
transform 1 0 115230 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2505
timestamp 1712078602
transform 1 0 115782 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2517
timestamp 1712078602
transform 1 0 116334 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2529
timestamp 1712078602
transform 1 0 116886 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2541
timestamp 1712078602
transform 1 0 117438 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2547
timestamp 1712078602
transform 1 0 117714 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2549
timestamp 1712078602
transform 1 0 117806 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2561
timestamp 1712078602
transform 1 0 118358 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2573
timestamp 1712078602
transform 1 0 118910 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2585
timestamp 1712078602
transform 1 0 119462 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2597
timestamp 1712078602
transform 1 0 120014 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2603
timestamp 1712078602
transform 1 0 120290 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2605
timestamp 1712078602
transform 1 0 120382 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2617
timestamp 1712078602
transform 1 0 120934 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2629
timestamp 1712078602
transform 1 0 121486 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2641
timestamp 1712078602
transform 1 0 122038 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2653
timestamp 1712078602
transform 1 0 122590 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2659
timestamp 1712078602
transform 1 0 122866 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2661
timestamp 1712078602
transform 1 0 122958 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2673
timestamp 1712078602
transform 1 0 123510 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2685
timestamp 1712078602
transform 1 0 124062 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2697
timestamp 1712078602
transform 1 0 124614 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2709
timestamp 1712078602
transform 1 0 125166 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2715
timestamp 1712078602
transform 1 0 125442 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2717
timestamp 1712078602
transform 1 0 125534 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2729
timestamp 1712078602
transform 1 0 126086 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2741
timestamp 1712078602
transform 1 0 126638 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2753
timestamp 1712078602
transform 1 0 127190 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2765
timestamp 1712078602
transform 1 0 127742 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2771
timestamp 1712078602
transform 1 0 128018 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2773
timestamp 1712078602
transform 1 0 128110 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2785
timestamp 1712078602
transform 1 0 128662 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2797
timestamp 1712078602
transform 1 0 129214 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2809
timestamp 1712078602
transform 1 0 129766 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2821
timestamp 1712078602
transform 1 0 130318 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2827
timestamp 1712078602
transform 1 0 130594 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2829
timestamp 1712078602
transform 1 0 130686 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2841
timestamp 1712078602
transform 1 0 131238 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2853
timestamp 1712078602
transform 1 0 131790 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2865
timestamp 1712078602
transform 1 0 132342 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2877
timestamp 1712078602
transform 1 0 132894 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2883
timestamp 1712078602
transform 1 0 133170 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2885
timestamp 1712078602
transform 1 0 133262 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2897
timestamp 1712078602
transform 1 0 133814 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2909
timestamp 1712078602
transform 1 0 134366 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2921
timestamp 1712078602
transform 1 0 134918 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2933
timestamp 1712078602
transform 1 0 135470 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2939
timestamp 1712078602
transform 1 0 135746 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2941
timestamp 1712078602
transform 1 0 135838 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2953
timestamp 1712078602
transform 1 0 136390 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2965
timestamp 1712078602
transform 1 0 136942 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2977
timestamp 1712078602
transform 1 0 137494 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_2989
timestamp 1712078602
transform 1 0 138046 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_2995
timestamp 1712078602
transform 1 0 138322 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_2997
timestamp 1712078602
transform 1 0 138414 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3009
timestamp 1712078602
transform 1 0 138966 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3021
timestamp 1712078602
transform 1 0 139518 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3033
timestamp 1712078602
transform 1 0 140070 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_3045
timestamp 1712078602
transform 1 0 140622 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_3051
timestamp 1712078602
transform 1 0 140898 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3053
timestamp 1712078602
transform 1 0 140990 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3065
timestamp 1712078602
transform 1 0 141542 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3077
timestamp 1712078602
transform 1 0 142094 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3089
timestamp 1712078602
transform 1 0 142646 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_3101
timestamp 1712078602
transform 1 0 143198 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_3107
timestamp 1712078602
transform 1 0 143474 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3109
timestamp 1712078602
transform 1 0 143566 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3121
timestamp 1712078602
transform 1 0 144118 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3133
timestamp 1712078602
transform 1 0 144670 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3145
timestamp 1712078602
transform 1 0 145222 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_3157
timestamp 1712078602
transform 1 0 145774 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_3163
timestamp 1712078602
transform 1 0 146050 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3165
timestamp 1712078602
transform 1 0 146142 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3177
timestamp 1712078602
transform 1 0 146694 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3189
timestamp 1712078602
transform 1 0 147246 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3201
timestamp 1712078602
transform 1 0 147798 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_3213
timestamp 1712078602
transform 1 0 148350 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_3219
timestamp 1712078602
transform 1 0 148626 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3221
timestamp 1712078602
transform 1 0 148718 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3233
timestamp 1712078602
transform 1 0 149270 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3245
timestamp 1712078602
transform 1 0 149822 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3257
timestamp 1712078602
transform 1 0 150374 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_3269
timestamp 1712078602
transform 1 0 150926 0 1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_2_3275
timestamp 1712078602
transform 1 0 151202 0 1 1632
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3277
timestamp 1712078602
transform 1 0 151294 0 1 1632
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_2_3289
timestamp 1712078602
transform 1 0 151846 0 1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_2_3301 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 152398 0 1 1632
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1712078602
transform 1 0 690 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1712078602
transform 1 0 1242 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1712078602
transform 1 0 1794 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1712078602
transform 1 0 2346 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1712078602
transform 1 0 2898 0 -1 2176
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1712078602
transform 1 0 3082 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1712078602
transform 1 0 3174 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1712078602
transform 1 0 3726 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1712078602
transform 1 0 4278 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1712078602
transform 1 0 4830 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1712078602
transform 1 0 5382 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1712078602
transform 1 0 5658 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1712078602
transform 1 0 5750 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1712078602
transform 1 0 6302 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1712078602
transform 1 0 6854 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1712078602
transform 1 0 7406 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1712078602
transform 1 0 7958 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1712078602
transform 1 0 8234 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1712078602
transform 1 0 8326 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1712078602
transform 1 0 8878 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1712078602
transform 1 0 9430 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1712078602
transform 1 0 9982 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1712078602
transform 1 0 10534 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1712078602
transform 1 0 10810 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1712078602
transform 1 0 10902 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1712078602
transform 1 0 11454 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1712078602
transform 1 0 12006 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1712078602
transform 1 0 12558 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1712078602
transform 1 0 13110 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1712078602
transform 1 0 13386 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1712078602
transform 1 0 13478 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1712078602
transform 1 0 14030 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1712078602
transform 1 0 14582 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1712078602
transform 1 0 15134 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1712078602
transform 1 0 15686 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1712078602
transform 1 0 15962 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1712078602
transform 1 0 16054 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1712078602
transform 1 0 16606 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1712078602
transform 1 0 17158 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1712078602
transform 1 0 17710 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1712078602
transform 1 0 18262 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1712078602
transform 1 0 18538 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1712078602
transform 1 0 18630 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1712078602
transform 1 0 19182 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1712078602
transform 1 0 19734 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1712078602
transform 1 0 20286 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1712078602
transform 1 0 20838 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1712078602
transform 1 0 21114 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1712078602
transform 1 0 21206 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1712078602
transform 1 0 21758 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1712078602
transform 1 0 22310 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1712078602
transform 1 0 22862 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1712078602
transform 1 0 23414 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1712078602
transform 1 0 23690 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1712078602
transform 1 0 23782 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1712078602
transform 1 0 24334 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1712078602
transform 1 0 24886 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1712078602
transform 1 0 25438 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1712078602
transform 1 0 25990 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1712078602
transform 1 0 26266 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1712078602
transform 1 0 26358 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1712078602
transform 1 0 26910 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1712078602
transform 1 0 27462 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1712078602
transform 1 0 28014 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1712078602
transform 1 0 28566 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1712078602
transform 1 0 28842 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1712078602
transform 1 0 28934 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1712078602
transform 1 0 29486 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1712078602
transform 1 0 30038 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1712078602
transform 1 0 30590 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1712078602
transform 1 0 31142 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1712078602
transform 1 0 31418 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1712078602
transform 1 0 31510 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1712078602
transform 1 0 32062 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1712078602
transform 1 0 32614 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1712078602
transform 1 0 33166 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1712078602
transform 1 0 33718 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1712078602
transform 1 0 33994 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1712078602
transform 1 0 34086 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1712078602
transform 1 0 34638 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1712078602
transform 1 0 35190 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1712078602
transform 1 0 35742 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1712078602
transform 1 0 36294 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1712078602
transform 1 0 36570 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1712078602
transform 1 0 36662 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1712078602
transform 1 0 37214 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1712078602
transform 1 0 37766 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1712078602
transform 1 0 38318 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1712078602
transform 1 0 38870 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1712078602
transform 1 0 39146 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1712078602
transform 1 0 39238 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1712078602
transform 1 0 39790 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1712078602
transform 1 0 40342 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1712078602
transform 1 0 40894 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1712078602
transform 1 0 41446 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1712078602
transform 1 0 41722 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1712078602
transform 1 0 41814 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1712078602
transform 1 0 42366 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1712078602
transform 1 0 42918 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1712078602
transform 1 0 43470 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1712078602
transform 1 0 44022 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1712078602
transform 1 0 44298 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1712078602
transform 1 0 44390 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1712078602
transform 1 0 44942 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1712078602
transform 1 0 45494 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1712078602
transform 1 0 46046 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1712078602
transform 1 0 46598 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1712078602
transform 1 0 46874 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1712078602
transform 1 0 46966 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1712078602
transform 1 0 47518 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1712078602
transform 1 0 48070 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1712078602
transform 1 0 48622 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1712078602
transform 1 0 49174 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1712078602
transform 1 0 49450 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1712078602
transform 1 0 49542 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1712078602
transform 1 0 50094 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1712078602
transform 1 0 50646 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1712078602
transform 1 0 51198 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1712078602
transform 1 0 51750 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1712078602
transform 1 0 52026 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1712078602
transform 1 0 52118 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1712078602
transform 1 0 52670 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1712078602
transform 1 0 53222 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1712078602
transform 1 0 53774 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1712078602
transform 1 0 54326 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1712078602
transform 1 0 54602 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1712078602
transform 1 0 54694 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1712078602
transform 1 0 55246 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1712078602
transform 1 0 55798 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1712078602
transform 1 0 56350 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1712078602
transform 1 0 56902 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1712078602
transform 1 0 57178 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1712078602
transform 1 0 57270 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1712078602
transform 1 0 57822 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1712078602
transform 1 0 58374 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1269
timestamp 1712078602
transform 1 0 58926 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1281
timestamp 1712078602
transform 1 0 59478 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1287
timestamp 1712078602
transform 1 0 59754 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1289
timestamp 1712078602
transform 1 0 59846 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1301
timestamp 1712078602
transform 1 0 60398 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1313
timestamp 1712078602
transform 1 0 60950 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1325
timestamp 1712078602
transform 1 0 61502 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1337
timestamp 1712078602
transform 1 0 62054 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1343
timestamp 1712078602
transform 1 0 62330 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1345
timestamp 1712078602
transform 1 0 62422 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1357
timestamp 1712078602
transform 1 0 62974 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1369
timestamp 1712078602
transform 1 0 63526 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1381
timestamp 1712078602
transform 1 0 64078 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1393
timestamp 1712078602
transform 1 0 64630 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1712078602
transform 1 0 64906 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1712078602
transform 1 0 64998 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1712078602
transform 1 0 65550 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1712078602
transform 1 0 66102 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1712078602
transform 1 0 66654 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1712078602
transform 1 0 67206 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1712078602
transform 1 0 67482 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1712078602
transform 1 0 67574 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1712078602
transform 1 0 68126 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1481
timestamp 1712078602
transform 1 0 68678 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1493
timestamp 1712078602
transform 1 0 69230 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1505
timestamp 1712078602
transform 1 0 69782 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1712078602
transform 1 0 70058 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1513
timestamp 1712078602
transform 1 0 70150 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1525
timestamp 1712078602
transform 1 0 70702 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1537
timestamp 1712078602
transform 1 0 71254 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1549
timestamp 1712078602
transform 1 0 71806 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1561
timestamp 1712078602
transform 1 0 72358 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1567
timestamp 1712078602
transform 1 0 72634 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1569
timestamp 1712078602
transform 1 0 72726 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1581
timestamp 1712078602
transform 1 0 73278 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1593
timestamp 1712078602
transform 1 0 73830 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1605
timestamp 1712078602
transform 1 0 74382 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1617
timestamp 1712078602
transform 1 0 74934 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1712078602
transform 1 0 75210 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1625
timestamp 1712078602
transform 1 0 75302 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1637
timestamp 1712078602
transform 1 0 75854 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1649
timestamp 1712078602
transform 1 0 76406 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1661
timestamp 1712078602
transform 1 0 76958 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1673
timestamp 1712078602
transform 1 0 77510 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1679
timestamp 1712078602
transform 1 0 77786 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1681
timestamp 1712078602
transform 1 0 77878 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1693
timestamp 1712078602
transform 1 0 78430 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1705
timestamp 1712078602
transform 1 0 78982 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1717
timestamp 1712078602
transform 1 0 79534 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1729
timestamp 1712078602
transform 1 0 80086 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1735
timestamp 1712078602
transform 1 0 80362 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1737
timestamp 1712078602
transform 1 0 80454 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1749
timestamp 1712078602
transform 1 0 81006 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1761
timestamp 1712078602
transform 1 0 81558 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1773
timestamp 1712078602
transform 1 0 82110 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1785
timestamp 1712078602
transform 1 0 82662 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1791
timestamp 1712078602
transform 1 0 82938 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1793
timestamp 1712078602
transform 1 0 83030 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1805
timestamp 1712078602
transform 1 0 83582 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1817
timestamp 1712078602
transform 1 0 84134 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1829
timestamp 1712078602
transform 1 0 84686 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1841
timestamp 1712078602
transform 1 0 85238 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1847
timestamp 1712078602
transform 1 0 85514 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1849
timestamp 1712078602
transform 1 0 85606 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1861
timestamp 1712078602
transform 1 0 86158 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1873
timestamp 1712078602
transform 1 0 86710 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1885
timestamp 1712078602
transform 1 0 87262 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1897
timestamp 1712078602
transform 1 0 87814 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1903
timestamp 1712078602
transform 1 0 88090 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1905
timestamp 1712078602
transform 1 0 88182 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1917
timestamp 1712078602
transform 1 0 88734 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1929
timestamp 1712078602
transform 1 0 89286 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1941
timestamp 1712078602
transform 1 0 89838 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_1953
timestamp 1712078602
transform 1 0 90390 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_1959
timestamp 1712078602
transform 1 0 90666 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1961
timestamp 1712078602
transform 1 0 90758 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1973
timestamp 1712078602
transform 1 0 91310 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1985
timestamp 1712078602
transform 1 0 91862 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_1997
timestamp 1712078602
transform 1 0 92414 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2009
timestamp 1712078602
transform 1 0 92966 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2015
timestamp 1712078602
transform 1 0 93242 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2017
timestamp 1712078602
transform 1 0 93334 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2029
timestamp 1712078602
transform 1 0 93886 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2041
timestamp 1712078602
transform 1 0 94438 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2053
timestamp 1712078602
transform 1 0 94990 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2065
timestamp 1712078602
transform 1 0 95542 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2071
timestamp 1712078602
transform 1 0 95818 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2073
timestamp 1712078602
transform 1 0 95910 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2085
timestamp 1712078602
transform 1 0 96462 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2097
timestamp 1712078602
transform 1 0 97014 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2109
timestamp 1712078602
transform 1 0 97566 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2121
timestamp 1712078602
transform 1 0 98118 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2127
timestamp 1712078602
transform 1 0 98394 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2129
timestamp 1712078602
transform 1 0 98486 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2141
timestamp 1712078602
transform 1 0 99038 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2153
timestamp 1712078602
transform 1 0 99590 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2165
timestamp 1712078602
transform 1 0 100142 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2177
timestamp 1712078602
transform 1 0 100694 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2183
timestamp 1712078602
transform 1 0 100970 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2185
timestamp 1712078602
transform 1 0 101062 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2197
timestamp 1712078602
transform 1 0 101614 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2209
timestamp 1712078602
transform 1 0 102166 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2221
timestamp 1712078602
transform 1 0 102718 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2233
timestamp 1712078602
transform 1 0 103270 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2239
timestamp 1712078602
transform 1 0 103546 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2241
timestamp 1712078602
transform 1 0 103638 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2253
timestamp 1712078602
transform 1 0 104190 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2265
timestamp 1712078602
transform 1 0 104742 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2277
timestamp 1712078602
transform 1 0 105294 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2289
timestamp 1712078602
transform 1 0 105846 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2295
timestamp 1712078602
transform 1 0 106122 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2297
timestamp 1712078602
transform 1 0 106214 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2309
timestamp 1712078602
transform 1 0 106766 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2321
timestamp 1712078602
transform 1 0 107318 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2333
timestamp 1712078602
transform 1 0 107870 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2345
timestamp 1712078602
transform 1 0 108422 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2351
timestamp 1712078602
transform 1 0 108698 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2353
timestamp 1712078602
transform 1 0 108790 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2365
timestamp 1712078602
transform 1 0 109342 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2377
timestamp 1712078602
transform 1 0 109894 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2389
timestamp 1712078602
transform 1 0 110446 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2401
timestamp 1712078602
transform 1 0 110998 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2407
timestamp 1712078602
transform 1 0 111274 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2409
timestamp 1712078602
transform 1 0 111366 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2421
timestamp 1712078602
transform 1 0 111918 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2433
timestamp 1712078602
transform 1 0 112470 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2445
timestamp 1712078602
transform 1 0 113022 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2457
timestamp 1712078602
transform 1 0 113574 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2463
timestamp 1712078602
transform 1 0 113850 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2465
timestamp 1712078602
transform 1 0 113942 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2477
timestamp 1712078602
transform 1 0 114494 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2489
timestamp 1712078602
transform 1 0 115046 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2501
timestamp 1712078602
transform 1 0 115598 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2513
timestamp 1712078602
transform 1 0 116150 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2519
timestamp 1712078602
transform 1 0 116426 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2521
timestamp 1712078602
transform 1 0 116518 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2533
timestamp 1712078602
transform 1 0 117070 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2545
timestamp 1712078602
transform 1 0 117622 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2557
timestamp 1712078602
transform 1 0 118174 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2569
timestamp 1712078602
transform 1 0 118726 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2575
timestamp 1712078602
transform 1 0 119002 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2577
timestamp 1712078602
transform 1 0 119094 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2589
timestamp 1712078602
transform 1 0 119646 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2601
timestamp 1712078602
transform 1 0 120198 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2613
timestamp 1712078602
transform 1 0 120750 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2625
timestamp 1712078602
transform 1 0 121302 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2631
timestamp 1712078602
transform 1 0 121578 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2633
timestamp 1712078602
transform 1 0 121670 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2645
timestamp 1712078602
transform 1 0 122222 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2657
timestamp 1712078602
transform 1 0 122774 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2669
timestamp 1712078602
transform 1 0 123326 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2681
timestamp 1712078602
transform 1 0 123878 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2687
timestamp 1712078602
transform 1 0 124154 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2689
timestamp 1712078602
transform 1 0 124246 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2701
timestamp 1712078602
transform 1 0 124798 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2713
timestamp 1712078602
transform 1 0 125350 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2725
timestamp 1712078602
transform 1 0 125902 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2737
timestamp 1712078602
transform 1 0 126454 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2743
timestamp 1712078602
transform 1 0 126730 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2745
timestamp 1712078602
transform 1 0 126822 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2757
timestamp 1712078602
transform 1 0 127374 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2769
timestamp 1712078602
transform 1 0 127926 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2781
timestamp 1712078602
transform 1 0 128478 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2793
timestamp 1712078602
transform 1 0 129030 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2799
timestamp 1712078602
transform 1 0 129306 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2801
timestamp 1712078602
transform 1 0 129398 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2813
timestamp 1712078602
transform 1 0 129950 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2825
timestamp 1712078602
transform 1 0 130502 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2837
timestamp 1712078602
transform 1 0 131054 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2849
timestamp 1712078602
transform 1 0 131606 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2855
timestamp 1712078602
transform 1 0 131882 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2857
timestamp 1712078602
transform 1 0 131974 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2869
timestamp 1712078602
transform 1 0 132526 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2881
timestamp 1712078602
transform 1 0 133078 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2893
timestamp 1712078602
transform 1 0 133630 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2905
timestamp 1712078602
transform 1 0 134182 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2911
timestamp 1712078602
transform 1 0 134458 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2913
timestamp 1712078602
transform 1 0 134550 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2925
timestamp 1712078602
transform 1 0 135102 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2937
timestamp 1712078602
transform 1 0 135654 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2949
timestamp 1712078602
transform 1 0 136206 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_2961
timestamp 1712078602
transform 1 0 136758 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_2967
timestamp 1712078602
transform 1 0 137034 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2969
timestamp 1712078602
transform 1 0 137126 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2981
timestamp 1712078602
transform 1 0 137678 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_2993
timestamp 1712078602
transform 1 0 138230 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3005
timestamp 1712078602
transform 1 0 138782 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_3017
timestamp 1712078602
transform 1 0 139334 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_3023
timestamp 1712078602
transform 1 0 139610 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3025
timestamp 1712078602
transform 1 0 139702 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3037
timestamp 1712078602
transform 1 0 140254 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3049
timestamp 1712078602
transform 1 0 140806 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3061
timestamp 1712078602
transform 1 0 141358 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_3073
timestamp 1712078602
transform 1 0 141910 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_3079
timestamp 1712078602
transform 1 0 142186 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3081
timestamp 1712078602
transform 1 0 142278 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3093
timestamp 1712078602
transform 1 0 142830 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3105
timestamp 1712078602
transform 1 0 143382 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3117
timestamp 1712078602
transform 1 0 143934 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_3129
timestamp 1712078602
transform 1 0 144486 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_3135
timestamp 1712078602
transform 1 0 144762 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3137
timestamp 1712078602
transform 1 0 144854 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3149
timestamp 1712078602
transform 1 0 145406 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3161
timestamp 1712078602
transform 1 0 145958 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3173
timestamp 1712078602
transform 1 0 146510 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_3185
timestamp 1712078602
transform 1 0 147062 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_3191
timestamp 1712078602
transform 1 0 147338 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3193
timestamp 1712078602
transform 1 0 147430 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3205
timestamp 1712078602
transform 1 0 147982 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3217
timestamp 1712078602
transform 1 0 148534 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3229
timestamp 1712078602
transform 1 0 149086 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_3241
timestamp 1712078602
transform 1 0 149638 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_3247
timestamp 1712078602
transform 1 0 149914 0 -1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3249
timestamp 1712078602
transform 1 0 150006 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3261
timestamp 1712078602
transform 1 0 150558 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3273
timestamp 1712078602
transform 1 0 151110 0 -1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_3_3285
timestamp 1712078602
transform 1 0 151662 0 -1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_3_3297
timestamp 1712078602
transform 1 0 152214 0 -1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_3_3303
timestamp 1712078602
transform 1 0 152490 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_3_3305
timestamp 1712078602
transform 1 0 152582 0 -1 2176
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1712078602
transform 1 0 690 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1712078602
transform 1 0 1242 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1712078602
transform 1 0 1794 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1712078602
transform 1 0 1886 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1712078602
transform 1 0 2438 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1712078602
transform 1 0 2990 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1712078602
transform 1 0 3542 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1712078602
transform 1 0 4094 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1712078602
transform 1 0 4370 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1712078602
transform 1 0 4462 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1712078602
transform 1 0 5014 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1712078602
transform 1 0 5566 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1712078602
transform 1 0 6118 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1712078602
transform 1 0 6670 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1712078602
transform 1 0 6946 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1712078602
transform 1 0 7038 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1712078602
transform 1 0 7590 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1712078602
transform 1 0 8142 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1712078602
transform 1 0 8694 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1712078602
transform 1 0 9246 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1712078602
transform 1 0 9522 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1712078602
transform 1 0 9614 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1712078602
transform 1 0 10166 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1712078602
transform 1 0 10718 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1712078602
transform 1 0 11270 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1712078602
transform 1 0 11822 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1712078602
transform 1 0 12098 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1712078602
transform 1 0 12190 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1712078602
transform 1 0 12742 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1712078602
transform 1 0 13294 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1712078602
transform 1 0 13846 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1712078602
transform 1 0 14398 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1712078602
transform 1 0 14674 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1712078602
transform 1 0 14766 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1712078602
transform 1 0 15318 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1712078602
transform 1 0 15870 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1712078602
transform 1 0 16422 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1712078602
transform 1 0 16974 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1712078602
transform 1 0 17250 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1712078602
transform 1 0 17342 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1712078602
transform 1 0 17894 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1712078602
transform 1 0 18446 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1712078602
transform 1 0 18998 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1712078602
transform 1 0 19550 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1712078602
transform 1 0 19826 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1712078602
transform 1 0 19918 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1712078602
transform 1 0 20470 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1712078602
transform 1 0 21022 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1712078602
transform 1 0 21574 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1712078602
transform 1 0 22126 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1712078602
transform 1 0 22402 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1712078602
transform 1 0 22494 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1712078602
transform 1 0 23046 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1712078602
transform 1 0 23598 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1712078602
transform 1 0 24150 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1712078602
transform 1 0 24702 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1712078602
transform 1 0 24978 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1712078602
transform 1 0 25070 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1712078602
transform 1 0 25622 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1712078602
transform 1 0 26174 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1712078602
transform 1 0 26726 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1712078602
transform 1 0 27278 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1712078602
transform 1 0 27554 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1712078602
transform 1 0 27646 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1712078602
transform 1 0 28198 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1712078602
transform 1 0 28750 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1712078602
transform 1 0 29302 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1712078602
transform 1 0 29854 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1712078602
transform 1 0 30130 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1712078602
transform 1 0 30222 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1712078602
transform 1 0 30774 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1712078602
transform 1 0 31326 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1712078602
transform 1 0 31878 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1712078602
transform 1 0 32430 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1712078602
transform 1 0 32706 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1712078602
transform 1 0 32798 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1712078602
transform 1 0 33350 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1712078602
transform 1 0 33902 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1712078602
transform 1 0 34454 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1712078602
transform 1 0 35006 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1712078602
transform 1 0 35282 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1712078602
transform 1 0 35374 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1712078602
transform 1 0 35926 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1712078602
transform 1 0 36478 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1712078602
transform 1 0 37030 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1712078602
transform 1 0 37582 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1712078602
transform 1 0 37858 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1712078602
transform 1 0 37950 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1712078602
transform 1 0 38502 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1712078602
transform 1 0 39054 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1712078602
transform 1 0 39606 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1712078602
transform 1 0 40158 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1712078602
transform 1 0 40434 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1712078602
transform 1 0 40526 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1712078602
transform 1 0 41078 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1712078602
transform 1 0 41630 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1712078602
transform 1 0 42182 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1712078602
transform 1 0 42734 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1712078602
transform 1 0 43010 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1712078602
transform 1 0 43102 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1712078602
transform 1 0 43654 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1712078602
transform 1 0 44206 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1712078602
transform 1 0 44758 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1712078602
transform 1 0 45310 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1712078602
transform 1 0 45586 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1712078602
transform 1 0 45678 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1712078602
transform 1 0 46230 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1712078602
transform 1 0 46782 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1712078602
transform 1 0 47334 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1712078602
transform 1 0 47886 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1712078602
transform 1 0 48162 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1712078602
transform 1 0 48254 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1712078602
transform 1 0 48806 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1712078602
transform 1 0 49358 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1712078602
transform 1 0 49910 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1712078602
transform 1 0 50462 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1712078602
transform 1 0 50738 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1712078602
transform 1 0 50830 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1712078602
transform 1 0 51382 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1712078602
transform 1 0 51934 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1712078602
transform 1 0 52486 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1712078602
transform 1 0 53038 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1712078602
transform 1 0 53314 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1712078602
transform 1 0 53406 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1712078602
transform 1 0 53958 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1712078602
transform 1 0 54510 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1712078602
transform 1 0 55062 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1712078602
transform 1 0 55614 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1712078602
transform 1 0 55890 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1712078602
transform 1 0 55982 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1712078602
transform 1 0 56534 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1712078602
transform 1 0 57086 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1712078602
transform 1 0 57638 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1712078602
transform 1 0 58190 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1712078602
transform 1 0 58466 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1712078602
transform 1 0 58558 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1273
timestamp 1712078602
transform 1 0 59110 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1285
timestamp 1712078602
transform 1 0 59662 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1297
timestamp 1712078602
transform 1 0 60214 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1309
timestamp 1712078602
transform 1 0 60766 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1315
timestamp 1712078602
transform 1 0 61042 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1317
timestamp 1712078602
transform 1 0 61134 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1329
timestamp 1712078602
transform 1 0 61686 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1341
timestamp 1712078602
transform 1 0 62238 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1353
timestamp 1712078602
transform 1 0 62790 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1365
timestamp 1712078602
transform 1 0 63342 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1371
timestamp 1712078602
transform 1 0 63618 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1373
timestamp 1712078602
transform 1 0 63710 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1385
timestamp 1712078602
transform 1 0 64262 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1397
timestamp 1712078602
transform 1 0 64814 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1409
timestamp 1712078602
transform 1 0 65366 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1421
timestamp 1712078602
transform 1 0 65918 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1427
timestamp 1712078602
transform 1 0 66194 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1712078602
transform 1 0 66286 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1441
timestamp 1712078602
transform 1 0 66838 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1453
timestamp 1712078602
transform 1 0 67390 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1465
timestamp 1712078602
transform 1 0 67942 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1477
timestamp 1712078602
transform 1 0 68494 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1483
timestamp 1712078602
transform 1 0 68770 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1485
timestamp 1712078602
transform 1 0 68862 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1497
timestamp 1712078602
transform 1 0 69414 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1509
timestamp 1712078602
transform 1 0 69966 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1521
timestamp 1712078602
transform 1 0 70518 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1533
timestamp 1712078602
transform 1 0 71070 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1539
timestamp 1712078602
transform 1 0 71346 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1712078602
transform 1 0 71438 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1712078602
transform 1 0 71990 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1565
timestamp 1712078602
transform 1 0 72542 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1577
timestamp 1712078602
transform 1 0 73094 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1589
timestamp 1712078602
transform 1 0 73646 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1712078602
transform 1 0 73922 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1597
timestamp 1712078602
transform 1 0 74014 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1609
timestamp 1712078602
transform 1 0 74566 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1621
timestamp 1712078602
transform 1 0 75118 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1633
timestamp 1712078602
transform 1 0 75670 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1645
timestamp 1712078602
transform 1 0 76222 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1651
timestamp 1712078602
transform 1 0 76498 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1653
timestamp 1712078602
transform 1 0 76590 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1665
timestamp 1712078602
transform 1 0 77142 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1677
timestamp 1712078602
transform 1 0 77694 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1689
timestamp 1712078602
transform 1 0 78246 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1701
timestamp 1712078602
transform 1 0 78798 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1707
timestamp 1712078602
transform 1 0 79074 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1709
timestamp 1712078602
transform 1 0 79166 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1721
timestamp 1712078602
transform 1 0 79718 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1733
timestamp 1712078602
transform 1 0 80270 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1745
timestamp 1712078602
transform 1 0 80822 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1757
timestamp 1712078602
transform 1 0 81374 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1763
timestamp 1712078602
transform 1 0 81650 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1765
timestamp 1712078602
transform 1 0 81742 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1777
timestamp 1712078602
transform 1 0 82294 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1789
timestamp 1712078602
transform 1 0 82846 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1801
timestamp 1712078602
transform 1 0 83398 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1813
timestamp 1712078602
transform 1 0 83950 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1819
timestamp 1712078602
transform 1 0 84226 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1821
timestamp 1712078602
transform 1 0 84318 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1833
timestamp 1712078602
transform 1 0 84870 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1845
timestamp 1712078602
transform 1 0 85422 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1857
timestamp 1712078602
transform 1 0 85974 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1869
timestamp 1712078602
transform 1 0 86526 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1875
timestamp 1712078602
transform 1 0 86802 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1877
timestamp 1712078602
transform 1 0 86894 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1889
timestamp 1712078602
transform 1 0 87446 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1901
timestamp 1712078602
transform 1 0 87998 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1913
timestamp 1712078602
transform 1 0 88550 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1925
timestamp 1712078602
transform 1 0 89102 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1931
timestamp 1712078602
transform 1 0 89378 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1933
timestamp 1712078602
transform 1 0 89470 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1945
timestamp 1712078602
transform 1 0 90022 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1957
timestamp 1712078602
transform 1 0 90574 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1969
timestamp 1712078602
transform 1 0 91126 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_1981
timestamp 1712078602
transform 1 0 91678 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_1987
timestamp 1712078602
transform 1 0 91954 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_1989
timestamp 1712078602
transform 1 0 92046 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2001
timestamp 1712078602
transform 1 0 92598 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2013
timestamp 1712078602
transform 1 0 93150 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2025
timestamp 1712078602
transform 1 0 93702 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2037
timestamp 1712078602
transform 1 0 94254 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2043
timestamp 1712078602
transform 1 0 94530 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2045
timestamp 1712078602
transform 1 0 94622 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2057
timestamp 1712078602
transform 1 0 95174 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2069
timestamp 1712078602
transform 1 0 95726 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2081
timestamp 1712078602
transform 1 0 96278 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2093
timestamp 1712078602
transform 1 0 96830 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2099
timestamp 1712078602
transform 1 0 97106 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2101
timestamp 1712078602
transform 1 0 97198 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2113
timestamp 1712078602
transform 1 0 97750 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2125
timestamp 1712078602
transform 1 0 98302 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2137
timestamp 1712078602
transform 1 0 98854 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2149
timestamp 1712078602
transform 1 0 99406 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2155
timestamp 1712078602
transform 1 0 99682 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2157
timestamp 1712078602
transform 1 0 99774 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2169
timestamp 1712078602
transform 1 0 100326 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2181
timestamp 1712078602
transform 1 0 100878 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2193
timestamp 1712078602
transform 1 0 101430 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2205
timestamp 1712078602
transform 1 0 101982 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2211
timestamp 1712078602
transform 1 0 102258 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2213
timestamp 1712078602
transform 1 0 102350 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2225
timestamp 1712078602
transform 1 0 102902 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2237
timestamp 1712078602
transform 1 0 103454 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2249
timestamp 1712078602
transform 1 0 104006 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2261
timestamp 1712078602
transform 1 0 104558 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2267
timestamp 1712078602
transform 1 0 104834 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2269
timestamp 1712078602
transform 1 0 104926 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2281
timestamp 1712078602
transform 1 0 105478 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2293
timestamp 1712078602
transform 1 0 106030 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2305
timestamp 1712078602
transform 1 0 106582 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2317
timestamp 1712078602
transform 1 0 107134 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2323
timestamp 1712078602
transform 1 0 107410 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2325
timestamp 1712078602
transform 1 0 107502 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2337
timestamp 1712078602
transform 1 0 108054 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2349
timestamp 1712078602
transform 1 0 108606 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2361
timestamp 1712078602
transform 1 0 109158 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2373
timestamp 1712078602
transform 1 0 109710 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2379
timestamp 1712078602
transform 1 0 109986 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2381
timestamp 1712078602
transform 1 0 110078 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2393
timestamp 1712078602
transform 1 0 110630 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2405
timestamp 1712078602
transform 1 0 111182 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2417
timestamp 1712078602
transform 1 0 111734 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2429
timestamp 1712078602
transform 1 0 112286 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2435
timestamp 1712078602
transform 1 0 112562 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2437
timestamp 1712078602
transform 1 0 112654 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2449
timestamp 1712078602
transform 1 0 113206 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2461
timestamp 1712078602
transform 1 0 113758 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2473
timestamp 1712078602
transform 1 0 114310 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2485
timestamp 1712078602
transform 1 0 114862 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2491
timestamp 1712078602
transform 1 0 115138 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2493
timestamp 1712078602
transform 1 0 115230 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2505
timestamp 1712078602
transform 1 0 115782 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2517
timestamp 1712078602
transform 1 0 116334 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2529
timestamp 1712078602
transform 1 0 116886 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2541
timestamp 1712078602
transform 1 0 117438 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2547
timestamp 1712078602
transform 1 0 117714 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2549
timestamp 1712078602
transform 1 0 117806 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2561
timestamp 1712078602
transform 1 0 118358 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2573
timestamp 1712078602
transform 1 0 118910 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2585
timestamp 1712078602
transform 1 0 119462 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2597
timestamp 1712078602
transform 1 0 120014 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2603
timestamp 1712078602
transform 1 0 120290 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2605
timestamp 1712078602
transform 1 0 120382 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2617
timestamp 1712078602
transform 1 0 120934 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2629
timestamp 1712078602
transform 1 0 121486 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2641
timestamp 1712078602
transform 1 0 122038 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2653
timestamp 1712078602
transform 1 0 122590 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2659
timestamp 1712078602
transform 1 0 122866 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2661
timestamp 1712078602
transform 1 0 122958 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2673
timestamp 1712078602
transform 1 0 123510 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2685
timestamp 1712078602
transform 1 0 124062 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2697
timestamp 1712078602
transform 1 0 124614 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2709
timestamp 1712078602
transform 1 0 125166 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2715
timestamp 1712078602
transform 1 0 125442 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2717
timestamp 1712078602
transform 1 0 125534 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2729
timestamp 1712078602
transform 1 0 126086 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2741
timestamp 1712078602
transform 1 0 126638 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2753
timestamp 1712078602
transform 1 0 127190 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2765
timestamp 1712078602
transform 1 0 127742 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2771
timestamp 1712078602
transform 1 0 128018 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2773
timestamp 1712078602
transform 1 0 128110 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2785
timestamp 1712078602
transform 1 0 128662 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2797
timestamp 1712078602
transform 1 0 129214 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2809
timestamp 1712078602
transform 1 0 129766 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2821
timestamp 1712078602
transform 1 0 130318 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2827
timestamp 1712078602
transform 1 0 130594 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2829
timestamp 1712078602
transform 1 0 130686 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2841
timestamp 1712078602
transform 1 0 131238 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2853
timestamp 1712078602
transform 1 0 131790 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2865
timestamp 1712078602
transform 1 0 132342 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2877
timestamp 1712078602
transform 1 0 132894 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2883
timestamp 1712078602
transform 1 0 133170 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2885
timestamp 1712078602
transform 1 0 133262 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2897
timestamp 1712078602
transform 1 0 133814 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2909
timestamp 1712078602
transform 1 0 134366 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2921
timestamp 1712078602
transform 1 0 134918 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2933
timestamp 1712078602
transform 1 0 135470 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2939
timestamp 1712078602
transform 1 0 135746 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2941
timestamp 1712078602
transform 1 0 135838 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2953
timestamp 1712078602
transform 1 0 136390 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2965
timestamp 1712078602
transform 1 0 136942 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2977
timestamp 1712078602
transform 1 0 137494 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_2989
timestamp 1712078602
transform 1 0 138046 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_2995
timestamp 1712078602
transform 1 0 138322 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_2997
timestamp 1712078602
transform 1 0 138414 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3009
timestamp 1712078602
transform 1 0 138966 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3021
timestamp 1712078602
transform 1 0 139518 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3033
timestamp 1712078602
transform 1 0 140070 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_3045
timestamp 1712078602
transform 1 0 140622 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_3051
timestamp 1712078602
transform 1 0 140898 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3053
timestamp 1712078602
transform 1 0 140990 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3065
timestamp 1712078602
transform 1 0 141542 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3077
timestamp 1712078602
transform 1 0 142094 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3089
timestamp 1712078602
transform 1 0 142646 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_3101
timestamp 1712078602
transform 1 0 143198 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_3107
timestamp 1712078602
transform 1 0 143474 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3109
timestamp 1712078602
transform 1 0 143566 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3121
timestamp 1712078602
transform 1 0 144118 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3133
timestamp 1712078602
transform 1 0 144670 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3145
timestamp 1712078602
transform 1 0 145222 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_3157
timestamp 1712078602
transform 1 0 145774 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_3163
timestamp 1712078602
transform 1 0 146050 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3165
timestamp 1712078602
transform 1 0 146142 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3177
timestamp 1712078602
transform 1 0 146694 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3189
timestamp 1712078602
transform 1 0 147246 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3201
timestamp 1712078602
transform 1 0 147798 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_3213
timestamp 1712078602
transform 1 0 148350 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_3219
timestamp 1712078602
transform 1 0 148626 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3221
timestamp 1712078602
transform 1 0 148718 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3233
timestamp 1712078602
transform 1 0 149270 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3245
timestamp 1712078602
transform 1 0 149822 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3257
timestamp 1712078602
transform 1 0 150374 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_4_3269
timestamp 1712078602
transform 1 0 150926 0 1 2176
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_4_3275
timestamp 1712078602
transform 1 0 151202 0 1 2176
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3277
timestamp 1712078602
transform 1 0 151294 0 1 2176
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_4_3289
timestamp 1712078602
transform 1 0 151846 0 1 2176
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_4_3301
timestamp 1712078602
transform 1 0 152398 0 1 2176
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1712078602
transform 1 0 690 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1712078602
transform 1 0 1242 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1712078602
transform 1 0 1794 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1712078602
transform 1 0 2346 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1712078602
transform 1 0 2898 0 -1 2720
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1712078602
transform 1 0 3082 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1712078602
transform 1 0 3174 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1712078602
transform 1 0 3726 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1712078602
transform 1 0 4278 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1712078602
transform 1 0 4830 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1712078602
transform 1 0 5382 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1712078602
transform 1 0 5658 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1712078602
transform 1 0 5750 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1712078602
transform 1 0 6302 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1712078602
transform 1 0 6854 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1712078602
transform 1 0 7406 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1712078602
transform 1 0 7958 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1712078602
transform 1 0 8234 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1712078602
transform 1 0 8326 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1712078602
transform 1 0 8878 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1712078602
transform 1 0 9430 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1712078602
transform 1 0 9982 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1712078602
transform 1 0 10534 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1712078602
transform 1 0 10810 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1712078602
transform 1 0 10902 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1712078602
transform 1 0 11454 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1712078602
transform 1 0 12006 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1712078602
transform 1 0 12558 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1712078602
transform 1 0 13110 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1712078602
transform 1 0 13386 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1712078602
transform 1 0 13478 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1712078602
transform 1 0 14030 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1712078602
transform 1 0 14582 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1712078602
transform 1 0 15134 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1712078602
transform 1 0 15686 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1712078602
transform 1 0 15962 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1712078602
transform 1 0 16054 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1712078602
transform 1 0 16606 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1712078602
transform 1 0 17158 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1712078602
transform 1 0 17710 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1712078602
transform 1 0 18262 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1712078602
transform 1 0 18538 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1712078602
transform 1 0 18630 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1712078602
transform 1 0 19182 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1712078602
transform 1 0 19734 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1712078602
transform 1 0 20286 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1712078602
transform 1 0 20838 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1712078602
transform 1 0 21114 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1712078602
transform 1 0 21206 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1712078602
transform 1 0 21758 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1712078602
transform 1 0 22310 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1712078602
transform 1 0 22862 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1712078602
transform 1 0 23414 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1712078602
transform 1 0 23690 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1712078602
transform 1 0 23782 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1712078602
transform 1 0 24334 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1712078602
transform 1 0 24886 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1712078602
transform 1 0 25438 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1712078602
transform 1 0 25990 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1712078602
transform 1 0 26266 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1712078602
transform 1 0 26358 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1712078602
transform 1 0 26910 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1712078602
transform 1 0 27462 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1712078602
transform 1 0 28014 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1712078602
transform 1 0 28566 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1712078602
transform 1 0 28842 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1712078602
transform 1 0 28934 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1712078602
transform 1 0 29486 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1712078602
transform 1 0 30038 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1712078602
transform 1 0 30590 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1712078602
transform 1 0 31142 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1712078602
transform 1 0 31418 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1712078602
transform 1 0 31510 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1712078602
transform 1 0 32062 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1712078602
transform 1 0 32614 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1712078602
transform 1 0 33166 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1712078602
transform 1 0 33718 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1712078602
transform 1 0 33994 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1712078602
transform 1 0 34086 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1712078602
transform 1 0 34638 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1712078602
transform 1 0 35190 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1712078602
transform 1 0 35742 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1712078602
transform 1 0 36294 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1712078602
transform 1 0 36570 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1712078602
transform 1 0 36662 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1712078602
transform 1 0 37214 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1712078602
transform 1 0 37766 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1712078602
transform 1 0 38318 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1712078602
transform 1 0 38870 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1712078602
transform 1 0 39146 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1712078602
transform 1 0 39238 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1712078602
transform 1 0 39790 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1712078602
transform 1 0 40342 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1712078602
transform 1 0 40894 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1712078602
transform 1 0 41446 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1712078602
transform 1 0 41722 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1712078602
transform 1 0 41814 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1712078602
transform 1 0 42366 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1712078602
transform 1 0 42918 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1712078602
transform 1 0 43470 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1712078602
transform 1 0 44022 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1712078602
transform 1 0 44298 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1712078602
transform 1 0 44390 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1712078602
transform 1 0 44942 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1712078602
transform 1 0 45494 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1712078602
transform 1 0 46046 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1712078602
transform 1 0 46598 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1712078602
transform 1 0 46874 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1712078602
transform 1 0 46966 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1712078602
transform 1 0 47518 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1712078602
transform 1 0 48070 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1712078602
transform 1 0 48622 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1712078602
transform 1 0 49174 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1712078602
transform 1 0 49450 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1712078602
transform 1 0 49542 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1712078602
transform 1 0 50094 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1712078602
transform 1 0 50646 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1712078602
transform 1 0 51198 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1712078602
transform 1 0 51750 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1712078602
transform 1 0 52026 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1712078602
transform 1 0 52118 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1712078602
transform 1 0 52670 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1712078602
transform 1 0 53222 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1712078602
transform 1 0 53774 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1712078602
transform 1 0 54326 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1712078602
transform 1 0 54602 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1712078602
transform 1 0 54694 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1712078602
transform 1 0 55246 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1712078602
transform 1 0 55798 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1712078602
transform 1 0 56350 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1712078602
transform 1 0 56902 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1712078602
transform 1 0 57178 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1712078602
transform 1 0 57270 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1712078602
transform 1 0 57822 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1712078602
transform 1 0 58374 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1269
timestamp 1712078602
transform 1 0 58926 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1281
timestamp 1712078602
transform 1 0 59478 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1712078602
transform 1 0 59754 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1289
timestamp 1712078602
transform 1 0 59846 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1301
timestamp 1712078602
transform 1 0 60398 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1313
timestamp 1712078602
transform 1 0 60950 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1325
timestamp 1712078602
transform 1 0 61502 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1337
timestamp 1712078602
transform 1 0 62054 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1343
timestamp 1712078602
transform 1 0 62330 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1345
timestamp 1712078602
transform 1 0 62422 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1357
timestamp 1712078602
transform 1 0 62974 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1369
timestamp 1712078602
transform 1 0 63526 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1381
timestamp 1712078602
transform 1 0 64078 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1393
timestamp 1712078602
transform 1 0 64630 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1399
timestamp 1712078602
transform 1 0 64906 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1401
timestamp 1712078602
transform 1 0 64998 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1413
timestamp 1712078602
transform 1 0 65550 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1425
timestamp 1712078602
transform 1 0 66102 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1437
timestamp 1712078602
transform 1 0 66654 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1449
timestamp 1712078602
transform 1 0 67206 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1455
timestamp 1712078602
transform 1 0 67482 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1457
timestamp 1712078602
transform 1 0 67574 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1469
timestamp 1712078602
transform 1 0 68126 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1481
timestamp 1712078602
transform 1 0 68678 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1493
timestamp 1712078602
transform 1 0 69230 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1505
timestamp 1712078602
transform 1 0 69782 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1511
timestamp 1712078602
transform 1 0 70058 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1513
timestamp 1712078602
transform 1 0 70150 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1525
timestamp 1712078602
transform 1 0 70702 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1537
timestamp 1712078602
transform 1 0 71254 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1549
timestamp 1712078602
transform 1 0 71806 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1561
timestamp 1712078602
transform 1 0 72358 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1567
timestamp 1712078602
transform 1 0 72634 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1569
timestamp 1712078602
transform 1 0 72726 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1581
timestamp 1712078602
transform 1 0 73278 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1593
timestamp 1712078602
transform 1 0 73830 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1605
timestamp 1712078602
transform 1 0 74382 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1617
timestamp 1712078602
transform 1 0 74934 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1712078602
transform 1 0 75210 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1625
timestamp 1712078602
transform 1 0 75302 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1637
timestamp 1712078602
transform 1 0 75854 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1649
timestamp 1712078602
transform 1 0 76406 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1661
timestamp 1712078602
transform 1 0 76958 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1712078602
transform 1 0 77510 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1712078602
transform 1 0 77786 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1681
timestamp 1712078602
transform 1 0 77878 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1693
timestamp 1712078602
transform 1 0 78430 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1705
timestamp 1712078602
transform 1 0 78982 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1717
timestamp 1712078602
transform 1 0 79534 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1729
timestamp 1712078602
transform 1 0 80086 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1735
timestamp 1712078602
transform 1 0 80362 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1737
timestamp 1712078602
transform 1 0 80454 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1749
timestamp 1712078602
transform 1 0 81006 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1761
timestamp 1712078602
transform 1 0 81558 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1773
timestamp 1712078602
transform 1 0 82110 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1785
timestamp 1712078602
transform 1 0 82662 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1791
timestamp 1712078602
transform 1 0 82938 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1793
timestamp 1712078602
transform 1 0 83030 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1805
timestamp 1712078602
transform 1 0 83582 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1817
timestamp 1712078602
transform 1 0 84134 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1829
timestamp 1712078602
transform 1 0 84686 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1841
timestamp 1712078602
transform 1 0 85238 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1847
timestamp 1712078602
transform 1 0 85514 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1849
timestamp 1712078602
transform 1 0 85606 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1861
timestamp 1712078602
transform 1 0 86158 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1873
timestamp 1712078602
transform 1 0 86710 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1885
timestamp 1712078602
transform 1 0 87262 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1897
timestamp 1712078602
transform 1 0 87814 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1903
timestamp 1712078602
transform 1 0 88090 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1905
timestamp 1712078602
transform 1 0 88182 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1917
timestamp 1712078602
transform 1 0 88734 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1929
timestamp 1712078602
transform 1 0 89286 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1941
timestamp 1712078602
transform 1 0 89838 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_1953
timestamp 1712078602
transform 1 0 90390 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_1959
timestamp 1712078602
transform 1 0 90666 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1961
timestamp 1712078602
transform 1 0 90758 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1973
timestamp 1712078602
transform 1 0 91310 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1985
timestamp 1712078602
transform 1 0 91862 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_1997
timestamp 1712078602
transform 1 0 92414 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2009
timestamp 1712078602
transform 1 0 92966 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2015
timestamp 1712078602
transform 1 0 93242 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2017
timestamp 1712078602
transform 1 0 93334 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2029
timestamp 1712078602
transform 1 0 93886 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2041
timestamp 1712078602
transform 1 0 94438 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2053
timestamp 1712078602
transform 1 0 94990 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2065
timestamp 1712078602
transform 1 0 95542 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2071
timestamp 1712078602
transform 1 0 95818 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2073
timestamp 1712078602
transform 1 0 95910 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2085
timestamp 1712078602
transform 1 0 96462 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2097
timestamp 1712078602
transform 1 0 97014 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2109
timestamp 1712078602
transform 1 0 97566 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2121
timestamp 1712078602
transform 1 0 98118 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2127
timestamp 1712078602
transform 1 0 98394 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2129
timestamp 1712078602
transform 1 0 98486 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2141
timestamp 1712078602
transform 1 0 99038 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2153
timestamp 1712078602
transform 1 0 99590 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2165
timestamp 1712078602
transform 1 0 100142 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2177
timestamp 1712078602
transform 1 0 100694 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2183
timestamp 1712078602
transform 1 0 100970 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2185
timestamp 1712078602
transform 1 0 101062 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2197
timestamp 1712078602
transform 1 0 101614 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2209
timestamp 1712078602
transform 1 0 102166 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2221
timestamp 1712078602
transform 1 0 102718 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2233
timestamp 1712078602
transform 1 0 103270 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2239
timestamp 1712078602
transform 1 0 103546 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2241
timestamp 1712078602
transform 1 0 103638 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2253
timestamp 1712078602
transform 1 0 104190 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2265
timestamp 1712078602
transform 1 0 104742 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2277
timestamp 1712078602
transform 1 0 105294 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2289
timestamp 1712078602
transform 1 0 105846 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2295
timestamp 1712078602
transform 1 0 106122 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2297
timestamp 1712078602
transform 1 0 106214 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2309
timestamp 1712078602
transform 1 0 106766 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2321
timestamp 1712078602
transform 1 0 107318 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2333
timestamp 1712078602
transform 1 0 107870 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2345
timestamp 1712078602
transform 1 0 108422 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2351
timestamp 1712078602
transform 1 0 108698 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2353
timestamp 1712078602
transform 1 0 108790 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2365
timestamp 1712078602
transform 1 0 109342 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2377
timestamp 1712078602
transform 1 0 109894 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2389
timestamp 1712078602
transform 1 0 110446 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2401
timestamp 1712078602
transform 1 0 110998 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2407
timestamp 1712078602
transform 1 0 111274 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2409
timestamp 1712078602
transform 1 0 111366 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2421
timestamp 1712078602
transform 1 0 111918 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2433
timestamp 1712078602
transform 1 0 112470 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2445
timestamp 1712078602
transform 1 0 113022 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2457
timestamp 1712078602
transform 1 0 113574 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2463
timestamp 1712078602
transform 1 0 113850 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2465
timestamp 1712078602
transform 1 0 113942 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2477
timestamp 1712078602
transform 1 0 114494 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2489
timestamp 1712078602
transform 1 0 115046 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2501
timestamp 1712078602
transform 1 0 115598 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2513
timestamp 1712078602
transform 1 0 116150 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2519
timestamp 1712078602
transform 1 0 116426 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2521
timestamp 1712078602
transform 1 0 116518 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2533
timestamp 1712078602
transform 1 0 117070 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2545
timestamp 1712078602
transform 1 0 117622 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2557
timestamp 1712078602
transform 1 0 118174 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2569
timestamp 1712078602
transform 1 0 118726 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2575
timestamp 1712078602
transform 1 0 119002 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2577
timestamp 1712078602
transform 1 0 119094 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2589
timestamp 1712078602
transform 1 0 119646 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2601
timestamp 1712078602
transform 1 0 120198 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2613
timestamp 1712078602
transform 1 0 120750 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2625
timestamp 1712078602
transform 1 0 121302 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2631
timestamp 1712078602
transform 1 0 121578 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2633
timestamp 1712078602
transform 1 0 121670 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2645
timestamp 1712078602
transform 1 0 122222 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2657
timestamp 1712078602
transform 1 0 122774 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2669
timestamp 1712078602
transform 1 0 123326 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2681
timestamp 1712078602
transform 1 0 123878 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2687
timestamp 1712078602
transform 1 0 124154 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2689
timestamp 1712078602
transform 1 0 124246 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2701
timestamp 1712078602
transform 1 0 124798 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2713
timestamp 1712078602
transform 1 0 125350 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2725
timestamp 1712078602
transform 1 0 125902 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2737
timestamp 1712078602
transform 1 0 126454 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2743
timestamp 1712078602
transform 1 0 126730 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2745
timestamp 1712078602
transform 1 0 126822 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2757
timestamp 1712078602
transform 1 0 127374 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2769
timestamp 1712078602
transform 1 0 127926 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2781
timestamp 1712078602
transform 1 0 128478 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2793
timestamp 1712078602
transform 1 0 129030 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2799
timestamp 1712078602
transform 1 0 129306 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2801
timestamp 1712078602
transform 1 0 129398 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2813
timestamp 1712078602
transform 1 0 129950 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2825
timestamp 1712078602
transform 1 0 130502 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2837
timestamp 1712078602
transform 1 0 131054 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2849
timestamp 1712078602
transform 1 0 131606 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2855
timestamp 1712078602
transform 1 0 131882 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2857
timestamp 1712078602
transform 1 0 131974 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2869
timestamp 1712078602
transform 1 0 132526 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2881
timestamp 1712078602
transform 1 0 133078 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2893
timestamp 1712078602
transform 1 0 133630 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2905
timestamp 1712078602
transform 1 0 134182 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2911
timestamp 1712078602
transform 1 0 134458 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2913
timestamp 1712078602
transform 1 0 134550 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2925
timestamp 1712078602
transform 1 0 135102 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2937
timestamp 1712078602
transform 1 0 135654 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2949
timestamp 1712078602
transform 1 0 136206 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_2961
timestamp 1712078602
transform 1 0 136758 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_2967
timestamp 1712078602
transform 1 0 137034 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2969
timestamp 1712078602
transform 1 0 137126 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2981
timestamp 1712078602
transform 1 0 137678 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_2993
timestamp 1712078602
transform 1 0 138230 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3005
timestamp 1712078602
transform 1 0 138782 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_3017
timestamp 1712078602
transform 1 0 139334 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_3023
timestamp 1712078602
transform 1 0 139610 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3025
timestamp 1712078602
transform 1 0 139702 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3037
timestamp 1712078602
transform 1 0 140254 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3049
timestamp 1712078602
transform 1 0 140806 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3061
timestamp 1712078602
transform 1 0 141358 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_3073
timestamp 1712078602
transform 1 0 141910 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_3079
timestamp 1712078602
transform 1 0 142186 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3081
timestamp 1712078602
transform 1 0 142278 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3093
timestamp 1712078602
transform 1 0 142830 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3105
timestamp 1712078602
transform 1 0 143382 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3117
timestamp 1712078602
transform 1 0 143934 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_3129
timestamp 1712078602
transform 1 0 144486 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_3135
timestamp 1712078602
transform 1 0 144762 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3137
timestamp 1712078602
transform 1 0 144854 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3149
timestamp 1712078602
transform 1 0 145406 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3161
timestamp 1712078602
transform 1 0 145958 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3173
timestamp 1712078602
transform 1 0 146510 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_3185
timestamp 1712078602
transform 1 0 147062 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_3191
timestamp 1712078602
transform 1 0 147338 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3193
timestamp 1712078602
transform 1 0 147430 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3205
timestamp 1712078602
transform 1 0 147982 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3217
timestamp 1712078602
transform 1 0 148534 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3229
timestamp 1712078602
transform 1 0 149086 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_3241
timestamp 1712078602
transform 1 0 149638 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_3247
timestamp 1712078602
transform 1 0 149914 0 -1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3249
timestamp 1712078602
transform 1 0 150006 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3261
timestamp 1712078602
transform 1 0 150558 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3273
timestamp 1712078602
transform 1 0 151110 0 -1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_5_3285
timestamp 1712078602
transform 1 0 151662 0 -1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_5_3297
timestamp 1712078602
transform 1 0 152214 0 -1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_5_3303
timestamp 1712078602
transform 1 0 152490 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_5_3305
timestamp 1712078602
transform 1 0 152582 0 -1 2720
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1712078602
transform 1 0 690 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1712078602
transform 1 0 1242 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1712078602
transform 1 0 1794 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1712078602
transform 1 0 1886 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1712078602
transform 1 0 2438 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1712078602
transform 1 0 2990 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1712078602
transform 1 0 3542 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1712078602
transform 1 0 4094 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1712078602
transform 1 0 4370 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1712078602
transform 1 0 4462 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1712078602
transform 1 0 5014 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1712078602
transform 1 0 5566 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1712078602
transform 1 0 6118 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1712078602
transform 1 0 6670 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1712078602
transform 1 0 6946 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1712078602
transform 1 0 7038 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1712078602
transform 1 0 7590 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1712078602
transform 1 0 8142 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1712078602
transform 1 0 8694 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1712078602
transform 1 0 9246 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1712078602
transform 1 0 9522 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1712078602
transform 1 0 9614 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1712078602
transform 1 0 10166 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1712078602
transform 1 0 10718 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1712078602
transform 1 0 11270 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1712078602
transform 1 0 11822 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1712078602
transform 1 0 12098 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1712078602
transform 1 0 12190 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1712078602
transform 1 0 12742 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1712078602
transform 1 0 13294 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1712078602
transform 1 0 13846 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1712078602
transform 1 0 14398 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1712078602
transform 1 0 14674 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1712078602
transform 1 0 14766 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1712078602
transform 1 0 15318 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1712078602
transform 1 0 15870 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1712078602
transform 1 0 16422 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1712078602
transform 1 0 16974 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1712078602
transform 1 0 17250 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1712078602
transform 1 0 17342 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1712078602
transform 1 0 17894 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1712078602
transform 1 0 18446 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1712078602
transform 1 0 18998 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1712078602
transform 1 0 19550 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1712078602
transform 1 0 19826 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1712078602
transform 1 0 19918 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1712078602
transform 1 0 20470 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1712078602
transform 1 0 21022 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1712078602
transform 1 0 21574 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1712078602
transform 1 0 22126 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1712078602
transform 1 0 22402 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1712078602
transform 1 0 22494 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1712078602
transform 1 0 23046 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1712078602
transform 1 0 23598 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1712078602
transform 1 0 24150 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1712078602
transform 1 0 24702 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1712078602
transform 1 0 24978 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1712078602
transform 1 0 25070 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1712078602
transform 1 0 25622 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1712078602
transform 1 0 26174 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1712078602
transform 1 0 26726 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1712078602
transform 1 0 27278 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1712078602
transform 1 0 27554 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1712078602
transform 1 0 27646 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1712078602
transform 1 0 28198 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1712078602
transform 1 0 28750 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1712078602
transform 1 0 29302 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1712078602
transform 1 0 29854 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1712078602
transform 1 0 30130 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1712078602
transform 1 0 30222 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1712078602
transform 1 0 30774 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1712078602
transform 1 0 31326 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1712078602
transform 1 0 31878 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1712078602
transform 1 0 32430 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1712078602
transform 1 0 32706 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1712078602
transform 1 0 32798 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1712078602
transform 1 0 33350 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1712078602
transform 1 0 33902 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1712078602
transform 1 0 34454 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1712078602
transform 1 0 35006 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1712078602
transform 1 0 35282 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1712078602
transform 1 0 35374 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1712078602
transform 1 0 35926 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1712078602
transform 1 0 36478 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1712078602
transform 1 0 37030 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1712078602
transform 1 0 37582 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1712078602
transform 1 0 37858 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1712078602
transform 1 0 37950 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1712078602
transform 1 0 38502 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1712078602
transform 1 0 39054 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1712078602
transform 1 0 39606 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1712078602
transform 1 0 40158 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1712078602
transform 1 0 40434 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1712078602
transform 1 0 40526 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1712078602
transform 1 0 41078 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1712078602
transform 1 0 41630 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1712078602
transform 1 0 42182 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1712078602
transform 1 0 42734 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1712078602
transform 1 0 43010 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1712078602
transform 1 0 43102 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1712078602
transform 1 0 43654 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1712078602
transform 1 0 44206 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1712078602
transform 1 0 44758 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1712078602
transform 1 0 45310 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1712078602
transform 1 0 45586 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1712078602
transform 1 0 45678 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1712078602
transform 1 0 46230 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1712078602
transform 1 0 46782 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1712078602
transform 1 0 47334 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1712078602
transform 1 0 47886 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1712078602
transform 1 0 48162 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1712078602
transform 1 0 48254 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1712078602
transform 1 0 48806 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1712078602
transform 1 0 49358 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1712078602
transform 1 0 49910 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1712078602
transform 1 0 50462 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1712078602
transform 1 0 50738 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1712078602
transform 1 0 50830 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1712078602
transform 1 0 51382 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1712078602
transform 1 0 51934 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1712078602
transform 1 0 52486 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1712078602
transform 1 0 53038 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1712078602
transform 1 0 53314 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1712078602
transform 1 0 53406 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1712078602
transform 1 0 53958 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1712078602
transform 1 0 54510 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1712078602
transform 1 0 55062 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1712078602
transform 1 0 55614 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1712078602
transform 1 0 55890 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1712078602
transform 1 0 55982 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1712078602
transform 1 0 56534 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1712078602
transform 1 0 57086 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1712078602
transform 1 0 57638 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1712078602
transform 1 0 58190 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1712078602
transform 1 0 58466 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1712078602
transform 1 0 58558 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1273
timestamp 1712078602
transform 1 0 59110 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1285
timestamp 1712078602
transform 1 0 59662 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1297
timestamp 1712078602
transform 1 0 60214 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1309
timestamp 1712078602
transform 1 0 60766 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1315
timestamp 1712078602
transform 1 0 61042 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1317
timestamp 1712078602
transform 1 0 61134 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1329
timestamp 1712078602
transform 1 0 61686 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1341
timestamp 1712078602
transform 1 0 62238 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1353
timestamp 1712078602
transform 1 0 62790 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1365
timestamp 1712078602
transform 1 0 63342 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1371
timestamp 1712078602
transform 1 0 63618 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1373
timestamp 1712078602
transform 1 0 63710 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1385
timestamp 1712078602
transform 1 0 64262 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1397
timestamp 1712078602
transform 1 0 64814 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1409
timestamp 1712078602
transform 1 0 65366 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1421
timestamp 1712078602
transform 1 0 65918 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1427
timestamp 1712078602
transform 1 0 66194 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1429
timestamp 1712078602
transform 1 0 66286 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1441
timestamp 1712078602
transform 1 0 66838 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1453
timestamp 1712078602
transform 1 0 67390 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1465
timestamp 1712078602
transform 1 0 67942 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1477
timestamp 1712078602
transform 1 0 68494 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1483
timestamp 1712078602
transform 1 0 68770 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1485
timestamp 1712078602
transform 1 0 68862 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1497
timestamp 1712078602
transform 1 0 69414 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1509
timestamp 1712078602
transform 1 0 69966 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1521
timestamp 1712078602
transform 1 0 70518 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1712078602
transform 1 0 71070 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1712078602
transform 1 0 71346 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1712078602
transform 1 0 71438 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1712078602
transform 1 0 71990 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1712078602
transform 1 0 72542 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1712078602
transform 1 0 73094 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1712078602
transform 1 0 73646 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1712078602
transform 1 0 73922 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1597
timestamp 1712078602
transform 1 0 74014 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1609
timestamp 1712078602
transform 1 0 74566 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1621
timestamp 1712078602
transform 1 0 75118 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1633
timestamp 1712078602
transform 1 0 75670 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1645
timestamp 1712078602
transform 1 0 76222 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1651
timestamp 1712078602
transform 1 0 76498 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1653
timestamp 1712078602
transform 1 0 76590 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1665
timestamp 1712078602
transform 1 0 77142 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1677
timestamp 1712078602
transform 1 0 77694 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1689
timestamp 1712078602
transform 1 0 78246 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1701
timestamp 1712078602
transform 1 0 78798 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1707
timestamp 1712078602
transform 1 0 79074 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1709
timestamp 1712078602
transform 1 0 79166 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1721
timestamp 1712078602
transform 1 0 79718 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1733
timestamp 1712078602
transform 1 0 80270 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1745
timestamp 1712078602
transform 1 0 80822 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1757
timestamp 1712078602
transform 1 0 81374 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1763
timestamp 1712078602
transform 1 0 81650 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1765
timestamp 1712078602
transform 1 0 81742 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1777
timestamp 1712078602
transform 1 0 82294 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1789
timestamp 1712078602
transform 1 0 82846 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1801
timestamp 1712078602
transform 1 0 83398 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1813
timestamp 1712078602
transform 1 0 83950 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1819
timestamp 1712078602
transform 1 0 84226 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1821
timestamp 1712078602
transform 1 0 84318 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1833
timestamp 1712078602
transform 1 0 84870 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1845
timestamp 1712078602
transform 1 0 85422 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1857
timestamp 1712078602
transform 1 0 85974 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1869
timestamp 1712078602
transform 1 0 86526 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1875
timestamp 1712078602
transform 1 0 86802 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1877
timestamp 1712078602
transform 1 0 86894 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1889
timestamp 1712078602
transform 1 0 87446 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1901
timestamp 1712078602
transform 1 0 87998 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1913
timestamp 1712078602
transform 1 0 88550 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1925
timestamp 1712078602
transform 1 0 89102 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1931
timestamp 1712078602
transform 1 0 89378 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1933
timestamp 1712078602
transform 1 0 89470 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1945
timestamp 1712078602
transform 1 0 90022 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1957
timestamp 1712078602
transform 1 0 90574 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1969
timestamp 1712078602
transform 1 0 91126 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_1981
timestamp 1712078602
transform 1 0 91678 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_1987
timestamp 1712078602
transform 1 0 91954 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_1989
timestamp 1712078602
transform 1 0 92046 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2001
timestamp 1712078602
transform 1 0 92598 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2013
timestamp 1712078602
transform 1 0 93150 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2025
timestamp 1712078602
transform 1 0 93702 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2037
timestamp 1712078602
transform 1 0 94254 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2043
timestamp 1712078602
transform 1 0 94530 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2045
timestamp 1712078602
transform 1 0 94622 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2057
timestamp 1712078602
transform 1 0 95174 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2069
timestamp 1712078602
transform 1 0 95726 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2081
timestamp 1712078602
transform 1 0 96278 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2093
timestamp 1712078602
transform 1 0 96830 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2099
timestamp 1712078602
transform 1 0 97106 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2101
timestamp 1712078602
transform 1 0 97198 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2113
timestamp 1712078602
transform 1 0 97750 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2125
timestamp 1712078602
transform 1 0 98302 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2137
timestamp 1712078602
transform 1 0 98854 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2149
timestamp 1712078602
transform 1 0 99406 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2155
timestamp 1712078602
transform 1 0 99682 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2157
timestamp 1712078602
transform 1 0 99774 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2169
timestamp 1712078602
transform 1 0 100326 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2181
timestamp 1712078602
transform 1 0 100878 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2193
timestamp 1712078602
transform 1 0 101430 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2205
timestamp 1712078602
transform 1 0 101982 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2211
timestamp 1712078602
transform 1 0 102258 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2213
timestamp 1712078602
transform 1 0 102350 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2225
timestamp 1712078602
transform 1 0 102902 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2237
timestamp 1712078602
transform 1 0 103454 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2249
timestamp 1712078602
transform 1 0 104006 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2261
timestamp 1712078602
transform 1 0 104558 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2267
timestamp 1712078602
transform 1 0 104834 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2269
timestamp 1712078602
transform 1 0 104926 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2281
timestamp 1712078602
transform 1 0 105478 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2293
timestamp 1712078602
transform 1 0 106030 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2305
timestamp 1712078602
transform 1 0 106582 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2317
timestamp 1712078602
transform 1 0 107134 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2323
timestamp 1712078602
transform 1 0 107410 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2325
timestamp 1712078602
transform 1 0 107502 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2337
timestamp 1712078602
transform 1 0 108054 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2349
timestamp 1712078602
transform 1 0 108606 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2361
timestamp 1712078602
transform 1 0 109158 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2373
timestamp 1712078602
transform 1 0 109710 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2379
timestamp 1712078602
transform 1 0 109986 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2381
timestamp 1712078602
transform 1 0 110078 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2393
timestamp 1712078602
transform 1 0 110630 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2405
timestamp 1712078602
transform 1 0 111182 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2417
timestamp 1712078602
transform 1 0 111734 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2429
timestamp 1712078602
transform 1 0 112286 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2435
timestamp 1712078602
transform 1 0 112562 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2437
timestamp 1712078602
transform 1 0 112654 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2449
timestamp 1712078602
transform 1 0 113206 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2461
timestamp 1712078602
transform 1 0 113758 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2473
timestamp 1712078602
transform 1 0 114310 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2485
timestamp 1712078602
transform 1 0 114862 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2491
timestamp 1712078602
transform 1 0 115138 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2493
timestamp 1712078602
transform 1 0 115230 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2505
timestamp 1712078602
transform 1 0 115782 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2517
timestamp 1712078602
transform 1 0 116334 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2529
timestamp 1712078602
transform 1 0 116886 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2541
timestamp 1712078602
transform 1 0 117438 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2547
timestamp 1712078602
transform 1 0 117714 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2549
timestamp 1712078602
transform 1 0 117806 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2561
timestamp 1712078602
transform 1 0 118358 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2573
timestamp 1712078602
transform 1 0 118910 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2585
timestamp 1712078602
transform 1 0 119462 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2597
timestamp 1712078602
transform 1 0 120014 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2603
timestamp 1712078602
transform 1 0 120290 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2605
timestamp 1712078602
transform 1 0 120382 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2617
timestamp 1712078602
transform 1 0 120934 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2629
timestamp 1712078602
transform 1 0 121486 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2641
timestamp 1712078602
transform 1 0 122038 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2653
timestamp 1712078602
transform 1 0 122590 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2659
timestamp 1712078602
transform 1 0 122866 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2661
timestamp 1712078602
transform 1 0 122958 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2673
timestamp 1712078602
transform 1 0 123510 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2685
timestamp 1712078602
transform 1 0 124062 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2697
timestamp 1712078602
transform 1 0 124614 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2709
timestamp 1712078602
transform 1 0 125166 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2715
timestamp 1712078602
transform 1 0 125442 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2717
timestamp 1712078602
transform 1 0 125534 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2729
timestamp 1712078602
transform 1 0 126086 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2741
timestamp 1712078602
transform 1 0 126638 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2753
timestamp 1712078602
transform 1 0 127190 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2765
timestamp 1712078602
transform 1 0 127742 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2771
timestamp 1712078602
transform 1 0 128018 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2773
timestamp 1712078602
transform 1 0 128110 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2785
timestamp 1712078602
transform 1 0 128662 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2797
timestamp 1712078602
transform 1 0 129214 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2809
timestamp 1712078602
transform 1 0 129766 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2821
timestamp 1712078602
transform 1 0 130318 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2827
timestamp 1712078602
transform 1 0 130594 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2829
timestamp 1712078602
transform 1 0 130686 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2841
timestamp 1712078602
transform 1 0 131238 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2853
timestamp 1712078602
transform 1 0 131790 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2865
timestamp 1712078602
transform 1 0 132342 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2877
timestamp 1712078602
transform 1 0 132894 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2883
timestamp 1712078602
transform 1 0 133170 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2885
timestamp 1712078602
transform 1 0 133262 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2897
timestamp 1712078602
transform 1 0 133814 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2909
timestamp 1712078602
transform 1 0 134366 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2921
timestamp 1712078602
transform 1 0 134918 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2933
timestamp 1712078602
transform 1 0 135470 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2939
timestamp 1712078602
transform 1 0 135746 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2941
timestamp 1712078602
transform 1 0 135838 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2953
timestamp 1712078602
transform 1 0 136390 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2965
timestamp 1712078602
transform 1 0 136942 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2977
timestamp 1712078602
transform 1 0 137494 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_2989
timestamp 1712078602
transform 1 0 138046 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_2995
timestamp 1712078602
transform 1 0 138322 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_2997
timestamp 1712078602
transform 1 0 138414 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3009
timestamp 1712078602
transform 1 0 138966 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3021
timestamp 1712078602
transform 1 0 139518 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3033
timestamp 1712078602
transform 1 0 140070 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_3045
timestamp 1712078602
transform 1 0 140622 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_3051
timestamp 1712078602
transform 1 0 140898 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3053
timestamp 1712078602
transform 1 0 140990 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3065
timestamp 1712078602
transform 1 0 141542 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3077
timestamp 1712078602
transform 1 0 142094 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3089
timestamp 1712078602
transform 1 0 142646 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_3101
timestamp 1712078602
transform 1 0 143198 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_3107
timestamp 1712078602
transform 1 0 143474 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3109
timestamp 1712078602
transform 1 0 143566 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3121
timestamp 1712078602
transform 1 0 144118 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3133
timestamp 1712078602
transform 1 0 144670 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3145
timestamp 1712078602
transform 1 0 145222 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_3157
timestamp 1712078602
transform 1 0 145774 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_3163
timestamp 1712078602
transform 1 0 146050 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3165
timestamp 1712078602
transform 1 0 146142 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3177
timestamp 1712078602
transform 1 0 146694 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3189
timestamp 1712078602
transform 1 0 147246 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3201
timestamp 1712078602
transform 1 0 147798 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_3213
timestamp 1712078602
transform 1 0 148350 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_3219
timestamp 1712078602
transform 1 0 148626 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3221
timestamp 1712078602
transform 1 0 148718 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3233
timestamp 1712078602
transform 1 0 149270 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3245
timestamp 1712078602
transform 1 0 149822 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3257
timestamp 1712078602
transform 1 0 150374 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_6_3269
timestamp 1712078602
transform 1 0 150926 0 1 2720
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_6_3275
timestamp 1712078602
transform 1 0 151202 0 1 2720
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3277
timestamp 1712078602
transform 1 0 151294 0 1 2720
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_6_3289
timestamp 1712078602
transform 1 0 151846 0 1 2720
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_6_3301
timestamp 1712078602
transform 1 0 152398 0 1 2720
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1712078602
transform 1 0 690 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1712078602
transform 1 0 1242 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1712078602
transform 1 0 1794 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1712078602
transform 1 0 2346 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1712078602
transform 1 0 2898 0 -1 3264
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1712078602
transform 1 0 3082 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1712078602
transform 1 0 3174 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1712078602
transform 1 0 3726 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1712078602
transform 1 0 4278 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1712078602
transform 1 0 4830 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1712078602
transform 1 0 5382 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1712078602
transform 1 0 5658 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1712078602
transform 1 0 5750 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1712078602
transform 1 0 6302 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1712078602
transform 1 0 6854 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1712078602
transform 1 0 7406 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1712078602
transform 1 0 7958 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1712078602
transform 1 0 8234 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1712078602
transform 1 0 8326 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1712078602
transform 1 0 8878 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1712078602
transform 1 0 9430 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1712078602
transform 1 0 9982 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1712078602
transform 1 0 10534 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1712078602
transform 1 0 10810 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1712078602
transform 1 0 10902 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1712078602
transform 1 0 11454 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1712078602
transform 1 0 12006 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1712078602
transform 1 0 12558 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1712078602
transform 1 0 13110 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1712078602
transform 1 0 13386 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1712078602
transform 1 0 13478 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1712078602
transform 1 0 14030 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1712078602
transform 1 0 14582 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1712078602
transform 1 0 15134 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1712078602
transform 1 0 15686 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1712078602
transform 1 0 15962 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1712078602
transform 1 0 16054 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1712078602
transform 1 0 16606 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1712078602
transform 1 0 17158 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1712078602
transform 1 0 17710 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1712078602
transform 1 0 18262 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1712078602
transform 1 0 18538 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1712078602
transform 1 0 18630 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1712078602
transform 1 0 19182 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1712078602
transform 1 0 19734 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1712078602
transform 1 0 20286 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1712078602
transform 1 0 20838 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1712078602
transform 1 0 21114 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1712078602
transform 1 0 21206 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1712078602
transform 1 0 21758 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1712078602
transform 1 0 22310 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1712078602
transform 1 0 22862 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1712078602
transform 1 0 23414 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1712078602
transform 1 0 23690 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1712078602
transform 1 0 23782 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1712078602
transform 1 0 24334 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1712078602
transform 1 0 24886 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1712078602
transform 1 0 25438 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1712078602
transform 1 0 25990 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1712078602
transform 1 0 26266 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1712078602
transform 1 0 26358 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1712078602
transform 1 0 26910 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1712078602
transform 1 0 27462 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1712078602
transform 1 0 28014 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1712078602
transform 1 0 28566 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1712078602
transform 1 0 28842 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1712078602
transform 1 0 28934 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1712078602
transform 1 0 29486 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1712078602
transform 1 0 30038 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1712078602
transform 1 0 30590 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1712078602
transform 1 0 31142 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1712078602
transform 1 0 31418 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1712078602
transform 1 0 31510 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1712078602
transform 1 0 32062 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1712078602
transform 1 0 32614 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1712078602
transform 1 0 33166 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1712078602
transform 1 0 33718 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1712078602
transform 1 0 33994 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1712078602
transform 1 0 34086 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1712078602
transform 1 0 34638 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1712078602
transform 1 0 35190 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1712078602
transform 1 0 35742 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1712078602
transform 1 0 36294 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1712078602
transform 1 0 36570 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1712078602
transform 1 0 36662 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1712078602
transform 1 0 37214 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1712078602
transform 1 0 37766 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1712078602
transform 1 0 38318 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1712078602
transform 1 0 38870 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1712078602
transform 1 0 39146 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1712078602
transform 1 0 39238 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1712078602
transform 1 0 39790 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1712078602
transform 1 0 40342 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1712078602
transform 1 0 40894 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1712078602
transform 1 0 41446 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1712078602
transform 1 0 41722 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1712078602
transform 1 0 41814 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1712078602
transform 1 0 42366 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1712078602
transform 1 0 42918 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1712078602
transform 1 0 43470 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1712078602
transform 1 0 44022 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1712078602
transform 1 0 44298 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1712078602
transform 1 0 44390 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1712078602
transform 1 0 44942 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1712078602
transform 1 0 45494 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1712078602
transform 1 0 46046 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1712078602
transform 1 0 46598 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1712078602
transform 1 0 46874 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1712078602
transform 1 0 46966 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1712078602
transform 1 0 47518 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1712078602
transform 1 0 48070 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1712078602
transform 1 0 48622 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1712078602
transform 1 0 49174 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1712078602
transform 1 0 49450 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1712078602
transform 1 0 49542 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1712078602
transform 1 0 50094 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1712078602
transform 1 0 50646 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1712078602
transform 1 0 51198 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1712078602
transform 1 0 51750 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1712078602
transform 1 0 52026 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1712078602
transform 1 0 52118 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1712078602
transform 1 0 52670 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1712078602
transform 1 0 53222 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1712078602
transform 1 0 53774 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1712078602
transform 1 0 54326 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1712078602
transform 1 0 54602 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1712078602
transform 1 0 54694 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1712078602
transform 1 0 55246 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1712078602
transform 1 0 55798 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1712078602
transform 1 0 56350 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1712078602
transform 1 0 56902 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1712078602
transform 1 0 57178 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1712078602
transform 1 0 57270 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1712078602
transform 1 0 57822 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1712078602
transform 1 0 58374 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1269
timestamp 1712078602
transform 1 0 58926 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1281
timestamp 1712078602
transform 1 0 59478 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1287
timestamp 1712078602
transform 1 0 59754 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1289
timestamp 1712078602
transform 1 0 59846 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1301
timestamp 1712078602
transform 1 0 60398 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1313
timestamp 1712078602
transform 1 0 60950 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1325
timestamp 1712078602
transform 1 0 61502 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1337
timestamp 1712078602
transform 1 0 62054 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1343
timestamp 1712078602
transform 1 0 62330 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1345
timestamp 1712078602
transform 1 0 62422 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1357
timestamp 1712078602
transform 1 0 62974 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1369
timestamp 1712078602
transform 1 0 63526 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1381
timestamp 1712078602
transform 1 0 64078 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1393
timestamp 1712078602
transform 1 0 64630 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1399
timestamp 1712078602
transform 1 0 64906 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1712078602
transform 1 0 64998 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1413
timestamp 1712078602
transform 1 0 65550 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1425
timestamp 1712078602
transform 1 0 66102 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1437
timestamp 1712078602
transform 1 0 66654 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1449
timestamp 1712078602
transform 1 0 67206 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1455
timestamp 1712078602
transform 1 0 67482 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1712078602
transform 1 0 67574 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1712078602
transform 1 0 68126 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1712078602
transform 1 0 68678 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1712078602
transform 1 0 69230 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1712078602
transform 1 0 69782 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1712078602
transform 1 0 70058 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1712078602
transform 1 0 70150 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1712078602
transform 1 0 70702 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1712078602
transform 1 0 71254 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1712078602
transform 1 0 71806 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1712078602
transform 1 0 72358 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1712078602
transform 1 0 72634 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1712078602
transform 1 0 72726 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1712078602
transform 1 0 73278 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1593
timestamp 1712078602
transform 1 0 73830 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1605
timestamp 1712078602
transform 1 0 74382 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1617
timestamp 1712078602
transform 1 0 74934 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1712078602
transform 1 0 75210 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1625
timestamp 1712078602
transform 1 0 75302 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1637
timestamp 1712078602
transform 1 0 75854 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1649
timestamp 1712078602
transform 1 0 76406 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1661
timestamp 1712078602
transform 1 0 76958 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1673
timestamp 1712078602
transform 1 0 77510 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1712078602
transform 1 0 77786 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1681
timestamp 1712078602
transform 1 0 77878 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1693
timestamp 1712078602
transform 1 0 78430 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1705
timestamp 1712078602
transform 1 0 78982 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1717
timestamp 1712078602
transform 1 0 79534 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1729
timestamp 1712078602
transform 1 0 80086 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1735
timestamp 1712078602
transform 1 0 80362 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1737
timestamp 1712078602
transform 1 0 80454 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1749
timestamp 1712078602
transform 1 0 81006 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1761
timestamp 1712078602
transform 1 0 81558 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1773
timestamp 1712078602
transform 1 0 82110 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1785
timestamp 1712078602
transform 1 0 82662 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1791
timestamp 1712078602
transform 1 0 82938 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1793
timestamp 1712078602
transform 1 0 83030 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1805
timestamp 1712078602
transform 1 0 83582 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1817
timestamp 1712078602
transform 1 0 84134 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1829
timestamp 1712078602
transform 1 0 84686 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1841
timestamp 1712078602
transform 1 0 85238 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1847
timestamp 1712078602
transform 1 0 85514 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1849
timestamp 1712078602
transform 1 0 85606 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1861
timestamp 1712078602
transform 1 0 86158 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1873
timestamp 1712078602
transform 1 0 86710 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1885
timestamp 1712078602
transform 1 0 87262 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1897
timestamp 1712078602
transform 1 0 87814 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1903
timestamp 1712078602
transform 1 0 88090 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1905
timestamp 1712078602
transform 1 0 88182 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1917
timestamp 1712078602
transform 1 0 88734 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1929
timestamp 1712078602
transform 1 0 89286 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1941
timestamp 1712078602
transform 1 0 89838 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_1953
timestamp 1712078602
transform 1 0 90390 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_1959
timestamp 1712078602
transform 1 0 90666 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1961
timestamp 1712078602
transform 1 0 90758 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1973
timestamp 1712078602
transform 1 0 91310 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1985
timestamp 1712078602
transform 1 0 91862 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_1997
timestamp 1712078602
transform 1 0 92414 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2009
timestamp 1712078602
transform 1 0 92966 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2015
timestamp 1712078602
transform 1 0 93242 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2017
timestamp 1712078602
transform 1 0 93334 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2029
timestamp 1712078602
transform 1 0 93886 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2041
timestamp 1712078602
transform 1 0 94438 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2053
timestamp 1712078602
transform 1 0 94990 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2065
timestamp 1712078602
transform 1 0 95542 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2071
timestamp 1712078602
transform 1 0 95818 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2073
timestamp 1712078602
transform 1 0 95910 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2085
timestamp 1712078602
transform 1 0 96462 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2097
timestamp 1712078602
transform 1 0 97014 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2109
timestamp 1712078602
transform 1 0 97566 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2121
timestamp 1712078602
transform 1 0 98118 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2127
timestamp 1712078602
transform 1 0 98394 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2129
timestamp 1712078602
transform 1 0 98486 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2141
timestamp 1712078602
transform 1 0 99038 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2153
timestamp 1712078602
transform 1 0 99590 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2165
timestamp 1712078602
transform 1 0 100142 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2177
timestamp 1712078602
transform 1 0 100694 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2183
timestamp 1712078602
transform 1 0 100970 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2185
timestamp 1712078602
transform 1 0 101062 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2197
timestamp 1712078602
transform 1 0 101614 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2209
timestamp 1712078602
transform 1 0 102166 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2221
timestamp 1712078602
transform 1 0 102718 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2233
timestamp 1712078602
transform 1 0 103270 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2239
timestamp 1712078602
transform 1 0 103546 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2241
timestamp 1712078602
transform 1 0 103638 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2253
timestamp 1712078602
transform 1 0 104190 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2265
timestamp 1712078602
transform 1 0 104742 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2277
timestamp 1712078602
transform 1 0 105294 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2289
timestamp 1712078602
transform 1 0 105846 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2295
timestamp 1712078602
transform 1 0 106122 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2297
timestamp 1712078602
transform 1 0 106214 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2309
timestamp 1712078602
transform 1 0 106766 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2321
timestamp 1712078602
transform 1 0 107318 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2333
timestamp 1712078602
transform 1 0 107870 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2345
timestamp 1712078602
transform 1 0 108422 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2351
timestamp 1712078602
transform 1 0 108698 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2353
timestamp 1712078602
transform 1 0 108790 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2365
timestamp 1712078602
transform 1 0 109342 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2377
timestamp 1712078602
transform 1 0 109894 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2389
timestamp 1712078602
transform 1 0 110446 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2401
timestamp 1712078602
transform 1 0 110998 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2407
timestamp 1712078602
transform 1 0 111274 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2409
timestamp 1712078602
transform 1 0 111366 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2421
timestamp 1712078602
transform 1 0 111918 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2433
timestamp 1712078602
transform 1 0 112470 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2445
timestamp 1712078602
transform 1 0 113022 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2457
timestamp 1712078602
transform 1 0 113574 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2463
timestamp 1712078602
transform 1 0 113850 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2465
timestamp 1712078602
transform 1 0 113942 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2477
timestamp 1712078602
transform 1 0 114494 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2489
timestamp 1712078602
transform 1 0 115046 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2501
timestamp 1712078602
transform 1 0 115598 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2513
timestamp 1712078602
transform 1 0 116150 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2519
timestamp 1712078602
transform 1 0 116426 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2521
timestamp 1712078602
transform 1 0 116518 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2533
timestamp 1712078602
transform 1 0 117070 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2545
timestamp 1712078602
transform 1 0 117622 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2557
timestamp 1712078602
transform 1 0 118174 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2569
timestamp 1712078602
transform 1 0 118726 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2575
timestamp 1712078602
transform 1 0 119002 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2577
timestamp 1712078602
transform 1 0 119094 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2589
timestamp 1712078602
transform 1 0 119646 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2601
timestamp 1712078602
transform 1 0 120198 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2613
timestamp 1712078602
transform 1 0 120750 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2625
timestamp 1712078602
transform 1 0 121302 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2631
timestamp 1712078602
transform 1 0 121578 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2633
timestamp 1712078602
transform 1 0 121670 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2645
timestamp 1712078602
transform 1 0 122222 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2657
timestamp 1712078602
transform 1 0 122774 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2669
timestamp 1712078602
transform 1 0 123326 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2681
timestamp 1712078602
transform 1 0 123878 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2687
timestamp 1712078602
transform 1 0 124154 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2689
timestamp 1712078602
transform 1 0 124246 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2701
timestamp 1712078602
transform 1 0 124798 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2713
timestamp 1712078602
transform 1 0 125350 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2725
timestamp 1712078602
transform 1 0 125902 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2737
timestamp 1712078602
transform 1 0 126454 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2743
timestamp 1712078602
transform 1 0 126730 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2745
timestamp 1712078602
transform 1 0 126822 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2757
timestamp 1712078602
transform 1 0 127374 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2769
timestamp 1712078602
transform 1 0 127926 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2781
timestamp 1712078602
transform 1 0 128478 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2793
timestamp 1712078602
transform 1 0 129030 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2799
timestamp 1712078602
transform 1 0 129306 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2801
timestamp 1712078602
transform 1 0 129398 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2813
timestamp 1712078602
transform 1 0 129950 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2825
timestamp 1712078602
transform 1 0 130502 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2837
timestamp 1712078602
transform 1 0 131054 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2849
timestamp 1712078602
transform 1 0 131606 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2855
timestamp 1712078602
transform 1 0 131882 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2857
timestamp 1712078602
transform 1 0 131974 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2869
timestamp 1712078602
transform 1 0 132526 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2881
timestamp 1712078602
transform 1 0 133078 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2893
timestamp 1712078602
transform 1 0 133630 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2905
timestamp 1712078602
transform 1 0 134182 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2911
timestamp 1712078602
transform 1 0 134458 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2913
timestamp 1712078602
transform 1 0 134550 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2925
timestamp 1712078602
transform 1 0 135102 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2937
timestamp 1712078602
transform 1 0 135654 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2949
timestamp 1712078602
transform 1 0 136206 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_2961
timestamp 1712078602
transform 1 0 136758 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_2967
timestamp 1712078602
transform 1 0 137034 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2969
timestamp 1712078602
transform 1 0 137126 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2981
timestamp 1712078602
transform 1 0 137678 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_2993
timestamp 1712078602
transform 1 0 138230 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3005
timestamp 1712078602
transform 1 0 138782 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_3017
timestamp 1712078602
transform 1 0 139334 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_3023
timestamp 1712078602
transform 1 0 139610 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3025
timestamp 1712078602
transform 1 0 139702 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3037
timestamp 1712078602
transform 1 0 140254 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3049
timestamp 1712078602
transform 1 0 140806 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3061
timestamp 1712078602
transform 1 0 141358 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_3073
timestamp 1712078602
transform 1 0 141910 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_3079
timestamp 1712078602
transform 1 0 142186 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3081
timestamp 1712078602
transform 1 0 142278 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3093
timestamp 1712078602
transform 1 0 142830 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3105
timestamp 1712078602
transform 1 0 143382 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3117
timestamp 1712078602
transform 1 0 143934 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_3129
timestamp 1712078602
transform 1 0 144486 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_3135
timestamp 1712078602
transform 1 0 144762 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3137
timestamp 1712078602
transform 1 0 144854 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3149
timestamp 1712078602
transform 1 0 145406 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3161
timestamp 1712078602
transform 1 0 145958 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3173
timestamp 1712078602
transform 1 0 146510 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_3185
timestamp 1712078602
transform 1 0 147062 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_3191
timestamp 1712078602
transform 1 0 147338 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3193
timestamp 1712078602
transform 1 0 147430 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3205
timestamp 1712078602
transform 1 0 147982 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3217
timestamp 1712078602
transform 1 0 148534 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3229
timestamp 1712078602
transform 1 0 149086 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_3241
timestamp 1712078602
transform 1 0 149638 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_7_3247
timestamp 1712078602
transform 1 0 149914 0 -1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3249
timestamp 1712078602
transform 1 0 150006 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3261
timestamp 1712078602
transform 1 0 150558 0 -1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_7_3273
timestamp 1712078602
transform 1 0 151110 0 -1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_7_3285
timestamp 1712078602
transform 1 0 151662 0 -1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_7_3300
timestamp 1712078602
transform 1 0 152352 0 -1 3264
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_7_3305
timestamp 1712078602
transform 1 0 152582 0 -1 3264
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1712078602
transform 1 0 690 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1712078602
transform 1 0 1242 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1712078602
transform 1 0 1794 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1712078602
transform 1 0 1886 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1712078602
transform 1 0 2438 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1712078602
transform 1 0 2990 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1712078602
transform 1 0 3542 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1712078602
transform 1 0 4094 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1712078602
transform 1 0 4370 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1712078602
transform 1 0 4462 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1712078602
transform 1 0 5014 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1712078602
transform 1 0 5566 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1712078602
transform 1 0 6118 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1712078602
transform 1 0 6670 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1712078602
transform 1 0 6946 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1712078602
transform 1 0 7038 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1712078602
transform 1 0 7590 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1712078602
transform 1 0 8142 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1712078602
transform 1 0 8694 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1712078602
transform 1 0 9246 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1712078602
transform 1 0 9522 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1712078602
transform 1 0 9614 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1712078602
transform 1 0 10166 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1712078602
transform 1 0 10718 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1712078602
transform 1 0 11270 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1712078602
transform 1 0 11822 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1712078602
transform 1 0 12098 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1712078602
transform 1 0 12190 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1712078602
transform 1 0 12742 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1712078602
transform 1 0 13294 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1712078602
transform 1 0 13846 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1712078602
transform 1 0 14398 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1712078602
transform 1 0 14674 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1712078602
transform 1 0 14766 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1712078602
transform 1 0 15318 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1712078602
transform 1 0 15870 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1712078602
transform 1 0 16422 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1712078602
transform 1 0 16974 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1712078602
transform 1 0 17250 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1712078602
transform 1 0 17342 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1712078602
transform 1 0 17894 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1712078602
transform 1 0 18446 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1712078602
transform 1 0 18998 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1712078602
transform 1 0 19550 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1712078602
transform 1 0 19826 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1712078602
transform 1 0 19918 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1712078602
transform 1 0 20470 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1712078602
transform 1 0 21022 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1712078602
transform 1 0 21574 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1712078602
transform 1 0 22126 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1712078602
transform 1 0 22402 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1712078602
transform 1 0 22494 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1712078602
transform 1 0 23046 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1712078602
transform 1 0 23598 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1712078602
transform 1 0 24150 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1712078602
transform 1 0 24702 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1712078602
transform 1 0 24978 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1712078602
transform 1 0 25070 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1712078602
transform 1 0 25622 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1712078602
transform 1 0 26174 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1712078602
transform 1 0 26726 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1712078602
transform 1 0 27278 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1712078602
transform 1 0 27554 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1712078602
transform 1 0 27646 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1712078602
transform 1 0 28198 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1712078602
transform 1 0 28750 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1712078602
transform 1 0 29302 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1712078602
transform 1 0 29854 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1712078602
transform 1 0 30130 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1712078602
transform 1 0 30222 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1712078602
transform 1 0 30774 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1712078602
transform 1 0 31326 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1712078602
transform 1 0 31878 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1712078602
transform 1 0 32430 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1712078602
transform 1 0 32706 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1712078602
transform 1 0 32798 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1712078602
transform 1 0 33350 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1712078602
transform 1 0 33902 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1712078602
transform 1 0 34454 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1712078602
transform 1 0 35006 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1712078602
transform 1 0 35282 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1712078602
transform 1 0 35374 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1712078602
transform 1 0 35926 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1712078602
transform 1 0 36478 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1712078602
transform 1 0 37030 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1712078602
transform 1 0 37582 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1712078602
transform 1 0 37858 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1712078602
transform 1 0 37950 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1712078602
transform 1 0 38502 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1712078602
transform 1 0 39054 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1712078602
transform 1 0 39606 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1712078602
transform 1 0 40158 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1712078602
transform 1 0 40434 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1712078602
transform 1 0 40526 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1712078602
transform 1 0 41078 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1712078602
transform 1 0 41630 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1712078602
transform 1 0 42182 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1712078602
transform 1 0 42734 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1712078602
transform 1 0 43010 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1712078602
transform 1 0 43102 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1712078602
transform 1 0 43654 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1712078602
transform 1 0 44206 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1712078602
transform 1 0 44758 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1712078602
transform 1 0 45310 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1712078602
transform 1 0 45586 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1712078602
transform 1 0 45678 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1712078602
transform 1 0 46230 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1712078602
transform 1 0 46782 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1712078602
transform 1 0 47334 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1712078602
transform 1 0 47886 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1712078602
transform 1 0 48162 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1712078602
transform 1 0 48254 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1712078602
transform 1 0 48806 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1712078602
transform 1 0 49358 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1712078602
transform 1 0 49910 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1712078602
transform 1 0 50462 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1712078602
transform 1 0 50738 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1712078602
transform 1 0 50830 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1712078602
transform 1 0 51382 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1712078602
transform 1 0 51934 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1712078602
transform 1 0 52486 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1712078602
transform 1 0 53038 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1712078602
transform 1 0 53314 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1712078602
transform 1 0 53406 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1712078602
transform 1 0 53958 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1712078602
transform 1 0 54510 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1712078602
transform 1 0 55062 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1712078602
transform 1 0 55614 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1712078602
transform 1 0 55890 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1712078602
transform 1 0 55982 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1712078602
transform 1 0 56534 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1712078602
transform 1 0 57086 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1712078602
transform 1 0 57638 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1712078602
transform 1 0 58190 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1712078602
transform 1 0 58466 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1712078602
transform 1 0 58558 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1273
timestamp 1712078602
transform 1 0 59110 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1285
timestamp 1712078602
transform 1 0 59662 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1297
timestamp 1712078602
transform 1 0 60214 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1712078602
transform 1 0 60766 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1712078602
transform 1 0 61042 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1317
timestamp 1712078602
transform 1 0 61134 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1329
timestamp 1712078602
transform 1 0 61686 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1341
timestamp 1712078602
transform 1 0 62238 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1353
timestamp 1712078602
transform 1 0 62790 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1365
timestamp 1712078602
transform 1 0 63342 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1371
timestamp 1712078602
transform 1 0 63618 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1712078602
transform 1 0 63710 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1712078602
transform 1 0 64262 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1712078602
transform 1 0 64814 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1712078602
transform 1 0 65366 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1712078602
transform 1 0 65918 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1712078602
transform 1 0 66194 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1712078602
transform 1 0 66286 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1712078602
transform 1 0 66838 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1712078602
transform 1 0 67390 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1712078602
transform 1 0 67942 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1712078602
transform 1 0 68494 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1712078602
transform 1 0 68770 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1712078602
transform 1 0 68862 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1712078602
transform 1 0 69414 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1712078602
transform 1 0 69966 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1712078602
transform 1 0 70518 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1712078602
transform 1 0 71070 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1712078602
transform 1 0 71346 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1712078602
transform 1 0 71438 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1712078602
transform 1 0 71990 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1712078602
transform 1 0 72542 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1712078602
transform 1 0 73094 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1712078602
transform 1 0 73646 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1712078602
transform 1 0 73922 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1597
timestamp 1712078602
transform 1 0 74014 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1609
timestamp 1712078602
transform 1 0 74566 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1621
timestamp 1712078602
transform 1 0 75118 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1633
timestamp 1712078602
transform 1 0 75670 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1645
timestamp 1712078602
transform 1 0 76222 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1651
timestamp 1712078602
transform 1 0 76498 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1653
timestamp 1712078602
transform 1 0 76590 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1665
timestamp 1712078602
transform 1 0 77142 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1677
timestamp 1712078602
transform 1 0 77694 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1689
timestamp 1712078602
transform 1 0 78246 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1701
timestamp 1712078602
transform 1 0 78798 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1707
timestamp 1712078602
transform 1 0 79074 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1709
timestamp 1712078602
transform 1 0 79166 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1721
timestamp 1712078602
transform 1 0 79718 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1733
timestamp 1712078602
transform 1 0 80270 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1745
timestamp 1712078602
transform 1 0 80822 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1757
timestamp 1712078602
transform 1 0 81374 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1763
timestamp 1712078602
transform 1 0 81650 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1765
timestamp 1712078602
transform 1 0 81742 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1777
timestamp 1712078602
transform 1 0 82294 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1789
timestamp 1712078602
transform 1 0 82846 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1801
timestamp 1712078602
transform 1 0 83398 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1813
timestamp 1712078602
transform 1 0 83950 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1819
timestamp 1712078602
transform 1 0 84226 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1821
timestamp 1712078602
transform 1 0 84318 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1833
timestamp 1712078602
transform 1 0 84870 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1845
timestamp 1712078602
transform 1 0 85422 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1857
timestamp 1712078602
transform 1 0 85974 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1869
timestamp 1712078602
transform 1 0 86526 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1875
timestamp 1712078602
transform 1 0 86802 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1877
timestamp 1712078602
transform 1 0 86894 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1889
timestamp 1712078602
transform 1 0 87446 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1901
timestamp 1712078602
transform 1 0 87998 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1913
timestamp 1712078602
transform 1 0 88550 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1925
timestamp 1712078602
transform 1 0 89102 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1931
timestamp 1712078602
transform 1 0 89378 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1933
timestamp 1712078602
transform 1 0 89470 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1945
timestamp 1712078602
transform 1 0 90022 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1957
timestamp 1712078602
transform 1 0 90574 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1969
timestamp 1712078602
transform 1 0 91126 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_1981
timestamp 1712078602
transform 1 0 91678 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_1987
timestamp 1712078602
transform 1 0 91954 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_1989
timestamp 1712078602
transform 1 0 92046 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2001
timestamp 1712078602
transform 1 0 92598 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2013
timestamp 1712078602
transform 1 0 93150 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2025
timestamp 1712078602
transform 1 0 93702 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2037
timestamp 1712078602
transform 1 0 94254 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2043
timestamp 1712078602
transform 1 0 94530 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2045
timestamp 1712078602
transform 1 0 94622 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2057
timestamp 1712078602
transform 1 0 95174 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2069
timestamp 1712078602
transform 1 0 95726 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2081
timestamp 1712078602
transform 1 0 96278 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2093
timestamp 1712078602
transform 1 0 96830 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2099
timestamp 1712078602
transform 1 0 97106 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2101
timestamp 1712078602
transform 1 0 97198 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2113
timestamp 1712078602
transform 1 0 97750 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2125
timestamp 1712078602
transform 1 0 98302 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2137
timestamp 1712078602
transform 1 0 98854 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2149
timestamp 1712078602
transform 1 0 99406 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2155
timestamp 1712078602
transform 1 0 99682 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2157
timestamp 1712078602
transform 1 0 99774 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2169
timestamp 1712078602
transform 1 0 100326 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2181
timestamp 1712078602
transform 1 0 100878 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2193
timestamp 1712078602
transform 1 0 101430 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2205
timestamp 1712078602
transform 1 0 101982 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2211
timestamp 1712078602
transform 1 0 102258 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2213
timestamp 1712078602
transform 1 0 102350 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2225
timestamp 1712078602
transform 1 0 102902 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2237
timestamp 1712078602
transform 1 0 103454 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2249
timestamp 1712078602
transform 1 0 104006 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2261
timestamp 1712078602
transform 1 0 104558 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2267
timestamp 1712078602
transform 1 0 104834 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2269
timestamp 1712078602
transform 1 0 104926 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2281
timestamp 1712078602
transform 1 0 105478 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2293
timestamp 1712078602
transform 1 0 106030 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2305
timestamp 1712078602
transform 1 0 106582 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2317
timestamp 1712078602
transform 1 0 107134 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2323
timestamp 1712078602
transform 1 0 107410 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2325
timestamp 1712078602
transform 1 0 107502 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2337
timestamp 1712078602
transform 1 0 108054 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2349
timestamp 1712078602
transform 1 0 108606 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2361
timestamp 1712078602
transform 1 0 109158 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2373
timestamp 1712078602
transform 1 0 109710 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2379
timestamp 1712078602
transform 1 0 109986 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2381
timestamp 1712078602
transform 1 0 110078 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2393
timestamp 1712078602
transform 1 0 110630 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2405
timestamp 1712078602
transform 1 0 111182 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2417
timestamp 1712078602
transform 1 0 111734 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2429
timestamp 1712078602
transform 1 0 112286 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2435
timestamp 1712078602
transform 1 0 112562 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2437
timestamp 1712078602
transform 1 0 112654 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2449
timestamp 1712078602
transform 1 0 113206 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2461
timestamp 1712078602
transform 1 0 113758 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2473
timestamp 1712078602
transform 1 0 114310 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2485
timestamp 1712078602
transform 1 0 114862 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2491
timestamp 1712078602
transform 1 0 115138 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2493
timestamp 1712078602
transform 1 0 115230 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2505
timestamp 1712078602
transform 1 0 115782 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2517
timestamp 1712078602
transform 1 0 116334 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2529
timestamp 1712078602
transform 1 0 116886 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2541
timestamp 1712078602
transform 1 0 117438 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2547
timestamp 1712078602
transform 1 0 117714 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2549
timestamp 1712078602
transform 1 0 117806 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2561
timestamp 1712078602
transform 1 0 118358 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2573
timestamp 1712078602
transform 1 0 118910 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2585
timestamp 1712078602
transform 1 0 119462 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2597
timestamp 1712078602
transform 1 0 120014 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2603
timestamp 1712078602
transform 1 0 120290 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2605
timestamp 1712078602
transform 1 0 120382 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2617
timestamp 1712078602
transform 1 0 120934 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2629
timestamp 1712078602
transform 1 0 121486 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2641
timestamp 1712078602
transform 1 0 122038 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2653
timestamp 1712078602
transform 1 0 122590 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2659
timestamp 1712078602
transform 1 0 122866 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2661
timestamp 1712078602
transform 1 0 122958 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2673
timestamp 1712078602
transform 1 0 123510 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2685
timestamp 1712078602
transform 1 0 124062 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2697
timestamp 1712078602
transform 1 0 124614 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2709
timestamp 1712078602
transform 1 0 125166 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2715
timestamp 1712078602
transform 1 0 125442 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2717
timestamp 1712078602
transform 1 0 125534 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2729
timestamp 1712078602
transform 1 0 126086 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2741
timestamp 1712078602
transform 1 0 126638 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2753
timestamp 1712078602
transform 1 0 127190 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2765
timestamp 1712078602
transform 1 0 127742 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2771
timestamp 1712078602
transform 1 0 128018 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2773
timestamp 1712078602
transform 1 0 128110 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2785
timestamp 1712078602
transform 1 0 128662 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2797
timestamp 1712078602
transform 1 0 129214 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2809
timestamp 1712078602
transform 1 0 129766 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2821
timestamp 1712078602
transform 1 0 130318 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2827
timestamp 1712078602
transform 1 0 130594 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2829
timestamp 1712078602
transform 1 0 130686 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2841
timestamp 1712078602
transform 1 0 131238 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2853
timestamp 1712078602
transform 1 0 131790 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2865
timestamp 1712078602
transform 1 0 132342 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2877
timestamp 1712078602
transform 1 0 132894 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2883
timestamp 1712078602
transform 1 0 133170 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2885
timestamp 1712078602
transform 1 0 133262 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2897
timestamp 1712078602
transform 1 0 133814 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2909
timestamp 1712078602
transform 1 0 134366 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2921
timestamp 1712078602
transform 1 0 134918 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2933
timestamp 1712078602
transform 1 0 135470 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2939
timestamp 1712078602
transform 1 0 135746 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2941
timestamp 1712078602
transform 1 0 135838 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2953
timestamp 1712078602
transform 1 0 136390 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2965
timestamp 1712078602
transform 1 0 136942 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2977
timestamp 1712078602
transform 1 0 137494 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_2989
timestamp 1712078602
transform 1 0 138046 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_2995
timestamp 1712078602
transform 1 0 138322 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_2997
timestamp 1712078602
transform 1 0 138414 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3009
timestamp 1712078602
transform 1 0 138966 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3021
timestamp 1712078602
transform 1 0 139518 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3033
timestamp 1712078602
transform 1 0 140070 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_3045
timestamp 1712078602
transform 1 0 140622 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_3051
timestamp 1712078602
transform 1 0 140898 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3053
timestamp 1712078602
transform 1 0 140990 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3065
timestamp 1712078602
transform 1 0 141542 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3077
timestamp 1712078602
transform 1 0 142094 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3089
timestamp 1712078602
transform 1 0 142646 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_3101
timestamp 1712078602
transform 1 0 143198 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_3107
timestamp 1712078602
transform 1 0 143474 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3109
timestamp 1712078602
transform 1 0 143566 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3121
timestamp 1712078602
transform 1 0 144118 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3133
timestamp 1712078602
transform 1 0 144670 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3145
timestamp 1712078602
transform 1 0 145222 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_3157
timestamp 1712078602
transform 1 0 145774 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_3163
timestamp 1712078602
transform 1 0 146050 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3165
timestamp 1712078602
transform 1 0 146142 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3177
timestamp 1712078602
transform 1 0 146694 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3189
timestamp 1712078602
transform 1 0 147246 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3201
timestamp 1712078602
transform 1 0 147798 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_3213
timestamp 1712078602
transform 1 0 148350 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_3219
timestamp 1712078602
transform 1 0 148626 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3221
timestamp 1712078602
transform 1 0 148718 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3233
timestamp 1712078602
transform 1 0 149270 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3245
timestamp 1712078602
transform 1 0 149822 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3257
timestamp 1712078602
transform 1 0 150374 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_8_3269
timestamp 1712078602
transform 1 0 150926 0 1 3264
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_8_3275
timestamp 1712078602
transform 1 0 151202 0 1 3264
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3277
timestamp 1712078602
transform 1 0 151294 0 1 3264
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_8_3289
timestamp 1712078602
transform 1 0 151846 0 1 3264
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_8_3301
timestamp 1712078602
transform 1 0 152398 0 1 3264
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1712078602
transform 1 0 690 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1712078602
transform 1 0 1242 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1712078602
transform 1 0 1794 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1712078602
transform 1 0 2346 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1712078602
transform 1 0 2898 0 -1 3808
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1712078602
transform 1 0 3082 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1712078602
transform 1 0 3174 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1712078602
transform 1 0 3726 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1712078602
transform 1 0 4278 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1712078602
transform 1 0 4830 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1712078602
transform 1 0 5382 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1712078602
transform 1 0 5658 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1712078602
transform 1 0 5750 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1712078602
transform 1 0 6302 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1712078602
transform 1 0 6854 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1712078602
transform 1 0 7406 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1712078602
transform 1 0 7958 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1712078602
transform 1 0 8234 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1712078602
transform 1 0 8326 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1712078602
transform 1 0 8878 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1712078602
transform 1 0 9430 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1712078602
transform 1 0 9982 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1712078602
transform 1 0 10534 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1712078602
transform 1 0 10810 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1712078602
transform 1 0 10902 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1712078602
transform 1 0 11454 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1712078602
transform 1 0 12006 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1712078602
transform 1 0 12558 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1712078602
transform 1 0 13110 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1712078602
transform 1 0 13386 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1712078602
transform 1 0 13478 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1712078602
transform 1 0 14030 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1712078602
transform 1 0 14582 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1712078602
transform 1 0 15134 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1712078602
transform 1 0 15686 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1712078602
transform 1 0 15962 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1712078602
transform 1 0 16054 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1712078602
transform 1 0 16606 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1712078602
transform 1 0 17158 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1712078602
transform 1 0 17710 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1712078602
transform 1 0 18262 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1712078602
transform 1 0 18538 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1712078602
transform 1 0 18630 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1712078602
transform 1 0 19182 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1712078602
transform 1 0 19734 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1712078602
transform 1 0 20286 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1712078602
transform 1 0 20838 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1712078602
transform 1 0 21114 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1712078602
transform 1 0 21206 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1712078602
transform 1 0 21758 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1712078602
transform 1 0 22310 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1712078602
transform 1 0 22862 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1712078602
transform 1 0 23414 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1712078602
transform 1 0 23690 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1712078602
transform 1 0 23782 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1712078602
transform 1 0 24334 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1712078602
transform 1 0 24886 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1712078602
transform 1 0 25438 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1712078602
transform 1 0 25990 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1712078602
transform 1 0 26266 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1712078602
transform 1 0 26358 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1712078602
transform 1 0 26910 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1712078602
transform 1 0 27462 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1712078602
transform 1 0 28014 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1712078602
transform 1 0 28566 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1712078602
transform 1 0 28842 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1712078602
transform 1 0 28934 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1712078602
transform 1 0 29486 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1712078602
transform 1 0 30038 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1712078602
transform 1 0 30590 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1712078602
transform 1 0 31142 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1712078602
transform 1 0 31418 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1712078602
transform 1 0 31510 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1712078602
transform 1 0 32062 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1712078602
transform 1 0 32614 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1712078602
transform 1 0 33166 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1712078602
transform 1 0 33718 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1712078602
transform 1 0 33994 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1712078602
transform 1 0 34086 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1712078602
transform 1 0 34638 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1712078602
transform 1 0 35190 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1712078602
transform 1 0 35742 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1712078602
transform 1 0 36294 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1712078602
transform 1 0 36570 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1712078602
transform 1 0 36662 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1712078602
transform 1 0 37214 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1712078602
transform 1 0 37766 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1712078602
transform 1 0 38318 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1712078602
transform 1 0 38870 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1712078602
transform 1 0 39146 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1712078602
transform 1 0 39238 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1712078602
transform 1 0 39790 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_865
timestamp 1712078602
transform 1 0 40342 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1712078602
transform 1 0 40894 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1712078602
transform 1 0 41446 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1712078602
transform 1 0 41722 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1712078602
transform 1 0 41814 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1712078602
transform 1 0 42366 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_921
timestamp 1712078602
transform 1 0 42918 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_933
timestamp 1712078602
transform 1 0 43470 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_945
timestamp 1712078602
transform 1 0 44022 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_951
timestamp 1712078602
transform 1 0 44298 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1712078602
transform 1 0 44390 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1712078602
transform 1 0 44942 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_977
timestamp 1712078602
transform 1 0 45494 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_989
timestamp 1712078602
transform 1 0 46046 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1001
timestamp 1712078602
transform 1 0 46598 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1007
timestamp 1712078602
transform 1 0 46874 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1712078602
transform 1 0 46966 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1712078602
transform 1 0 47518 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1033
timestamp 1712078602
transform 1 0 48070 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1045
timestamp 1712078602
transform 1 0 48622 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1057
timestamp 1712078602
transform 1 0 49174 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1712078602
transform 1 0 49450 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1712078602
transform 1 0 49542 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1712078602
transform 1 0 50094 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1089
timestamp 1712078602
transform 1 0 50646 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1101
timestamp 1712078602
transform 1 0 51198 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1712078602
transform 1 0 51750 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1712078602
transform 1 0 52026 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1712078602
transform 1 0 52118 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1712078602
transform 1 0 52670 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1145
timestamp 1712078602
transform 1 0 53222 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1157
timestamp 1712078602
transform 1 0 53774 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1712078602
transform 1 0 54326 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1712078602
transform 1 0 54602 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1712078602
transform 1 0 54694 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1712078602
transform 1 0 55246 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1201
timestamp 1712078602
transform 1 0 55798 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1213
timestamp 1712078602
transform 1 0 56350 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1225
timestamp 1712078602
transform 1 0 56902 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1231
timestamp 1712078602
transform 1 0 57178 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1712078602
transform 1 0 57270 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1712078602
transform 1 0 57822 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1257
timestamp 1712078602
transform 1 0 58374 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1269
timestamp 1712078602
transform 1 0 58926 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1281
timestamp 1712078602
transform 1 0 59478 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1287
timestamp 1712078602
transform 1 0 59754 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1289
timestamp 1712078602
transform 1 0 59846 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1301
timestamp 1712078602
transform 1 0 60398 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1313
timestamp 1712078602
transform 1 0 60950 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1325
timestamp 1712078602
transform 1 0 61502 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1337
timestamp 1712078602
transform 1 0 62054 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1343
timestamp 1712078602
transform 1 0 62330 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1345
timestamp 1712078602
transform 1 0 62422 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1357
timestamp 1712078602
transform 1 0 62974 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1369
timestamp 1712078602
transform 1 0 63526 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1381
timestamp 1712078602
transform 1 0 64078 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1393
timestamp 1712078602
transform 1 0 64630 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1399
timestamp 1712078602
transform 1 0 64906 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1712078602
transform 1 0 64998 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1712078602
transform 1 0 65550 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1425
timestamp 1712078602
transform 1 0 66102 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1437
timestamp 1712078602
transform 1 0 66654 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1449
timestamp 1712078602
transform 1 0 67206 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1455
timestamp 1712078602
transform 1 0 67482 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1712078602
transform 1 0 67574 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1712078602
transform 1 0 68126 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1481
timestamp 1712078602
transform 1 0 68678 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1493
timestamp 1712078602
transform 1 0 69230 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1505
timestamp 1712078602
transform 1 0 69782 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1511
timestamp 1712078602
transform 1 0 70058 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1712078602
transform 1 0 70150 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1712078602
transform 1 0 70702 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1537
timestamp 1712078602
transform 1 0 71254 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1549
timestamp 1712078602
transform 1 0 71806 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1561
timestamp 1712078602
transform 1 0 72358 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1567
timestamp 1712078602
transform 1 0 72634 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1712078602
transform 1 0 72726 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1712078602
transform 1 0 73278 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1593
timestamp 1712078602
transform 1 0 73830 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1605
timestamp 1712078602
transform 1 0 74382 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1617
timestamp 1712078602
transform 1 0 74934 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1623
timestamp 1712078602
transform 1 0 75210 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1625
timestamp 1712078602
transform 1 0 75302 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1637
timestamp 1712078602
transform 1 0 75854 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1649
timestamp 1712078602
transform 1 0 76406 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1661
timestamp 1712078602
transform 1 0 76958 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1673
timestamp 1712078602
transform 1 0 77510 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1679
timestamp 1712078602
transform 1 0 77786 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1681
timestamp 1712078602
transform 1 0 77878 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1693
timestamp 1712078602
transform 1 0 78430 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1705
timestamp 1712078602
transform 1 0 78982 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1717
timestamp 1712078602
transform 1 0 79534 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1729
timestamp 1712078602
transform 1 0 80086 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1735
timestamp 1712078602
transform 1 0 80362 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1737
timestamp 1712078602
transform 1 0 80454 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1749
timestamp 1712078602
transform 1 0 81006 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1761
timestamp 1712078602
transform 1 0 81558 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1773
timestamp 1712078602
transform 1 0 82110 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1785
timestamp 1712078602
transform 1 0 82662 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1791
timestamp 1712078602
transform 1 0 82938 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1793
timestamp 1712078602
transform 1 0 83030 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1805
timestamp 1712078602
transform 1 0 83582 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1817
timestamp 1712078602
transform 1 0 84134 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1829
timestamp 1712078602
transform 1 0 84686 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1841
timestamp 1712078602
transform 1 0 85238 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1847
timestamp 1712078602
transform 1 0 85514 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1849
timestamp 1712078602
transform 1 0 85606 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1861
timestamp 1712078602
transform 1 0 86158 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1873
timestamp 1712078602
transform 1 0 86710 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1885
timestamp 1712078602
transform 1 0 87262 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1897
timestamp 1712078602
transform 1 0 87814 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1903
timestamp 1712078602
transform 1 0 88090 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1905
timestamp 1712078602
transform 1 0 88182 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1917
timestamp 1712078602
transform 1 0 88734 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1929
timestamp 1712078602
transform 1 0 89286 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1941
timestamp 1712078602
transform 1 0 89838 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_1953
timestamp 1712078602
transform 1 0 90390 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_1959
timestamp 1712078602
transform 1 0 90666 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1961
timestamp 1712078602
transform 1 0 90758 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1973
timestamp 1712078602
transform 1 0 91310 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1985
timestamp 1712078602
transform 1 0 91862 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_1997
timestamp 1712078602
transform 1 0 92414 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2009
timestamp 1712078602
transform 1 0 92966 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2015
timestamp 1712078602
transform 1 0 93242 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2017
timestamp 1712078602
transform 1 0 93334 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2029
timestamp 1712078602
transform 1 0 93886 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2041
timestamp 1712078602
transform 1 0 94438 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2053
timestamp 1712078602
transform 1 0 94990 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2065
timestamp 1712078602
transform 1 0 95542 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2071
timestamp 1712078602
transform 1 0 95818 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2073
timestamp 1712078602
transform 1 0 95910 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2085
timestamp 1712078602
transform 1 0 96462 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2097
timestamp 1712078602
transform 1 0 97014 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2109
timestamp 1712078602
transform 1 0 97566 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2121
timestamp 1712078602
transform 1 0 98118 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2127
timestamp 1712078602
transform 1 0 98394 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2129
timestamp 1712078602
transform 1 0 98486 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2141
timestamp 1712078602
transform 1 0 99038 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2153
timestamp 1712078602
transform 1 0 99590 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2165
timestamp 1712078602
transform 1 0 100142 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2177
timestamp 1712078602
transform 1 0 100694 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2183
timestamp 1712078602
transform 1 0 100970 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2185
timestamp 1712078602
transform 1 0 101062 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2197
timestamp 1712078602
transform 1 0 101614 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2209
timestamp 1712078602
transform 1 0 102166 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2221
timestamp 1712078602
transform 1 0 102718 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2233
timestamp 1712078602
transform 1 0 103270 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2239
timestamp 1712078602
transform 1 0 103546 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2241
timestamp 1712078602
transform 1 0 103638 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2253
timestamp 1712078602
transform 1 0 104190 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2265
timestamp 1712078602
transform 1 0 104742 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2277
timestamp 1712078602
transform 1 0 105294 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2289
timestamp 1712078602
transform 1 0 105846 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2295
timestamp 1712078602
transform 1 0 106122 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2297
timestamp 1712078602
transform 1 0 106214 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2309
timestamp 1712078602
transform 1 0 106766 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2321
timestamp 1712078602
transform 1 0 107318 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2333
timestamp 1712078602
transform 1 0 107870 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2345
timestamp 1712078602
transform 1 0 108422 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2351
timestamp 1712078602
transform 1 0 108698 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2353
timestamp 1712078602
transform 1 0 108790 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2365
timestamp 1712078602
transform 1 0 109342 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2377
timestamp 1712078602
transform 1 0 109894 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2389
timestamp 1712078602
transform 1 0 110446 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2401
timestamp 1712078602
transform 1 0 110998 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2407
timestamp 1712078602
transform 1 0 111274 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2409
timestamp 1712078602
transform 1 0 111366 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2421
timestamp 1712078602
transform 1 0 111918 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2433
timestamp 1712078602
transform 1 0 112470 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2445
timestamp 1712078602
transform 1 0 113022 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2457
timestamp 1712078602
transform 1 0 113574 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2463
timestamp 1712078602
transform 1 0 113850 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2465
timestamp 1712078602
transform 1 0 113942 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2477
timestamp 1712078602
transform 1 0 114494 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2489
timestamp 1712078602
transform 1 0 115046 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2501
timestamp 1712078602
transform 1 0 115598 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2513
timestamp 1712078602
transform 1 0 116150 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2519
timestamp 1712078602
transform 1 0 116426 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2521
timestamp 1712078602
transform 1 0 116518 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2533
timestamp 1712078602
transform 1 0 117070 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2545
timestamp 1712078602
transform 1 0 117622 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2557
timestamp 1712078602
transform 1 0 118174 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2569
timestamp 1712078602
transform 1 0 118726 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2575
timestamp 1712078602
transform 1 0 119002 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2577
timestamp 1712078602
transform 1 0 119094 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2589
timestamp 1712078602
transform 1 0 119646 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2601
timestamp 1712078602
transform 1 0 120198 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2613
timestamp 1712078602
transform 1 0 120750 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2625
timestamp 1712078602
transform 1 0 121302 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2631
timestamp 1712078602
transform 1 0 121578 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2633
timestamp 1712078602
transform 1 0 121670 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2645
timestamp 1712078602
transform 1 0 122222 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2657
timestamp 1712078602
transform 1 0 122774 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2669
timestamp 1712078602
transform 1 0 123326 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2681
timestamp 1712078602
transform 1 0 123878 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2687
timestamp 1712078602
transform 1 0 124154 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2689
timestamp 1712078602
transform 1 0 124246 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2701
timestamp 1712078602
transform 1 0 124798 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2713
timestamp 1712078602
transform 1 0 125350 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2725
timestamp 1712078602
transform 1 0 125902 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2737
timestamp 1712078602
transform 1 0 126454 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2743
timestamp 1712078602
transform 1 0 126730 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2745
timestamp 1712078602
transform 1 0 126822 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2757
timestamp 1712078602
transform 1 0 127374 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2769
timestamp 1712078602
transform 1 0 127926 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2781
timestamp 1712078602
transform 1 0 128478 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2793
timestamp 1712078602
transform 1 0 129030 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2799
timestamp 1712078602
transform 1 0 129306 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2801
timestamp 1712078602
transform 1 0 129398 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2813
timestamp 1712078602
transform 1 0 129950 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2825
timestamp 1712078602
transform 1 0 130502 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2837
timestamp 1712078602
transform 1 0 131054 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2849
timestamp 1712078602
transform 1 0 131606 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2855
timestamp 1712078602
transform 1 0 131882 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2857
timestamp 1712078602
transform 1 0 131974 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2869
timestamp 1712078602
transform 1 0 132526 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2881
timestamp 1712078602
transform 1 0 133078 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2893
timestamp 1712078602
transform 1 0 133630 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2905
timestamp 1712078602
transform 1 0 134182 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2911
timestamp 1712078602
transform 1 0 134458 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2913
timestamp 1712078602
transform 1 0 134550 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2925
timestamp 1712078602
transform 1 0 135102 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2937
timestamp 1712078602
transform 1 0 135654 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2949
timestamp 1712078602
transform 1 0 136206 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_2961
timestamp 1712078602
transform 1 0 136758 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_2967
timestamp 1712078602
transform 1 0 137034 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2969
timestamp 1712078602
transform 1 0 137126 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2981
timestamp 1712078602
transform 1 0 137678 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_2993
timestamp 1712078602
transform 1 0 138230 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3005
timestamp 1712078602
transform 1 0 138782 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_3017
timestamp 1712078602
transform 1 0 139334 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_3023
timestamp 1712078602
transform 1 0 139610 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3025
timestamp 1712078602
transform 1 0 139702 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3037
timestamp 1712078602
transform 1 0 140254 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3049
timestamp 1712078602
transform 1 0 140806 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3061
timestamp 1712078602
transform 1 0 141358 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_3073
timestamp 1712078602
transform 1 0 141910 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_3079
timestamp 1712078602
transform 1 0 142186 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3081
timestamp 1712078602
transform 1 0 142278 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3093
timestamp 1712078602
transform 1 0 142830 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3105
timestamp 1712078602
transform 1 0 143382 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3117
timestamp 1712078602
transform 1 0 143934 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_3129
timestamp 1712078602
transform 1 0 144486 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_3135
timestamp 1712078602
transform 1 0 144762 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3137
timestamp 1712078602
transform 1 0 144854 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3149
timestamp 1712078602
transform 1 0 145406 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3161
timestamp 1712078602
transform 1 0 145958 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3173
timestamp 1712078602
transform 1 0 146510 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_3185
timestamp 1712078602
transform 1 0 147062 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_3191
timestamp 1712078602
transform 1 0 147338 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3193
timestamp 1712078602
transform 1 0 147430 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3205
timestamp 1712078602
transform 1 0 147982 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3217
timestamp 1712078602
transform 1 0 148534 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3229
timestamp 1712078602
transform 1 0 149086 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_3241
timestamp 1712078602
transform 1 0 149638 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_3247
timestamp 1712078602
transform 1 0 149914 0 -1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3249
timestamp 1712078602
transform 1 0 150006 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3261
timestamp 1712078602
transform 1 0 150558 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3273
timestamp 1712078602
transform 1 0 151110 0 -1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_9_3285
timestamp 1712078602
transform 1 0 151662 0 -1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_9_3297
timestamp 1712078602
transform 1 0 152214 0 -1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_9_3303
timestamp 1712078602
transform 1 0 152490 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_9_3305
timestamp 1712078602
transform 1 0 152582 0 -1 3808
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1712078602
transform 1 0 690 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1712078602
transform 1 0 1242 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1712078602
transform 1 0 1794 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1712078602
transform 1 0 1886 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1712078602
transform 1 0 2438 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1712078602
transform 1 0 2990 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1712078602
transform 1 0 3542 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1712078602
transform 1 0 4094 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1712078602
transform 1 0 4370 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1712078602
transform 1 0 4462 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1712078602
transform 1 0 5014 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1712078602
transform 1 0 5566 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1712078602
transform 1 0 6118 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1712078602
transform 1 0 6670 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1712078602
transform 1 0 6946 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1712078602
transform 1 0 7038 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1712078602
transform 1 0 7590 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1712078602
transform 1 0 8142 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1712078602
transform 1 0 8694 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1712078602
transform 1 0 9246 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1712078602
transform 1 0 9522 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1712078602
transform 1 0 9614 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1712078602
transform 1 0 10166 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1712078602
transform 1 0 10718 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1712078602
transform 1 0 11270 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1712078602
transform 1 0 11822 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1712078602
transform 1 0 12098 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1712078602
transform 1 0 12190 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1712078602
transform 1 0 12742 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1712078602
transform 1 0 13294 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1712078602
transform 1 0 13846 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1712078602
transform 1 0 14398 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1712078602
transform 1 0 14674 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1712078602
transform 1 0 14766 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1712078602
transform 1 0 15318 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1712078602
transform 1 0 15870 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1712078602
transform 1 0 16422 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1712078602
transform 1 0 16974 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1712078602
transform 1 0 17250 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1712078602
transform 1 0 17342 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1712078602
transform 1 0 17894 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1712078602
transform 1 0 18446 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1712078602
transform 1 0 18998 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1712078602
transform 1 0 19550 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1712078602
transform 1 0 19826 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1712078602
transform 1 0 19918 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1712078602
transform 1 0 20470 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1712078602
transform 1 0 21022 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1712078602
transform 1 0 21574 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1712078602
transform 1 0 22126 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1712078602
transform 1 0 22402 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1712078602
transform 1 0 22494 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1712078602
transform 1 0 23046 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1712078602
transform 1 0 23598 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1712078602
transform 1 0 24150 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1712078602
transform 1 0 24702 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1712078602
transform 1 0 24978 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1712078602
transform 1 0 25070 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1712078602
transform 1 0 25622 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1712078602
transform 1 0 26174 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1712078602
transform 1 0 26726 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1712078602
transform 1 0 27278 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1712078602
transform 1 0 27554 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1712078602
transform 1 0 27646 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1712078602
transform 1 0 28198 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1712078602
transform 1 0 28750 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1712078602
transform 1 0 29302 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1712078602
transform 1 0 29854 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1712078602
transform 1 0 30130 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1712078602
transform 1 0 30222 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1712078602
transform 1 0 30774 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1712078602
transform 1 0 31326 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1712078602
transform 1 0 31878 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1712078602
transform 1 0 32430 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1712078602
transform 1 0 32706 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1712078602
transform 1 0 32798 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1712078602
transform 1 0 33350 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1712078602
transform 1 0 33902 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1712078602
transform 1 0 34454 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1712078602
transform 1 0 35006 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1712078602
transform 1 0 35282 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1712078602
transform 1 0 35374 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1712078602
transform 1 0 35926 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1712078602
transform 1 0 36478 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1712078602
transform 1 0 37030 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1712078602
transform 1 0 37582 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1712078602
transform 1 0 37858 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_813
timestamp 1712078602
transform 1 0 37950 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_825
timestamp 1712078602
transform 1 0 38502 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_837
timestamp 1712078602
transform 1 0 39054 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_849
timestamp 1712078602
transform 1 0 39606 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1712078602
transform 1 0 40158 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1712078602
transform 1 0 40434 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_869
timestamp 1712078602
transform 1 0 40526 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_881
timestamp 1712078602
transform 1 0 41078 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_893
timestamp 1712078602
transform 1 0 41630 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_905
timestamp 1712078602
transform 1 0 42182 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1712078602
transform 1 0 42734 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1712078602
transform 1 0 43010 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_925
timestamp 1712078602
transform 1 0 43102 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_937
timestamp 1712078602
transform 1 0 43654 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_949
timestamp 1712078602
transform 1 0 44206 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_961
timestamp 1712078602
transform 1 0 44758 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1712078602
transform 1 0 45310 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1712078602
transform 1 0 45586 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_981
timestamp 1712078602
transform 1 0 45678 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_993
timestamp 1712078602
transform 1 0 46230 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1005
timestamp 1712078602
transform 1 0 46782 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1017
timestamp 1712078602
transform 1 0 47334 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1029
timestamp 1712078602
transform 1 0 47886 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1035
timestamp 1712078602
transform 1 0 48162 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1037
timestamp 1712078602
transform 1 0 48254 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1049
timestamp 1712078602
transform 1 0 48806 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1061
timestamp 1712078602
transform 1 0 49358 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1073
timestamp 1712078602
transform 1 0 49910 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1085
timestamp 1712078602
transform 1 0 50462 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1712078602
transform 1 0 50738 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1093
timestamp 1712078602
transform 1 0 50830 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1105
timestamp 1712078602
transform 1 0 51382 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1117
timestamp 1712078602
transform 1 0 51934 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1129
timestamp 1712078602
transform 1 0 52486 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1712078602
transform 1 0 53038 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1712078602
transform 1 0 53314 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1149
timestamp 1712078602
transform 1 0 53406 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1161
timestamp 1712078602
transform 1 0 53958 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1173
timestamp 1712078602
transform 1 0 54510 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1185
timestamp 1712078602
transform 1 0 55062 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1712078602
transform 1 0 55614 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1712078602
transform 1 0 55890 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1205
timestamp 1712078602
transform 1 0 55982 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1217
timestamp 1712078602
transform 1 0 56534 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1229
timestamp 1712078602
transform 1 0 57086 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1241
timestamp 1712078602
transform 1 0 57638 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1253
timestamp 1712078602
transform 1 0 58190 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1259
timestamp 1712078602
transform 1 0 58466 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1261
timestamp 1712078602
transform 1 0 58558 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1273
timestamp 1712078602
transform 1 0 59110 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1285
timestamp 1712078602
transform 1 0 59662 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1297
timestamp 1712078602
transform 1 0 60214 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1309
timestamp 1712078602
transform 1 0 60766 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1315
timestamp 1712078602
transform 1 0 61042 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1317
timestamp 1712078602
transform 1 0 61134 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1329
timestamp 1712078602
transform 1 0 61686 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1341
timestamp 1712078602
transform 1 0 62238 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1353
timestamp 1712078602
transform 1 0 62790 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1365
timestamp 1712078602
transform 1 0 63342 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1371
timestamp 1712078602
transform 1 0 63618 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1373
timestamp 1712078602
transform 1 0 63710 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1385
timestamp 1712078602
transform 1 0 64262 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1397
timestamp 1712078602
transform 1 0 64814 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1409
timestamp 1712078602
transform 1 0 65366 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1421
timestamp 1712078602
transform 1 0 65918 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1427
timestamp 1712078602
transform 1 0 66194 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1429
timestamp 1712078602
transform 1 0 66286 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1441
timestamp 1712078602
transform 1 0 66838 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1453
timestamp 1712078602
transform 1 0 67390 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1465
timestamp 1712078602
transform 1 0 67942 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1477
timestamp 1712078602
transform 1 0 68494 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1483
timestamp 1712078602
transform 1 0 68770 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1485
timestamp 1712078602
transform 1 0 68862 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1497
timestamp 1712078602
transform 1 0 69414 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1509
timestamp 1712078602
transform 1 0 69966 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1521
timestamp 1712078602
transform 1 0 70518 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1533
timestamp 1712078602
transform 1 0 71070 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1539
timestamp 1712078602
transform 1 0 71346 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1541
timestamp 1712078602
transform 1 0 71438 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1553
timestamp 1712078602
transform 1 0 71990 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1565
timestamp 1712078602
transform 1 0 72542 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1577
timestamp 1712078602
transform 1 0 73094 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1589
timestamp 1712078602
transform 1 0 73646 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1595
timestamp 1712078602
transform 1 0 73922 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1597
timestamp 1712078602
transform 1 0 74014 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1609
timestamp 1712078602
transform 1 0 74566 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1621
timestamp 1712078602
transform 1 0 75118 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1633
timestamp 1712078602
transform 1 0 75670 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1645
timestamp 1712078602
transform 1 0 76222 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1651
timestamp 1712078602
transform 1 0 76498 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1653
timestamp 1712078602
transform 1 0 76590 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1665
timestamp 1712078602
transform 1 0 77142 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1677
timestamp 1712078602
transform 1 0 77694 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1689
timestamp 1712078602
transform 1 0 78246 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1701
timestamp 1712078602
transform 1 0 78798 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1707
timestamp 1712078602
transform 1 0 79074 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1709
timestamp 1712078602
transform 1 0 79166 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1721
timestamp 1712078602
transform 1 0 79718 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1733
timestamp 1712078602
transform 1 0 80270 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1745
timestamp 1712078602
transform 1 0 80822 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1757
timestamp 1712078602
transform 1 0 81374 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1763
timestamp 1712078602
transform 1 0 81650 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1765
timestamp 1712078602
transform 1 0 81742 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1777
timestamp 1712078602
transform 1 0 82294 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1789
timestamp 1712078602
transform 1 0 82846 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1801
timestamp 1712078602
transform 1 0 83398 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1813
timestamp 1712078602
transform 1 0 83950 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1819
timestamp 1712078602
transform 1 0 84226 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1821
timestamp 1712078602
transform 1 0 84318 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1833
timestamp 1712078602
transform 1 0 84870 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1845
timestamp 1712078602
transform 1 0 85422 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1857
timestamp 1712078602
transform 1 0 85974 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1869
timestamp 1712078602
transform 1 0 86526 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1875
timestamp 1712078602
transform 1 0 86802 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1877
timestamp 1712078602
transform 1 0 86894 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1889
timestamp 1712078602
transform 1 0 87446 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1901
timestamp 1712078602
transform 1 0 87998 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1913
timestamp 1712078602
transform 1 0 88550 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1925
timestamp 1712078602
transform 1 0 89102 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1931
timestamp 1712078602
transform 1 0 89378 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1933
timestamp 1712078602
transform 1 0 89470 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1945
timestamp 1712078602
transform 1 0 90022 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1957
timestamp 1712078602
transform 1 0 90574 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1969
timestamp 1712078602
transform 1 0 91126 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_1981
timestamp 1712078602
transform 1 0 91678 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_1987
timestamp 1712078602
transform 1 0 91954 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_1989
timestamp 1712078602
transform 1 0 92046 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2001
timestamp 1712078602
transform 1 0 92598 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2013
timestamp 1712078602
transform 1 0 93150 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2025
timestamp 1712078602
transform 1 0 93702 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2037
timestamp 1712078602
transform 1 0 94254 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2043
timestamp 1712078602
transform 1 0 94530 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2045
timestamp 1712078602
transform 1 0 94622 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2057
timestamp 1712078602
transform 1 0 95174 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2069
timestamp 1712078602
transform 1 0 95726 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2081
timestamp 1712078602
transform 1 0 96278 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2093
timestamp 1712078602
transform 1 0 96830 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2099
timestamp 1712078602
transform 1 0 97106 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2101
timestamp 1712078602
transform 1 0 97198 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2113
timestamp 1712078602
transform 1 0 97750 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2125
timestamp 1712078602
transform 1 0 98302 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2137
timestamp 1712078602
transform 1 0 98854 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2149
timestamp 1712078602
transform 1 0 99406 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2155
timestamp 1712078602
transform 1 0 99682 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2157
timestamp 1712078602
transform 1 0 99774 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2169
timestamp 1712078602
transform 1 0 100326 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2181
timestamp 1712078602
transform 1 0 100878 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2193
timestamp 1712078602
transform 1 0 101430 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2205
timestamp 1712078602
transform 1 0 101982 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2211
timestamp 1712078602
transform 1 0 102258 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2213
timestamp 1712078602
transform 1 0 102350 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2225
timestamp 1712078602
transform 1 0 102902 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2237
timestamp 1712078602
transform 1 0 103454 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2249
timestamp 1712078602
transform 1 0 104006 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2261
timestamp 1712078602
transform 1 0 104558 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2267
timestamp 1712078602
transform 1 0 104834 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2269
timestamp 1712078602
transform 1 0 104926 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2281
timestamp 1712078602
transform 1 0 105478 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2293
timestamp 1712078602
transform 1 0 106030 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2305
timestamp 1712078602
transform 1 0 106582 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2317
timestamp 1712078602
transform 1 0 107134 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2323
timestamp 1712078602
transform 1 0 107410 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2325
timestamp 1712078602
transform 1 0 107502 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2337
timestamp 1712078602
transform 1 0 108054 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2349
timestamp 1712078602
transform 1 0 108606 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2361
timestamp 1712078602
transform 1 0 109158 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2373
timestamp 1712078602
transform 1 0 109710 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2379
timestamp 1712078602
transform 1 0 109986 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2381
timestamp 1712078602
transform 1 0 110078 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2393
timestamp 1712078602
transform 1 0 110630 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2405
timestamp 1712078602
transform 1 0 111182 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2417
timestamp 1712078602
transform 1 0 111734 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2429
timestamp 1712078602
transform 1 0 112286 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2435
timestamp 1712078602
transform 1 0 112562 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2437
timestamp 1712078602
transform 1 0 112654 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2449
timestamp 1712078602
transform 1 0 113206 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2461
timestamp 1712078602
transform 1 0 113758 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2473
timestamp 1712078602
transform 1 0 114310 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2485
timestamp 1712078602
transform 1 0 114862 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2491
timestamp 1712078602
transform 1 0 115138 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2493
timestamp 1712078602
transform 1 0 115230 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2505
timestamp 1712078602
transform 1 0 115782 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2517
timestamp 1712078602
transform 1 0 116334 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2529
timestamp 1712078602
transform 1 0 116886 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2541
timestamp 1712078602
transform 1 0 117438 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2547
timestamp 1712078602
transform 1 0 117714 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2549
timestamp 1712078602
transform 1 0 117806 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2561
timestamp 1712078602
transform 1 0 118358 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2573
timestamp 1712078602
transform 1 0 118910 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2585
timestamp 1712078602
transform 1 0 119462 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2597
timestamp 1712078602
transform 1 0 120014 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2603
timestamp 1712078602
transform 1 0 120290 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2605
timestamp 1712078602
transform 1 0 120382 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2617
timestamp 1712078602
transform 1 0 120934 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2629
timestamp 1712078602
transform 1 0 121486 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2641
timestamp 1712078602
transform 1 0 122038 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2653
timestamp 1712078602
transform 1 0 122590 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2659
timestamp 1712078602
transform 1 0 122866 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2661
timestamp 1712078602
transform 1 0 122958 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2673
timestamp 1712078602
transform 1 0 123510 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2685
timestamp 1712078602
transform 1 0 124062 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2697
timestamp 1712078602
transform 1 0 124614 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2709
timestamp 1712078602
transform 1 0 125166 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2715
timestamp 1712078602
transform 1 0 125442 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2717
timestamp 1712078602
transform 1 0 125534 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2729
timestamp 1712078602
transform 1 0 126086 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2741
timestamp 1712078602
transform 1 0 126638 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2753
timestamp 1712078602
transform 1 0 127190 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2765
timestamp 1712078602
transform 1 0 127742 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2771
timestamp 1712078602
transform 1 0 128018 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2773
timestamp 1712078602
transform 1 0 128110 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2785
timestamp 1712078602
transform 1 0 128662 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2797
timestamp 1712078602
transform 1 0 129214 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2809
timestamp 1712078602
transform 1 0 129766 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2821
timestamp 1712078602
transform 1 0 130318 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2827
timestamp 1712078602
transform 1 0 130594 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2829
timestamp 1712078602
transform 1 0 130686 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2841
timestamp 1712078602
transform 1 0 131238 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2853
timestamp 1712078602
transform 1 0 131790 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2865
timestamp 1712078602
transform 1 0 132342 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2877
timestamp 1712078602
transform 1 0 132894 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2883
timestamp 1712078602
transform 1 0 133170 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2885
timestamp 1712078602
transform 1 0 133262 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2897
timestamp 1712078602
transform 1 0 133814 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2909
timestamp 1712078602
transform 1 0 134366 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2921
timestamp 1712078602
transform 1 0 134918 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2933
timestamp 1712078602
transform 1 0 135470 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2939
timestamp 1712078602
transform 1 0 135746 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2941
timestamp 1712078602
transform 1 0 135838 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2953
timestamp 1712078602
transform 1 0 136390 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2965
timestamp 1712078602
transform 1 0 136942 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2977
timestamp 1712078602
transform 1 0 137494 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_2989
timestamp 1712078602
transform 1 0 138046 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_2995
timestamp 1712078602
transform 1 0 138322 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_2997
timestamp 1712078602
transform 1 0 138414 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3009
timestamp 1712078602
transform 1 0 138966 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3021
timestamp 1712078602
transform 1 0 139518 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3033
timestamp 1712078602
transform 1 0 140070 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_3045
timestamp 1712078602
transform 1 0 140622 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_3051
timestamp 1712078602
transform 1 0 140898 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3053
timestamp 1712078602
transform 1 0 140990 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3065
timestamp 1712078602
transform 1 0 141542 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3077
timestamp 1712078602
transform 1 0 142094 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3089
timestamp 1712078602
transform 1 0 142646 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_3101
timestamp 1712078602
transform 1 0 143198 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_3107
timestamp 1712078602
transform 1 0 143474 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3109
timestamp 1712078602
transform 1 0 143566 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3121
timestamp 1712078602
transform 1 0 144118 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3133
timestamp 1712078602
transform 1 0 144670 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3145
timestamp 1712078602
transform 1 0 145222 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_3157
timestamp 1712078602
transform 1 0 145774 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_3163
timestamp 1712078602
transform 1 0 146050 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3165
timestamp 1712078602
transform 1 0 146142 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3177
timestamp 1712078602
transform 1 0 146694 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3189
timestamp 1712078602
transform 1 0 147246 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3201
timestamp 1712078602
transform 1 0 147798 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_3213
timestamp 1712078602
transform 1 0 148350 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_3219
timestamp 1712078602
transform 1 0 148626 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3221
timestamp 1712078602
transform 1 0 148718 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3233
timestamp 1712078602
transform 1 0 149270 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3245
timestamp 1712078602
transform 1 0 149822 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3257
timestamp 1712078602
transform 1 0 150374 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_10_3269
timestamp 1712078602
transform 1 0 150926 0 1 3808
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_10_3275
timestamp 1712078602
transform 1 0 151202 0 1 3808
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3277
timestamp 1712078602
transform 1 0 151294 0 1 3808
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_10_3289
timestamp 1712078602
transform 1 0 151846 0 1 3808
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_10_3301
timestamp 1712078602
transform 1 0 152398 0 1 3808
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_11_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 828 0 -1 4352
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_11_10
timestamp 1712078602
transform 1 0 1012 0 -1 4352
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_11_14
timestamp 1712078602
transform 1 0 1196 0 -1 4352
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp 1712078602
transform 1 0 1380 0 -1 4352
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_11_22
timestamp 1712078602
transform 1 0 1564 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1712078602
transform 1 0 2116 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1712078602
transform 1 0 2668 0 -1 4352
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1712078602
transform 1 0 3036 0 -1 4352
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1712078602
transform 1 0 3174 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1712078602
transform 1 0 3726 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1712078602
transform 1 0 4278 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1712078602
transform 1 0 4830 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1712078602
transform 1 0 5382 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1712078602
transform 1 0 5658 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1712078602
transform 1 0 5750 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1712078602
transform 1 0 6302 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1712078602
transform 1 0 6854 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1712078602
transform 1 0 7406 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1712078602
transform 1 0 7958 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1712078602
transform 1 0 8234 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1712078602
transform 1 0 8326 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1712078602
transform 1 0 8878 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1712078602
transform 1 0 9430 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1712078602
transform 1 0 9982 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1712078602
transform 1 0 10534 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1712078602
transform 1 0 10810 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1712078602
transform 1 0 10902 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1712078602
transform 1 0 11454 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1712078602
transform 1 0 12006 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1712078602
transform 1 0 12558 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1712078602
transform 1 0 13110 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1712078602
transform 1 0 13386 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1712078602
transform 1 0 13478 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1712078602
transform 1 0 14030 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1712078602
transform 1 0 14582 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1712078602
transform 1 0 15134 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1712078602
transform 1 0 15686 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1712078602
transform 1 0 15962 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1712078602
transform 1 0 16054 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1712078602
transform 1 0 16606 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1712078602
transform 1 0 17158 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1712078602
transform 1 0 17710 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1712078602
transform 1 0 18262 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1712078602
transform 1 0 18538 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1712078602
transform 1 0 18630 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1712078602
transform 1 0 19182 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1712078602
transform 1 0 19734 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1712078602
transform 1 0 20286 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1712078602
transform 1 0 20838 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1712078602
transform 1 0 21114 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1712078602
transform 1 0 21206 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1712078602
transform 1 0 21758 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1712078602
transform 1 0 22310 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1712078602
transform 1 0 22862 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1712078602
transform 1 0 23414 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1712078602
transform 1 0 23690 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1712078602
transform 1 0 23782 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1712078602
transform 1 0 24334 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1712078602
transform 1 0 24886 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1712078602
transform 1 0 25438 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1712078602
transform 1 0 25990 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1712078602
transform 1 0 26266 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1712078602
transform 1 0 26358 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1712078602
transform 1 0 26910 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1712078602
transform 1 0 27462 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1712078602
transform 1 0 28014 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1712078602
transform 1 0 28566 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1712078602
transform 1 0 28842 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1712078602
transform 1 0 28934 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1712078602
transform 1 0 29486 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1712078602
transform 1 0 30038 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1712078602
transform 1 0 30590 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1712078602
transform 1 0 31142 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1712078602
transform 1 0 31418 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1712078602
transform 1 0 31510 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1712078602
transform 1 0 32062 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1712078602
transform 1 0 32614 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1712078602
transform 1 0 33166 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1712078602
transform 1 0 33718 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1712078602
transform 1 0 33994 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1712078602
transform 1 0 34086 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1712078602
transform 1 0 34638 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1712078602
transform 1 0 35190 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1712078602
transform 1 0 35742 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1712078602
transform 1 0 36294 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1712078602
transform 1 0 36570 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1712078602
transform 1 0 36662 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1712078602
transform 1 0 37214 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1712078602
transform 1 0 37766 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_821
timestamp 1712078602
transform 1 0 38318 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1712078602
transform 1 0 38870 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1712078602
transform 1 0 39146 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1712078602
transform 1 0 39238 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1712078602
transform 1 0 39790 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1712078602
transform 1 0 40342 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1712078602
transform 1 0 40894 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1712078602
transform 1 0 41446 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1712078602
transform 1 0 41722 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1712078602
transform 1 0 41814 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_909
timestamp 1712078602
transform 1 0 42366 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_921
timestamp 1712078602
transform 1 0 42918 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_933
timestamp 1712078602
transform 1 0 43470 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1712078602
transform 1 0 44022 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1712078602
transform 1 0 44298 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_953
timestamp 1712078602
transform 1 0 44390 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_965
timestamp 1712078602
transform 1 0 44942 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_977
timestamp 1712078602
transform 1 0 45494 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_989
timestamp 1712078602
transform 1 0 46046 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1712078602
transform 1 0 46598 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1712078602
transform 1 0 46874 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1009
timestamp 1712078602
transform 1 0 46966 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1021
timestamp 1712078602
transform 1 0 47518 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1033
timestamp 1712078602
transform 1 0 48070 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1045
timestamp 1712078602
transform 1 0 48622 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1712078602
transform 1 0 49174 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1712078602
transform 1 0 49450 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1065
timestamp 1712078602
transform 1 0 49542 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1077
timestamp 1712078602
transform 1 0 50094 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1089
timestamp 1712078602
transform 1 0 50646 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1101
timestamp 1712078602
transform 1 0 51198 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1712078602
transform 1 0 51750 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1712078602
transform 1 0 52026 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1121
timestamp 1712078602
transform 1 0 52118 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1133
timestamp 1712078602
transform 1 0 52670 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1145
timestamp 1712078602
transform 1 0 53222 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1157
timestamp 1712078602
transform 1 0 53774 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1712078602
transform 1 0 54326 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1712078602
transform 1 0 54602 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1177
timestamp 1712078602
transform 1 0 54694 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1189
timestamp 1712078602
transform 1 0 55246 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1201
timestamp 1712078602
transform 1 0 55798 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1213
timestamp 1712078602
transform 1 0 56350 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1712078602
transform 1 0 56902 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1712078602
transform 1 0 57178 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1233
timestamp 1712078602
transform 1 0 57270 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1245
timestamp 1712078602
transform 1 0 57822 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1257
timestamp 1712078602
transform 1 0 58374 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1269
timestamp 1712078602
transform 1 0 58926 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1281
timestamp 1712078602
transform 1 0 59478 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1287
timestamp 1712078602
transform 1 0 59754 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1289
timestamp 1712078602
transform 1 0 59846 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1301
timestamp 1712078602
transform 1 0 60398 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1313
timestamp 1712078602
transform 1 0 60950 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1325
timestamp 1712078602
transform 1 0 61502 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1337
timestamp 1712078602
transform 1 0 62054 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1343
timestamp 1712078602
transform 1 0 62330 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1345
timestamp 1712078602
transform 1 0 62422 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1357
timestamp 1712078602
transform 1 0 62974 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1369
timestamp 1712078602
transform 1 0 63526 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1381
timestamp 1712078602
transform 1 0 64078 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1393
timestamp 1712078602
transform 1 0 64630 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1399
timestamp 1712078602
transform 1 0 64906 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1401
timestamp 1712078602
transform 1 0 64998 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1413
timestamp 1712078602
transform 1 0 65550 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1425
timestamp 1712078602
transform 1 0 66102 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1437
timestamp 1712078602
transform 1 0 66654 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1449
timestamp 1712078602
transform 1 0 67206 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1455
timestamp 1712078602
transform 1 0 67482 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1457
timestamp 1712078602
transform 1 0 67574 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1469
timestamp 1712078602
transform 1 0 68126 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1481
timestamp 1712078602
transform 1 0 68678 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1493
timestamp 1712078602
transform 1 0 69230 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1505
timestamp 1712078602
transform 1 0 69782 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1511
timestamp 1712078602
transform 1 0 70058 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1513
timestamp 1712078602
transform 1 0 70150 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1525
timestamp 1712078602
transform 1 0 70702 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1537
timestamp 1712078602
transform 1 0 71254 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1549
timestamp 1712078602
transform 1 0 71806 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1561
timestamp 1712078602
transform 1 0 72358 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1567
timestamp 1712078602
transform 1 0 72634 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1569
timestamp 1712078602
transform 1 0 72726 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1581
timestamp 1712078602
transform 1 0 73278 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1593
timestamp 1712078602
transform 1 0 73830 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1605
timestamp 1712078602
transform 1 0 74382 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1617
timestamp 1712078602
transform 1 0 74934 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1623
timestamp 1712078602
transform 1 0 75210 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1625
timestamp 1712078602
transform 1 0 75302 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1637
timestamp 1712078602
transform 1 0 75854 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1649
timestamp 1712078602
transform 1 0 76406 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1661
timestamp 1712078602
transform 1 0 76958 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1673
timestamp 1712078602
transform 1 0 77510 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1679
timestamp 1712078602
transform 1 0 77786 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1681
timestamp 1712078602
transform 1 0 77878 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1693
timestamp 1712078602
transform 1 0 78430 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1705
timestamp 1712078602
transform 1 0 78982 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1717
timestamp 1712078602
transform 1 0 79534 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1729
timestamp 1712078602
transform 1 0 80086 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1735
timestamp 1712078602
transform 1 0 80362 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1737
timestamp 1712078602
transform 1 0 80454 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1749
timestamp 1712078602
transform 1 0 81006 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1761
timestamp 1712078602
transform 1 0 81558 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1773
timestamp 1712078602
transform 1 0 82110 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1785
timestamp 1712078602
transform 1 0 82662 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1791
timestamp 1712078602
transform 1 0 82938 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1793
timestamp 1712078602
transform 1 0 83030 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1805
timestamp 1712078602
transform 1 0 83582 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1817
timestamp 1712078602
transform 1 0 84134 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1829
timestamp 1712078602
transform 1 0 84686 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1841
timestamp 1712078602
transform 1 0 85238 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1847
timestamp 1712078602
transform 1 0 85514 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1849
timestamp 1712078602
transform 1 0 85606 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1861
timestamp 1712078602
transform 1 0 86158 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1873
timestamp 1712078602
transform 1 0 86710 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1885
timestamp 1712078602
transform 1 0 87262 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1897
timestamp 1712078602
transform 1 0 87814 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1903
timestamp 1712078602
transform 1 0 88090 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1905
timestamp 1712078602
transform 1 0 88182 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1917
timestamp 1712078602
transform 1 0 88734 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1929
timestamp 1712078602
transform 1 0 89286 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1941
timestamp 1712078602
transform 1 0 89838 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_1953
timestamp 1712078602
transform 1 0 90390 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_1959
timestamp 1712078602
transform 1 0 90666 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1961
timestamp 1712078602
transform 1 0 90758 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1973
timestamp 1712078602
transform 1 0 91310 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1985
timestamp 1712078602
transform 1 0 91862 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_1997
timestamp 1712078602
transform 1 0 92414 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2009
timestamp 1712078602
transform 1 0 92966 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2015
timestamp 1712078602
transform 1 0 93242 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2017
timestamp 1712078602
transform 1 0 93334 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2029
timestamp 1712078602
transform 1 0 93886 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2041
timestamp 1712078602
transform 1 0 94438 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2053
timestamp 1712078602
transform 1 0 94990 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2065
timestamp 1712078602
transform 1 0 95542 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2071
timestamp 1712078602
transform 1 0 95818 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2073
timestamp 1712078602
transform 1 0 95910 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2085
timestamp 1712078602
transform 1 0 96462 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2097
timestamp 1712078602
transform 1 0 97014 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2109
timestamp 1712078602
transform 1 0 97566 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2121
timestamp 1712078602
transform 1 0 98118 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2127
timestamp 1712078602
transform 1 0 98394 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2129
timestamp 1712078602
transform 1 0 98486 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2141
timestamp 1712078602
transform 1 0 99038 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2153
timestamp 1712078602
transform 1 0 99590 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2165
timestamp 1712078602
transform 1 0 100142 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2177
timestamp 1712078602
transform 1 0 100694 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2183
timestamp 1712078602
transform 1 0 100970 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2185
timestamp 1712078602
transform 1 0 101062 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2197
timestamp 1712078602
transform 1 0 101614 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2209
timestamp 1712078602
transform 1 0 102166 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2221
timestamp 1712078602
transform 1 0 102718 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2233
timestamp 1712078602
transform 1 0 103270 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2239
timestamp 1712078602
transform 1 0 103546 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2241
timestamp 1712078602
transform 1 0 103638 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2253
timestamp 1712078602
transform 1 0 104190 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2265
timestamp 1712078602
transform 1 0 104742 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2277
timestamp 1712078602
transform 1 0 105294 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2289
timestamp 1712078602
transform 1 0 105846 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2295
timestamp 1712078602
transform 1 0 106122 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2297
timestamp 1712078602
transform 1 0 106214 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2309
timestamp 1712078602
transform 1 0 106766 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2321
timestamp 1712078602
transform 1 0 107318 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2333
timestamp 1712078602
transform 1 0 107870 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2345
timestamp 1712078602
transform 1 0 108422 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2351
timestamp 1712078602
transform 1 0 108698 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2353
timestamp 1712078602
transform 1 0 108790 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2365
timestamp 1712078602
transform 1 0 109342 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2377
timestamp 1712078602
transform 1 0 109894 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2389
timestamp 1712078602
transform 1 0 110446 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2401
timestamp 1712078602
transform 1 0 110998 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2407
timestamp 1712078602
transform 1 0 111274 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2409
timestamp 1712078602
transform 1 0 111366 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2421
timestamp 1712078602
transform 1 0 111918 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2433
timestamp 1712078602
transform 1 0 112470 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2445
timestamp 1712078602
transform 1 0 113022 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2457
timestamp 1712078602
transform 1 0 113574 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2463
timestamp 1712078602
transform 1 0 113850 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2465
timestamp 1712078602
transform 1 0 113942 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2477
timestamp 1712078602
transform 1 0 114494 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2489
timestamp 1712078602
transform 1 0 115046 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2501
timestamp 1712078602
transform 1 0 115598 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2513
timestamp 1712078602
transform 1 0 116150 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2519
timestamp 1712078602
transform 1 0 116426 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2521
timestamp 1712078602
transform 1 0 116518 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2533
timestamp 1712078602
transform 1 0 117070 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2545
timestamp 1712078602
transform 1 0 117622 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2557
timestamp 1712078602
transform 1 0 118174 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2569
timestamp 1712078602
transform 1 0 118726 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2575
timestamp 1712078602
transform 1 0 119002 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2577
timestamp 1712078602
transform 1 0 119094 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2589
timestamp 1712078602
transform 1 0 119646 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2601
timestamp 1712078602
transform 1 0 120198 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2613
timestamp 1712078602
transform 1 0 120750 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2625
timestamp 1712078602
transform 1 0 121302 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2631
timestamp 1712078602
transform 1 0 121578 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2633
timestamp 1712078602
transform 1 0 121670 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2645
timestamp 1712078602
transform 1 0 122222 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2657
timestamp 1712078602
transform 1 0 122774 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2669
timestamp 1712078602
transform 1 0 123326 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2681
timestamp 1712078602
transform 1 0 123878 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2687
timestamp 1712078602
transform 1 0 124154 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2689
timestamp 1712078602
transform 1 0 124246 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2701
timestamp 1712078602
transform 1 0 124798 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2713
timestamp 1712078602
transform 1 0 125350 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2725
timestamp 1712078602
transform 1 0 125902 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2737
timestamp 1712078602
transform 1 0 126454 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2743
timestamp 1712078602
transform 1 0 126730 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2745
timestamp 1712078602
transform 1 0 126822 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2757
timestamp 1712078602
transform 1 0 127374 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2769
timestamp 1712078602
transform 1 0 127926 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2781
timestamp 1712078602
transform 1 0 128478 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2793
timestamp 1712078602
transform 1 0 129030 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2799
timestamp 1712078602
transform 1 0 129306 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2801
timestamp 1712078602
transform 1 0 129398 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2813
timestamp 1712078602
transform 1 0 129950 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2825
timestamp 1712078602
transform 1 0 130502 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2837
timestamp 1712078602
transform 1 0 131054 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2849
timestamp 1712078602
transform 1 0 131606 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2855
timestamp 1712078602
transform 1 0 131882 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2857
timestamp 1712078602
transform 1 0 131974 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2869
timestamp 1712078602
transform 1 0 132526 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2881
timestamp 1712078602
transform 1 0 133078 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2893
timestamp 1712078602
transform 1 0 133630 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2905
timestamp 1712078602
transform 1 0 134182 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2911
timestamp 1712078602
transform 1 0 134458 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2913
timestamp 1712078602
transform 1 0 134550 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2925
timestamp 1712078602
transform 1 0 135102 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2937
timestamp 1712078602
transform 1 0 135654 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2949
timestamp 1712078602
transform 1 0 136206 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_2961
timestamp 1712078602
transform 1 0 136758 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_2967
timestamp 1712078602
transform 1 0 137034 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2969
timestamp 1712078602
transform 1 0 137126 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2981
timestamp 1712078602
transform 1 0 137678 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_2993
timestamp 1712078602
transform 1 0 138230 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3005
timestamp 1712078602
transform 1 0 138782 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_3017
timestamp 1712078602
transform 1 0 139334 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_3023
timestamp 1712078602
transform 1 0 139610 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3025
timestamp 1712078602
transform 1 0 139702 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3037
timestamp 1712078602
transform 1 0 140254 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3049
timestamp 1712078602
transform 1 0 140806 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3061
timestamp 1712078602
transform 1 0 141358 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_3073
timestamp 1712078602
transform 1 0 141910 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_3079
timestamp 1712078602
transform 1 0 142186 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3081
timestamp 1712078602
transform 1 0 142278 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3093
timestamp 1712078602
transform 1 0 142830 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3105
timestamp 1712078602
transform 1 0 143382 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3117
timestamp 1712078602
transform 1 0 143934 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_3129
timestamp 1712078602
transform 1 0 144486 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_3135
timestamp 1712078602
transform 1 0 144762 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3137
timestamp 1712078602
transform 1 0 144854 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3149
timestamp 1712078602
transform 1 0 145406 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3161
timestamp 1712078602
transform 1 0 145958 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3173
timestamp 1712078602
transform 1 0 146510 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_3185
timestamp 1712078602
transform 1 0 147062 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_3191
timestamp 1712078602
transform 1 0 147338 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3193
timestamp 1712078602
transform 1 0 147430 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3205
timestamp 1712078602
transform 1 0 147982 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3217
timestamp 1712078602
transform 1 0 148534 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3229
timestamp 1712078602
transform 1 0 149086 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_3241
timestamp 1712078602
transform 1 0 149638 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_3247
timestamp 1712078602
transform 1 0 149914 0 -1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3249
timestamp 1712078602
transform 1 0 150006 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3261
timestamp 1712078602
transform 1 0 150558 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3273
timestamp 1712078602
transform 1 0 151110 0 -1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_11_3285
timestamp 1712078602
transform 1 0 151662 0 -1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_11_3297
timestamp 1712078602
transform 1 0 152214 0 -1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_11_3303
timestamp 1712078602
transform 1 0 152490 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_11_3305
timestamp 1712078602
transform 1 0 152582 0 -1 4352
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1712078602
transform 1 0 690 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1712078602
transform 1 0 1242 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1712078602
transform 1 0 1794 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1712078602
transform 1 0 1886 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1712078602
transform 1 0 2438 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1712078602
transform 1 0 2990 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1712078602
transform 1 0 3542 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1712078602
transform 1 0 4094 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1712078602
transform 1 0 4370 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1712078602
transform 1 0 4462 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1712078602
transform 1 0 5014 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1712078602
transform 1 0 5566 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1712078602
transform 1 0 6118 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1712078602
transform 1 0 6670 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1712078602
transform 1 0 6946 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1712078602
transform 1 0 7038 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1712078602
transform 1 0 7590 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1712078602
transform 1 0 8142 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1712078602
transform 1 0 8694 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1712078602
transform 1 0 9246 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1712078602
transform 1 0 9522 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1712078602
transform 1 0 9614 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1712078602
transform 1 0 10166 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1712078602
transform 1 0 10718 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1712078602
transform 1 0 11270 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1712078602
transform 1 0 11822 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1712078602
transform 1 0 12098 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1712078602
transform 1 0 12190 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1712078602
transform 1 0 12742 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1712078602
transform 1 0 13294 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1712078602
transform 1 0 13846 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1712078602
transform 1 0 14398 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1712078602
transform 1 0 14674 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1712078602
transform 1 0 14766 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1712078602
transform 1 0 15318 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1712078602
transform 1 0 15870 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1712078602
transform 1 0 16422 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1712078602
transform 1 0 16974 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1712078602
transform 1 0 17250 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1712078602
transform 1 0 17342 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1712078602
transform 1 0 17894 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1712078602
transform 1 0 18446 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1712078602
transform 1 0 18998 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1712078602
transform 1 0 19550 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1712078602
transform 1 0 19826 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1712078602
transform 1 0 19918 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1712078602
transform 1 0 20470 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1712078602
transform 1 0 21022 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1712078602
transform 1 0 21574 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1712078602
transform 1 0 22126 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1712078602
transform 1 0 22402 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1712078602
transform 1 0 22494 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1712078602
transform 1 0 23046 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1712078602
transform 1 0 23598 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1712078602
transform 1 0 24150 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1712078602
transform 1 0 24702 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1712078602
transform 1 0 24978 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1712078602
transform 1 0 25070 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1712078602
transform 1 0 25622 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1712078602
transform 1 0 26174 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1712078602
transform 1 0 26726 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1712078602
transform 1 0 27278 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1712078602
transform 1 0 27554 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1712078602
transform 1 0 27646 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1712078602
transform 1 0 28198 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1712078602
transform 1 0 28750 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1712078602
transform 1 0 29302 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1712078602
transform 1 0 29854 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1712078602
transform 1 0 30130 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1712078602
transform 1 0 30222 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1712078602
transform 1 0 30774 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1712078602
transform 1 0 31326 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1712078602
transform 1 0 31878 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1712078602
transform 1 0 32430 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1712078602
transform 1 0 32706 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1712078602
transform 1 0 32798 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1712078602
transform 1 0 33350 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1712078602
transform 1 0 33902 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1712078602
transform 1 0 34454 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1712078602
transform 1 0 35006 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1712078602
transform 1 0 35282 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1712078602
transform 1 0 35374 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1712078602
transform 1 0 35926 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1712078602
transform 1 0 36478 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1712078602
transform 1 0 37030 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1712078602
transform 1 0 37582 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1712078602
transform 1 0 37858 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1712078602
transform 1 0 37950 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1712078602
transform 1 0 38502 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_837
timestamp 1712078602
transform 1 0 39054 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_849
timestamp 1712078602
transform 1 0 39606 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1712078602
transform 1 0 40158 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1712078602
transform 1 0 40434 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1712078602
transform 1 0 40526 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1712078602
transform 1 0 41078 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1712078602
transform 1 0 41630 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1712078602
transform 1 0 42182 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1712078602
transform 1 0 42734 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1712078602
transform 1 0 43010 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_925
timestamp 1712078602
transform 1 0 43102 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_937
timestamp 1712078602
transform 1 0 43654 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_949
timestamp 1712078602
transform 1 0 44206 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_961
timestamp 1712078602
transform 1 0 44758 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1712078602
transform 1 0 45310 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1712078602
transform 1 0 45586 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_981
timestamp 1712078602
transform 1 0 45678 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_993
timestamp 1712078602
transform 1 0 46230 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1005
timestamp 1712078602
transform 1 0 46782 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1017
timestamp 1712078602
transform 1 0 47334 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1712078602
transform 1 0 47886 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1712078602
transform 1 0 48162 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1037
timestamp 1712078602
transform 1 0 48254 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1049
timestamp 1712078602
transform 1 0 48806 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1061
timestamp 1712078602
transform 1 0 49358 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1073
timestamp 1712078602
transform 1 0 49910 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1712078602
transform 1 0 50462 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1712078602
transform 1 0 50738 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1093
timestamp 1712078602
transform 1 0 50830 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1105
timestamp 1712078602
transform 1 0 51382 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1117
timestamp 1712078602
transform 1 0 51934 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1129
timestamp 1712078602
transform 1 0 52486 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1712078602
transform 1 0 53038 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1712078602
transform 1 0 53314 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1149
timestamp 1712078602
transform 1 0 53406 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1161
timestamp 1712078602
transform 1 0 53958 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1173
timestamp 1712078602
transform 1 0 54510 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1185
timestamp 1712078602
transform 1 0 55062 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1712078602
transform 1 0 55614 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1712078602
transform 1 0 55890 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1205
timestamp 1712078602
transform 1 0 55982 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1217
timestamp 1712078602
transform 1 0 56534 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1229
timestamp 1712078602
transform 1 0 57086 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1241
timestamp 1712078602
transform 1 0 57638 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1712078602
transform 1 0 58190 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1712078602
transform 1 0 58466 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1261
timestamp 1712078602
transform 1 0 58558 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1273
timestamp 1712078602
transform 1 0 59110 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1285
timestamp 1712078602
transform 1 0 59662 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1297
timestamp 1712078602
transform 1 0 60214 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1309
timestamp 1712078602
transform 1 0 60766 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1315
timestamp 1712078602
transform 1 0 61042 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1317
timestamp 1712078602
transform 1 0 61134 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1329
timestamp 1712078602
transform 1 0 61686 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1341
timestamp 1712078602
transform 1 0 62238 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1353
timestamp 1712078602
transform 1 0 62790 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1365
timestamp 1712078602
transform 1 0 63342 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1371
timestamp 1712078602
transform 1 0 63618 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1373
timestamp 1712078602
transform 1 0 63710 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1385
timestamp 1712078602
transform 1 0 64262 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1397
timestamp 1712078602
transform 1 0 64814 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1409
timestamp 1712078602
transform 1 0 65366 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1421
timestamp 1712078602
transform 1 0 65918 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1427
timestamp 1712078602
transform 1 0 66194 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1429
timestamp 1712078602
transform 1 0 66286 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1441
timestamp 1712078602
transform 1 0 66838 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1453
timestamp 1712078602
transform 1 0 67390 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1465
timestamp 1712078602
transform 1 0 67942 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1477
timestamp 1712078602
transform 1 0 68494 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1483
timestamp 1712078602
transform 1 0 68770 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1485
timestamp 1712078602
transform 1 0 68862 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1497
timestamp 1712078602
transform 1 0 69414 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1509
timestamp 1712078602
transform 1 0 69966 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1521
timestamp 1712078602
transform 1 0 70518 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1533
timestamp 1712078602
transform 1 0 71070 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1539
timestamp 1712078602
transform 1 0 71346 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1541
timestamp 1712078602
transform 1 0 71438 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1553
timestamp 1712078602
transform 1 0 71990 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1565
timestamp 1712078602
transform 1 0 72542 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1577
timestamp 1712078602
transform 1 0 73094 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1589
timestamp 1712078602
transform 1 0 73646 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1595
timestamp 1712078602
transform 1 0 73922 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1597
timestamp 1712078602
transform 1 0 74014 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1609
timestamp 1712078602
transform 1 0 74566 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1621
timestamp 1712078602
transform 1 0 75118 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1633
timestamp 1712078602
transform 1 0 75670 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1645
timestamp 1712078602
transform 1 0 76222 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1651
timestamp 1712078602
transform 1 0 76498 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1653
timestamp 1712078602
transform 1 0 76590 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1665
timestamp 1712078602
transform 1 0 77142 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1677
timestamp 1712078602
transform 1 0 77694 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1689
timestamp 1712078602
transform 1 0 78246 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1701
timestamp 1712078602
transform 1 0 78798 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1707
timestamp 1712078602
transform 1 0 79074 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1709
timestamp 1712078602
transform 1 0 79166 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1721
timestamp 1712078602
transform 1 0 79718 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1733
timestamp 1712078602
transform 1 0 80270 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1745
timestamp 1712078602
transform 1 0 80822 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1757
timestamp 1712078602
transform 1 0 81374 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1763
timestamp 1712078602
transform 1 0 81650 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1765
timestamp 1712078602
transform 1 0 81742 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1777
timestamp 1712078602
transform 1 0 82294 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1789
timestamp 1712078602
transform 1 0 82846 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1801
timestamp 1712078602
transform 1 0 83398 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1813
timestamp 1712078602
transform 1 0 83950 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1819
timestamp 1712078602
transform 1 0 84226 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1821
timestamp 1712078602
transform 1 0 84318 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1833
timestamp 1712078602
transform 1 0 84870 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1845
timestamp 1712078602
transform 1 0 85422 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1857
timestamp 1712078602
transform 1 0 85974 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1869
timestamp 1712078602
transform 1 0 86526 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1875
timestamp 1712078602
transform 1 0 86802 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1877
timestamp 1712078602
transform 1 0 86894 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1889
timestamp 1712078602
transform 1 0 87446 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1901
timestamp 1712078602
transform 1 0 87998 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1913
timestamp 1712078602
transform 1 0 88550 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1925
timestamp 1712078602
transform 1 0 89102 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1931
timestamp 1712078602
transform 1 0 89378 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1933
timestamp 1712078602
transform 1 0 89470 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1945
timestamp 1712078602
transform 1 0 90022 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1957
timestamp 1712078602
transform 1 0 90574 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1969
timestamp 1712078602
transform 1 0 91126 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_1981
timestamp 1712078602
transform 1 0 91678 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_1987
timestamp 1712078602
transform 1 0 91954 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_1989
timestamp 1712078602
transform 1 0 92046 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2001
timestamp 1712078602
transform 1 0 92598 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2013
timestamp 1712078602
transform 1 0 93150 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2025
timestamp 1712078602
transform 1 0 93702 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2037
timestamp 1712078602
transform 1 0 94254 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2043
timestamp 1712078602
transform 1 0 94530 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2045
timestamp 1712078602
transform 1 0 94622 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2057
timestamp 1712078602
transform 1 0 95174 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2069
timestamp 1712078602
transform 1 0 95726 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2081
timestamp 1712078602
transform 1 0 96278 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2093
timestamp 1712078602
transform 1 0 96830 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2099
timestamp 1712078602
transform 1 0 97106 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2101
timestamp 1712078602
transform 1 0 97198 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2113
timestamp 1712078602
transform 1 0 97750 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2125
timestamp 1712078602
transform 1 0 98302 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2137
timestamp 1712078602
transform 1 0 98854 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2149
timestamp 1712078602
transform 1 0 99406 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2155
timestamp 1712078602
transform 1 0 99682 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2157
timestamp 1712078602
transform 1 0 99774 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2169
timestamp 1712078602
transform 1 0 100326 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2181
timestamp 1712078602
transform 1 0 100878 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2193
timestamp 1712078602
transform 1 0 101430 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2205
timestamp 1712078602
transform 1 0 101982 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2211
timestamp 1712078602
transform 1 0 102258 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2213
timestamp 1712078602
transform 1 0 102350 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2225
timestamp 1712078602
transform 1 0 102902 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2237
timestamp 1712078602
transform 1 0 103454 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2249
timestamp 1712078602
transform 1 0 104006 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2261
timestamp 1712078602
transform 1 0 104558 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2267
timestamp 1712078602
transform 1 0 104834 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2269
timestamp 1712078602
transform 1 0 104926 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2281
timestamp 1712078602
transform 1 0 105478 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2293
timestamp 1712078602
transform 1 0 106030 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2305
timestamp 1712078602
transform 1 0 106582 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2317
timestamp 1712078602
transform 1 0 107134 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2323
timestamp 1712078602
transform 1 0 107410 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2325
timestamp 1712078602
transform 1 0 107502 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2337
timestamp 1712078602
transform 1 0 108054 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2349
timestamp 1712078602
transform 1 0 108606 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2361
timestamp 1712078602
transform 1 0 109158 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2373
timestamp 1712078602
transform 1 0 109710 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2379
timestamp 1712078602
transform 1 0 109986 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2381
timestamp 1712078602
transform 1 0 110078 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2393
timestamp 1712078602
transform 1 0 110630 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2405
timestamp 1712078602
transform 1 0 111182 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2417
timestamp 1712078602
transform 1 0 111734 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2429
timestamp 1712078602
transform 1 0 112286 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2435
timestamp 1712078602
transform 1 0 112562 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2437
timestamp 1712078602
transform 1 0 112654 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2449
timestamp 1712078602
transform 1 0 113206 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2461
timestamp 1712078602
transform 1 0 113758 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2473
timestamp 1712078602
transform 1 0 114310 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2485
timestamp 1712078602
transform 1 0 114862 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2491
timestamp 1712078602
transform 1 0 115138 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2493
timestamp 1712078602
transform 1 0 115230 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2505
timestamp 1712078602
transform 1 0 115782 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2517
timestamp 1712078602
transform 1 0 116334 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2529
timestamp 1712078602
transform 1 0 116886 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2541
timestamp 1712078602
transform 1 0 117438 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2547
timestamp 1712078602
transform 1 0 117714 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2549
timestamp 1712078602
transform 1 0 117806 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2561
timestamp 1712078602
transform 1 0 118358 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2573
timestamp 1712078602
transform 1 0 118910 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2585
timestamp 1712078602
transform 1 0 119462 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2597
timestamp 1712078602
transform 1 0 120014 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2603
timestamp 1712078602
transform 1 0 120290 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2605
timestamp 1712078602
transform 1 0 120382 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2617
timestamp 1712078602
transform 1 0 120934 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2629
timestamp 1712078602
transform 1 0 121486 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2641
timestamp 1712078602
transform 1 0 122038 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2653
timestamp 1712078602
transform 1 0 122590 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2659
timestamp 1712078602
transform 1 0 122866 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2661
timestamp 1712078602
transform 1 0 122958 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2673
timestamp 1712078602
transform 1 0 123510 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2685
timestamp 1712078602
transform 1 0 124062 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2697
timestamp 1712078602
transform 1 0 124614 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2709
timestamp 1712078602
transform 1 0 125166 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2715
timestamp 1712078602
transform 1 0 125442 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2717
timestamp 1712078602
transform 1 0 125534 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2729
timestamp 1712078602
transform 1 0 126086 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2741
timestamp 1712078602
transform 1 0 126638 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2753
timestamp 1712078602
transform 1 0 127190 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2765
timestamp 1712078602
transform 1 0 127742 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2771
timestamp 1712078602
transform 1 0 128018 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2773
timestamp 1712078602
transform 1 0 128110 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2785
timestamp 1712078602
transform 1 0 128662 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2797
timestamp 1712078602
transform 1 0 129214 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2809
timestamp 1712078602
transform 1 0 129766 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2821
timestamp 1712078602
transform 1 0 130318 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2827
timestamp 1712078602
transform 1 0 130594 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2829
timestamp 1712078602
transform 1 0 130686 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2841
timestamp 1712078602
transform 1 0 131238 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2853
timestamp 1712078602
transform 1 0 131790 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2865
timestamp 1712078602
transform 1 0 132342 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2877
timestamp 1712078602
transform 1 0 132894 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2883
timestamp 1712078602
transform 1 0 133170 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2885
timestamp 1712078602
transform 1 0 133262 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2897
timestamp 1712078602
transform 1 0 133814 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2909
timestamp 1712078602
transform 1 0 134366 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2921
timestamp 1712078602
transform 1 0 134918 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2933
timestamp 1712078602
transform 1 0 135470 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2939
timestamp 1712078602
transform 1 0 135746 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2941
timestamp 1712078602
transform 1 0 135838 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2953
timestamp 1712078602
transform 1 0 136390 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2965
timestamp 1712078602
transform 1 0 136942 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2977
timestamp 1712078602
transform 1 0 137494 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_2989
timestamp 1712078602
transform 1 0 138046 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_2995
timestamp 1712078602
transform 1 0 138322 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_2997
timestamp 1712078602
transform 1 0 138414 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3009
timestamp 1712078602
transform 1 0 138966 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3021
timestamp 1712078602
transform 1 0 139518 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3033
timestamp 1712078602
transform 1 0 140070 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_3045
timestamp 1712078602
transform 1 0 140622 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_3051
timestamp 1712078602
transform 1 0 140898 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3053
timestamp 1712078602
transform 1 0 140990 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3065
timestamp 1712078602
transform 1 0 141542 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3077
timestamp 1712078602
transform 1 0 142094 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3089
timestamp 1712078602
transform 1 0 142646 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_3101
timestamp 1712078602
transform 1 0 143198 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_3107
timestamp 1712078602
transform 1 0 143474 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3109
timestamp 1712078602
transform 1 0 143566 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3121
timestamp 1712078602
transform 1 0 144118 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3133
timestamp 1712078602
transform 1 0 144670 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3145
timestamp 1712078602
transform 1 0 145222 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_3157
timestamp 1712078602
transform 1 0 145774 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_3163
timestamp 1712078602
transform 1 0 146050 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3165
timestamp 1712078602
transform 1 0 146142 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3177
timestamp 1712078602
transform 1 0 146694 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3189
timestamp 1712078602
transform 1 0 147246 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3201
timestamp 1712078602
transform 1 0 147798 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_3213
timestamp 1712078602
transform 1 0 148350 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_3219
timestamp 1712078602
transform 1 0 148626 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3221
timestamp 1712078602
transform 1 0 148718 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3233
timestamp 1712078602
transform 1 0 149270 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3245
timestamp 1712078602
transform 1 0 149822 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3257
timestamp 1712078602
transform 1 0 150374 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_12_3269
timestamp 1712078602
transform 1 0 150926 0 1 4352
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_12_3275
timestamp 1712078602
transform 1 0 151202 0 1 4352
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3277
timestamp 1712078602
transform 1 0 151294 0 1 4352
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_12_3289
timestamp 1712078602
transform 1 0 151846 0 1 4352
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_12_3301
timestamp 1712078602
transform 1 0 152398 0 1 4352
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1712078602
transform 1 0 690 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1712078602
transform 1 0 1242 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1712078602
transform 1 0 1794 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1712078602
transform 1 0 2346 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1712078602
transform 1 0 2898 0 -1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1712078602
transform 1 0 3082 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1712078602
transform 1 0 3174 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1712078602
transform 1 0 3726 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1712078602
transform 1 0 4278 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1712078602
transform 1 0 4830 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1712078602
transform 1 0 5382 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1712078602
transform 1 0 5658 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1712078602
transform 1 0 5750 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1712078602
transform 1 0 6302 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1712078602
transform 1 0 6854 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1712078602
transform 1 0 7406 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1712078602
transform 1 0 7958 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1712078602
transform 1 0 8234 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1712078602
transform 1 0 8326 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1712078602
transform 1 0 8878 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1712078602
transform 1 0 9430 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1712078602
transform 1 0 9982 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1712078602
transform 1 0 10534 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1712078602
transform 1 0 10810 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1712078602
transform 1 0 10902 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1712078602
transform 1 0 11454 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1712078602
transform 1 0 12006 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1712078602
transform 1 0 12558 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1712078602
transform 1 0 13110 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1712078602
transform 1 0 13386 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1712078602
transform 1 0 13478 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1712078602
transform 1 0 14030 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1712078602
transform 1 0 14582 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_13_317
timestamp 1712078602
transform 1 0 15134 0 -1 4896
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_13_325
timestamp 1712078602
transform 1 0 15502 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1712078602
transform 1 0 15686 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1712078602
transform 1 0 15962 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_13_340
timestamp 1712078602
transform 1 0 16192 0 -1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_13_347
timestamp 1712078602
transform 1 0 16514 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_359
timestamp 1712078602
transform 1 0 17066 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_371
timestamp 1712078602
transform 1 0 17618 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_13_383
timestamp 1712078602
transform 1 0 18170 0 -1 4896
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1712078602
transform 1 0 18538 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1712078602
transform 1 0 18630 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1712078602
transform 1 0 19182 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1712078602
transform 1 0 19734 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1712078602
transform 1 0 20286 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1712078602
transform 1 0 20838 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1712078602
transform 1 0 21114 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1712078602
transform 1 0 21206 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1712078602
transform 1 0 21758 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1712078602
transform 1 0 22310 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1712078602
transform 1 0 22862 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1712078602
transform 1 0 23414 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1712078602
transform 1 0 23690 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1712078602
transform 1 0 23782 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1712078602
transform 1 0 24334 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1712078602
transform 1 0 24886 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1712078602
transform 1 0 25438 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1712078602
transform 1 0 25990 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1712078602
transform 1 0 26266 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1712078602
transform 1 0 26358 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1712078602
transform 1 0 26910 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1712078602
transform 1 0 27462 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1712078602
transform 1 0 28014 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1712078602
transform 1 0 28566 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1712078602
transform 1 0 28842 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1712078602
transform 1 0 28934 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1712078602
transform 1 0 29486 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1712078602
transform 1 0 30038 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1712078602
transform 1 0 30590 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1712078602
transform 1 0 31142 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1712078602
transform 1 0 31418 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1712078602
transform 1 0 31510 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1712078602
transform 1 0 32062 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1712078602
transform 1 0 32614 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1712078602
transform 1 0 33166 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1712078602
transform 1 0 33718 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1712078602
transform 1 0 33994 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1712078602
transform 1 0 34086 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1712078602
transform 1 0 34638 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1712078602
transform 1 0 35190 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1712078602
transform 1 0 35742 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1712078602
transform 1 0 36294 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1712078602
transform 1 0 36570 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1712078602
transform 1 0 36662 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1712078602
transform 1 0 37214 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1712078602
transform 1 0 37766 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_821
timestamp 1712078602
transform 1 0 38318 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1712078602
transform 1 0 38870 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1712078602
transform 1 0 39146 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1712078602
transform 1 0 39238 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_853
timestamp 1712078602
transform 1 0 39790 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_865
timestamp 1712078602
transform 1 0 40342 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_877
timestamp 1712078602
transform 1 0 40894 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1712078602
transform 1 0 41446 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1712078602
transform 1 0 41722 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1712078602
transform 1 0 41814 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_909
timestamp 1712078602
transform 1 0 42366 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_921
timestamp 1712078602
transform 1 0 42918 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_933
timestamp 1712078602
transform 1 0 43470 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1712078602
transform 1 0 44022 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_951
timestamp 1712078602
transform 1 0 44298 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_953
timestamp 1712078602
transform 1 0 44390 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_965
timestamp 1712078602
transform 1 0 44942 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_977
timestamp 1712078602
transform 1 0 45494 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_989
timestamp 1712078602
transform 1 0 46046 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1001
timestamp 1712078602
transform 1 0 46598 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1712078602
transform 1 0 46874 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1009
timestamp 1712078602
transform 1 0 46966 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1021
timestamp 1712078602
transform 1 0 47518 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1033
timestamp 1712078602
transform 1 0 48070 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1045
timestamp 1712078602
transform 1 0 48622 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1057
timestamp 1712078602
transform 1 0 49174 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1063
timestamp 1712078602
transform 1 0 49450 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1065
timestamp 1712078602
transform 1 0 49542 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1077
timestamp 1712078602
transform 1 0 50094 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1089
timestamp 1712078602
transform 1 0 50646 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1101
timestamp 1712078602
transform 1 0 51198 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1712078602
transform 1 0 51750 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1712078602
transform 1 0 52026 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1121
timestamp 1712078602
transform 1 0 52118 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1133
timestamp 1712078602
transform 1 0 52670 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1145
timestamp 1712078602
transform 1 0 53222 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1157
timestamp 1712078602
transform 1 0 53774 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1712078602
transform 1 0 54326 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1712078602
transform 1 0 54602 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1177
timestamp 1712078602
transform 1 0 54694 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1189
timestamp 1712078602
transform 1 0 55246 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1201
timestamp 1712078602
transform 1 0 55798 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1213
timestamp 1712078602
transform 1 0 56350 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1225
timestamp 1712078602
transform 1 0 56902 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1231
timestamp 1712078602
transform 1 0 57178 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1233
timestamp 1712078602
transform 1 0 57270 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1245
timestamp 1712078602
transform 1 0 57822 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1257
timestamp 1712078602
transform 1 0 58374 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1269
timestamp 1712078602
transform 1 0 58926 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1281
timestamp 1712078602
transform 1 0 59478 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1287
timestamp 1712078602
transform 1 0 59754 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1289
timestamp 1712078602
transform 1 0 59846 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1301
timestamp 1712078602
transform 1 0 60398 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1313
timestamp 1712078602
transform 1 0 60950 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1325
timestamp 1712078602
transform 1 0 61502 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1337
timestamp 1712078602
transform 1 0 62054 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1343
timestamp 1712078602
transform 1 0 62330 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1345
timestamp 1712078602
transform 1 0 62422 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1357
timestamp 1712078602
transform 1 0 62974 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1369
timestamp 1712078602
transform 1 0 63526 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1381
timestamp 1712078602
transform 1 0 64078 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1393
timestamp 1712078602
transform 1 0 64630 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1399
timestamp 1712078602
transform 1 0 64906 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1401
timestamp 1712078602
transform 1 0 64998 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1413
timestamp 1712078602
transform 1 0 65550 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1425
timestamp 1712078602
transform 1 0 66102 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1437
timestamp 1712078602
transform 1 0 66654 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1449
timestamp 1712078602
transform 1 0 67206 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1455
timestamp 1712078602
transform 1 0 67482 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1457
timestamp 1712078602
transform 1 0 67574 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1469
timestamp 1712078602
transform 1 0 68126 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1481
timestamp 1712078602
transform 1 0 68678 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1493
timestamp 1712078602
transform 1 0 69230 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1505
timestamp 1712078602
transform 1 0 69782 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1511
timestamp 1712078602
transform 1 0 70058 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_13_1513
timestamp 1712078602
transform 1 0 70150 0 -1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1537
timestamp 1712078602
transform 1 0 71254 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1549
timestamp 1712078602
transform 1 0 71806 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1561
timestamp 1712078602
transform 1 0 72358 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1567
timestamp 1712078602
transform 1 0 72634 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1569
timestamp 1712078602
transform 1 0 72726 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1581
timestamp 1712078602
transform 1 0 73278 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1593
timestamp 1712078602
transform 1 0 73830 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1605
timestamp 1712078602
transform 1 0 74382 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1617
timestamp 1712078602
transform 1 0 74934 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1623
timestamp 1712078602
transform 1 0 75210 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1625
timestamp 1712078602
transform 1 0 75302 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1637
timestamp 1712078602
transform 1 0 75854 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1649
timestamp 1712078602
transform 1 0 76406 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1661
timestamp 1712078602
transform 1 0 76958 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1673
timestamp 1712078602
transform 1 0 77510 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1679
timestamp 1712078602
transform 1 0 77786 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_13_1681
timestamp 1712078602
transform 1 0 77878 0 -1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1705
timestamp 1712078602
transform 1 0 78982 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1717
timestamp 1712078602
transform 1 0 79534 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1729
timestamp 1712078602
transform 1 0 80086 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1735
timestamp 1712078602
transform 1 0 80362 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1737
timestamp 1712078602
transform 1 0 80454 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1749
timestamp 1712078602
transform 1 0 81006 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1761
timestamp 1712078602
transform 1 0 81558 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1773
timestamp 1712078602
transform 1 0 82110 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1785
timestamp 1712078602
transform 1 0 82662 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1791
timestamp 1712078602
transform 1 0 82938 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1793
timestamp 1712078602
transform 1 0 83030 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1805
timestamp 1712078602
transform 1 0 83582 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1817
timestamp 1712078602
transform 1 0 84134 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1829
timestamp 1712078602
transform 1 0 84686 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1841
timestamp 1712078602
transform 1 0 85238 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1847
timestamp 1712078602
transform 1 0 85514 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1849
timestamp 1712078602
transform 1 0 85606 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1861
timestamp 1712078602
transform 1 0 86158 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1873
timestamp 1712078602
transform 1 0 86710 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1885
timestamp 1712078602
transform 1 0 87262 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1897
timestamp 1712078602
transform 1 0 87814 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1903
timestamp 1712078602
transform 1 0 88090 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1905
timestamp 1712078602
transform 1 0 88182 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1917
timestamp 1712078602
transform 1 0 88734 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1929
timestamp 1712078602
transform 1 0 89286 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1941
timestamp 1712078602
transform 1 0 89838 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_1953
timestamp 1712078602
transform 1 0 90390 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_1959
timestamp 1712078602
transform 1 0 90666 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1961
timestamp 1712078602
transform 1 0 90758 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1973
timestamp 1712078602
transform 1 0 91310 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1985
timestamp 1712078602
transform 1 0 91862 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_1997
timestamp 1712078602
transform 1 0 92414 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2009
timestamp 1712078602
transform 1 0 92966 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2015
timestamp 1712078602
transform 1 0 93242 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2017
timestamp 1712078602
transform 1 0 93334 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2029
timestamp 1712078602
transform 1 0 93886 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2041
timestamp 1712078602
transform 1 0 94438 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2053
timestamp 1712078602
transform 1 0 94990 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2065
timestamp 1712078602
transform 1 0 95542 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2071
timestamp 1712078602
transform 1 0 95818 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_13_2073
timestamp 1712078602
transform 1 0 95910 0 -1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2077
timestamp 1712078602
transform 1 0 96094 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_13_2081
timestamp 1712078602
transform 1 0 96278 0 -1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2088
timestamp 1712078602
transform 1 0 96600 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2100
timestamp 1712078602
transform 1 0 97152 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2112
timestamp 1712078602
transform 1 0 97704 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_13_2124
timestamp 1712078602
transform 1 0 98256 0 -1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2129
timestamp 1712078602
transform 1 0 98486 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2141
timestamp 1712078602
transform 1 0 99038 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2153
timestamp 1712078602
transform 1 0 99590 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2165
timestamp 1712078602
transform 1 0 100142 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2177
timestamp 1712078602
transform 1 0 100694 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2183
timestamp 1712078602
transform 1 0 100970 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2185
timestamp 1712078602
transform 1 0 101062 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2197
timestamp 1712078602
transform 1 0 101614 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2209
timestamp 1712078602
transform 1 0 102166 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2221
timestamp 1712078602
transform 1 0 102718 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2233
timestamp 1712078602
transform 1 0 103270 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2239
timestamp 1712078602
transform 1 0 103546 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2241
timestamp 1712078602
transform 1 0 103638 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2253
timestamp 1712078602
transform 1 0 104190 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2265
timestamp 1712078602
transform 1 0 104742 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2277
timestamp 1712078602
transform 1 0 105294 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2289
timestamp 1712078602
transform 1 0 105846 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2295
timestamp 1712078602
transform 1 0 106122 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2297
timestamp 1712078602
transform 1 0 106214 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2309
timestamp 1712078602
transform 1 0 106766 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2321
timestamp 1712078602
transform 1 0 107318 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2333
timestamp 1712078602
transform 1 0 107870 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2345
timestamp 1712078602
transform 1 0 108422 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2351
timestamp 1712078602
transform 1 0 108698 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2353
timestamp 1712078602
transform 1 0 108790 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2365
timestamp 1712078602
transform 1 0 109342 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2377
timestamp 1712078602
transform 1 0 109894 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2389
timestamp 1712078602
transform 1 0 110446 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2401
timestamp 1712078602
transform 1 0 110998 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2407
timestamp 1712078602
transform 1 0 111274 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2409
timestamp 1712078602
transform 1 0 111366 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2421
timestamp 1712078602
transform 1 0 111918 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2433
timestamp 1712078602
transform 1 0 112470 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2445
timestamp 1712078602
transform 1 0 113022 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2457
timestamp 1712078602
transform 1 0 113574 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2463
timestamp 1712078602
transform 1 0 113850 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2465
timestamp 1712078602
transform 1 0 113942 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2477
timestamp 1712078602
transform 1 0 114494 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2489
timestamp 1712078602
transform 1 0 115046 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2501
timestamp 1712078602
transform 1 0 115598 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2513
timestamp 1712078602
transform 1 0 116150 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2519
timestamp 1712078602
transform 1 0 116426 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2521
timestamp 1712078602
transform 1 0 116518 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2533
timestamp 1712078602
transform 1 0 117070 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2545
timestamp 1712078602
transform 1 0 117622 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2557
timestamp 1712078602
transform 1 0 118174 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2569
timestamp 1712078602
transform 1 0 118726 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2575
timestamp 1712078602
transform 1 0 119002 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2577
timestamp 1712078602
transform 1 0 119094 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2589
timestamp 1712078602
transform 1 0 119646 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2601
timestamp 1712078602
transform 1 0 120198 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2613
timestamp 1712078602
transform 1 0 120750 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2625
timestamp 1712078602
transform 1 0 121302 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2631
timestamp 1712078602
transform 1 0 121578 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2633
timestamp 1712078602
transform 1 0 121670 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2645
timestamp 1712078602
transform 1 0 122222 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2657
timestamp 1712078602
transform 1 0 122774 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2669
timestamp 1712078602
transform 1 0 123326 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2681
timestamp 1712078602
transform 1 0 123878 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2687
timestamp 1712078602
transform 1 0 124154 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2689
timestamp 1712078602
transform 1 0 124246 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2701
timestamp 1712078602
transform 1 0 124798 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2713
timestamp 1712078602
transform 1 0 125350 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2725
timestamp 1712078602
transform 1 0 125902 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2737
timestamp 1712078602
transform 1 0 126454 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2743
timestamp 1712078602
transform 1 0 126730 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2745
timestamp 1712078602
transform 1 0 126822 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2757
timestamp 1712078602
transform 1 0 127374 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2769
timestamp 1712078602
transform 1 0 127926 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2781
timestamp 1712078602
transform 1 0 128478 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2793
timestamp 1712078602
transform 1 0 129030 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2799
timestamp 1712078602
transform 1 0 129306 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2801
timestamp 1712078602
transform 1 0 129398 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2813
timestamp 1712078602
transform 1 0 129950 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2825
timestamp 1712078602
transform 1 0 130502 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2837
timestamp 1712078602
transform 1 0 131054 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2849
timestamp 1712078602
transform 1 0 131606 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2855
timestamp 1712078602
transform 1 0 131882 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2857
timestamp 1712078602
transform 1 0 131974 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2869
timestamp 1712078602
transform 1 0 132526 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2881
timestamp 1712078602
transform 1 0 133078 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2893
timestamp 1712078602
transform 1 0 133630 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__decap_8  FILLER_13_2902
timestamp 1712078602
transform 1 0 134044 0 -1 4896
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_13_2910
timestamp 1712078602
transform 1 0 134412 0 -1 4896
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2913
timestamp 1712078602
transform 1 0 134550 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2925
timestamp 1712078602
transform 1 0 135102 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2937
timestamp 1712078602
transform 1 0 135654 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2949
timestamp 1712078602
transform 1 0 136206 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_2961
timestamp 1712078602
transform 1 0 136758 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_2967
timestamp 1712078602
transform 1 0 137034 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2969
timestamp 1712078602
transform 1 0 137126 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2981
timestamp 1712078602
transform 1 0 137678 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_2993
timestamp 1712078602
transform 1 0 138230 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3005
timestamp 1712078602
transform 1 0 138782 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_3017
timestamp 1712078602
transform 1 0 139334 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_3023
timestamp 1712078602
transform 1 0 139610 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3025
timestamp 1712078602
transform 1 0 139702 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3037
timestamp 1712078602
transform 1 0 140254 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3049
timestamp 1712078602
transform 1 0 140806 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3061
timestamp 1712078602
transform 1 0 141358 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_3073
timestamp 1712078602
transform 1 0 141910 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_3079
timestamp 1712078602
transform 1 0 142186 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3081
timestamp 1712078602
transform 1 0 142278 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3093
timestamp 1712078602
transform 1 0 142830 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3105
timestamp 1712078602
transform 1 0 143382 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3117
timestamp 1712078602
transform 1 0 143934 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_3129
timestamp 1712078602
transform 1 0 144486 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_3135
timestamp 1712078602
transform 1 0 144762 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3137
timestamp 1712078602
transform 1 0 144854 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3149
timestamp 1712078602
transform 1 0 145406 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3161
timestamp 1712078602
transform 1 0 145958 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3173
timestamp 1712078602
transform 1 0 146510 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_3185
timestamp 1712078602
transform 1 0 147062 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_3191
timestamp 1712078602
transform 1 0 147338 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3193
timestamp 1712078602
transform 1 0 147430 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3205
timestamp 1712078602
transform 1 0 147982 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3217
timestamp 1712078602
transform 1 0 148534 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3229
timestamp 1712078602
transform 1 0 149086 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_3241
timestamp 1712078602
transform 1 0 149638 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_3247
timestamp 1712078602
transform 1 0 149914 0 -1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3249
timestamp 1712078602
transform 1 0 150006 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3261
timestamp 1712078602
transform 1 0 150558 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3273
timestamp 1712078602
transform 1 0 151110 0 -1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_13_3285
timestamp 1712078602
transform 1 0 151662 0 -1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_13_3297
timestamp 1712078602
transform 1 0 152214 0 -1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_13_3303
timestamp 1712078602
transform 1 0 152490 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_13_3305
timestamp 1712078602
transform 1 0 152582 0 -1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1712078602
transform 1 0 690 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1712078602
transform 1 0 1242 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1712078602
transform 1 0 1794 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1712078602
transform 1 0 1886 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1712078602
transform 1 0 2438 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1712078602
transform 1 0 2990 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1712078602
transform 1 0 3542 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1712078602
transform 1 0 4094 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1712078602
transform 1 0 4370 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1712078602
transform 1 0 4462 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1712078602
transform 1 0 5014 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1712078602
transform 1 0 5566 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1712078602
transform 1 0 6118 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1712078602
transform 1 0 6670 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1712078602
transform 1 0 6946 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1712078602
transform 1 0 7038 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1712078602
transform 1 0 7590 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1712078602
transform 1 0 8142 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1712078602
transform 1 0 8694 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1712078602
transform 1 0 9246 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1712078602
transform 1 0 9522 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1712078602
transform 1 0 9614 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1712078602
transform 1 0 10166 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1712078602
transform 1 0 10718 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1712078602
transform 1 0 11270 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1712078602
transform 1 0 11822 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1712078602
transform 1 0 12098 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1712078602
transform 1 0 12190 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1712078602
transform 1 0 12742 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1712078602
transform 1 0 13294 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1712078602
transform 1 0 13846 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1712078602
transform 1 0 14398 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1712078602
transform 1 0 14674 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1712078602
transform 1 0 14766 0 1 4896
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_14_320
timestamp 1712078602
transform 1 0 15272 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_327
timestamp 1712078602
transform 1 0 15594 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_334
timestamp 1712078602
transform 1 0 15916 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_341
timestamp 1712078602
transform 1 0 16238 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_348
timestamp 1712078602
transform 1 0 16560 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1712078602
transform 1 0 16882 0 1 4896
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1712078602
transform 1 0 17250 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1712078602
transform 1 0 17342 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1712078602
transform 1 0 17894 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1712078602
transform 1 0 18446 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1712078602
transform 1 0 18998 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1712078602
transform 1 0 19550 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1712078602
transform 1 0 19826 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1712078602
transform 1 0 19918 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1712078602
transform 1 0 20470 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1712078602
transform 1 0 21022 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1712078602
transform 1 0 21574 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1712078602
transform 1 0 22126 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1712078602
transform 1 0 22402 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1712078602
transform 1 0 22494 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1712078602
transform 1 0 23046 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1712078602
transform 1 0 23598 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1712078602
transform 1 0 24150 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1712078602
transform 1 0 24702 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1712078602
transform 1 0 24978 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1712078602
transform 1 0 25070 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1712078602
transform 1 0 25622 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1712078602
transform 1 0 26174 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1712078602
transform 1 0 26726 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1712078602
transform 1 0 27278 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1712078602
transform 1 0 27554 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1712078602
transform 1 0 27646 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1712078602
transform 1 0 28198 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1712078602
transform 1 0 28750 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1712078602
transform 1 0 29302 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1712078602
transform 1 0 29854 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1712078602
transform 1 0 30130 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1712078602
transform 1 0 30222 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1712078602
transform 1 0 30774 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1712078602
transform 1 0 31326 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1712078602
transform 1 0 31878 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1712078602
transform 1 0 32430 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1712078602
transform 1 0 32706 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1712078602
transform 1 0 32798 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1712078602
transform 1 0 33350 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1712078602
transform 1 0 33902 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1712078602
transform 1 0 34454 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1712078602
transform 1 0 35006 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1712078602
transform 1 0 35282 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1712078602
transform 1 0 35374 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1712078602
transform 1 0 35926 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1712078602
transform 1 0 36478 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1712078602
transform 1 0 37030 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1712078602
transform 1 0 37582 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1712078602
transform 1 0 37858 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_813
timestamp 1712078602
transform 1 0 37950 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_825
timestamp 1712078602
transform 1 0 38502 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_837
timestamp 1712078602
transform 1 0 39054 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_849
timestamp 1712078602
transform 1 0 39606 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1712078602
transform 1 0 40158 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1712078602
transform 1 0 40434 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_869
timestamp 1712078602
transform 1 0 40526 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_881
timestamp 1712078602
transform 1 0 41078 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_893
timestamp 1712078602
transform 1 0 41630 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_905
timestamp 1712078602
transform 1 0 42182 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1712078602
transform 1 0 42734 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1712078602
transform 1 0 43010 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_925
timestamp 1712078602
transform 1 0 43102 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_937
timestamp 1712078602
transform 1 0 43654 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_949
timestamp 1712078602
transform 1 0 44206 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_961
timestamp 1712078602
transform 1 0 44758 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_973
timestamp 1712078602
transform 1 0 45310 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1712078602
transform 1 0 45586 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_981
timestamp 1712078602
transform 1 0 45678 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_993
timestamp 1712078602
transform 1 0 46230 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1005
timestamp 1712078602
transform 1 0 46782 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1017
timestamp 1712078602
transform 1 0 47334 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1029
timestamp 1712078602
transform 1 0 47886 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1035
timestamp 1712078602
transform 1 0 48162 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1037
timestamp 1712078602
transform 1 0 48254 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1049
timestamp 1712078602
transform 1 0 48806 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1061
timestamp 1712078602
transform 1 0 49358 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1073
timestamp 1712078602
transform 1 0 49910 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1085
timestamp 1712078602
transform 1 0 50462 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1091
timestamp 1712078602
transform 1 0 50738 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1093
timestamp 1712078602
transform 1 0 50830 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1105
timestamp 1712078602
transform 1 0 51382 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1117
timestamp 1712078602
transform 1 0 51934 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1129
timestamp 1712078602
transform 1 0 52486 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1712078602
transform 1 0 53038 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1712078602
transform 1 0 53314 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1149
timestamp 1712078602
transform 1 0 53406 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1161
timestamp 1712078602
transform 1 0 53958 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1173
timestamp 1712078602
transform 1 0 54510 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1185
timestamp 1712078602
transform 1 0 55062 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1197
timestamp 1712078602
transform 1 0 55614 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1203
timestamp 1712078602
transform 1 0 55890 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1205
timestamp 1712078602
transform 1 0 55982 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1217
timestamp 1712078602
transform 1 0 56534 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1229
timestamp 1712078602
transform 1 0 57086 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1241
timestamp 1712078602
transform 1 0 57638 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1253
timestamp 1712078602
transform 1 0 58190 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1259
timestamp 1712078602
transform 1 0 58466 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1261
timestamp 1712078602
transform 1 0 58558 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1273
timestamp 1712078602
transform 1 0 59110 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1285
timestamp 1712078602
transform 1 0 59662 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1297
timestamp 1712078602
transform 1 0 60214 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1309
timestamp 1712078602
transform 1 0 60766 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1315
timestamp 1712078602
transform 1 0 61042 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1317
timestamp 1712078602
transform 1 0 61134 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1329
timestamp 1712078602
transform 1 0 61686 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1341
timestamp 1712078602
transform 1 0 62238 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1353
timestamp 1712078602
transform 1 0 62790 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1365
timestamp 1712078602
transform 1 0 63342 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1371
timestamp 1712078602
transform 1 0 63618 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1373
timestamp 1712078602
transform 1 0 63710 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1385
timestamp 1712078602
transform 1 0 64262 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1397
timestamp 1712078602
transform 1 0 64814 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1409
timestamp 1712078602
transform 1 0 65366 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1421
timestamp 1712078602
transform 1 0 65918 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1427
timestamp 1712078602
transform 1 0 66194 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1429
timestamp 1712078602
transform 1 0 66286 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1441
timestamp 1712078602
transform 1 0 66838 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1453
timestamp 1712078602
transform 1 0 67390 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1465
timestamp 1712078602
transform 1 0 67942 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1477
timestamp 1712078602
transform 1 0 68494 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1483
timestamp 1712078602
transform 1 0 68770 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1485
timestamp 1712078602
transform 1 0 68862 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1497
timestamp 1712078602
transform 1 0 69414 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_14_1509
timestamp 1712078602
transform 1 0 69966 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1513
timestamp 1712078602
transform 1 0 70150 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1534
timestamp 1712078602
transform 1 0 71116 0 1 4896
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1541
timestamp 1712078602
transform 1 0 71438 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1553
timestamp 1712078602
transform 1 0 71990 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1565
timestamp 1712078602
transform 1 0 72542 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1577
timestamp 1712078602
transform 1 0 73094 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1589
timestamp 1712078602
transform 1 0 73646 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1595
timestamp 1712078602
transform 1 0 73922 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1597
timestamp 1712078602
transform 1 0 74014 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1609
timestamp 1712078602
transform 1 0 74566 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1621
timestamp 1712078602
transform 1 0 75118 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1633
timestamp 1712078602
transform 1 0 75670 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1645
timestamp 1712078602
transform 1 0 76222 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1651
timestamp 1712078602
transform 1 0 76498 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1653
timestamp 1712078602
transform 1 0 76590 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1665
timestamp 1712078602
transform 1 0 77142 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1677
timestamp 1712078602
transform 1 0 77694 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1683
timestamp 1712078602
transform 1 0 77970 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_14_1704
timestamp 1712078602
transform 1 0 78936 0 1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1709
timestamp 1712078602
transform 1 0 79166 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1721
timestamp 1712078602
transform 1 0 79718 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1733
timestamp 1712078602
transform 1 0 80270 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1745
timestamp 1712078602
transform 1 0 80822 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1757
timestamp 1712078602
transform 1 0 81374 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1763
timestamp 1712078602
transform 1 0 81650 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1765
timestamp 1712078602
transform 1 0 81742 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1777
timestamp 1712078602
transform 1 0 82294 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1789
timestamp 1712078602
transform 1 0 82846 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1801
timestamp 1712078602
transform 1 0 83398 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1813
timestamp 1712078602
transform 1 0 83950 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1819
timestamp 1712078602
transform 1 0 84226 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1821
timestamp 1712078602
transform 1 0 84318 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1833
timestamp 1712078602
transform 1 0 84870 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1845
timestamp 1712078602
transform 1 0 85422 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1857
timestamp 1712078602
transform 1 0 85974 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1869
timestamp 1712078602
transform 1 0 86526 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1875
timestamp 1712078602
transform 1 0 86802 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1877
timestamp 1712078602
transform 1 0 86894 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1889
timestamp 1712078602
transform 1 0 87446 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1901
timestamp 1712078602
transform 1 0 87998 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1913
timestamp 1712078602
transform 1 0 88550 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1925
timestamp 1712078602
transform 1 0 89102 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1931
timestamp 1712078602
transform 1 0 89378 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1933
timestamp 1712078602
transform 1 0 89470 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1945
timestamp 1712078602
transform 1 0 90022 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1957
timestamp 1712078602
transform 1 0 90574 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1969
timestamp 1712078602
transform 1 0 91126 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_1981
timestamp 1712078602
transform 1 0 91678 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_1987
timestamp 1712078602
transform 1 0 91954 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_1989
timestamp 1712078602
transform 1 0 92046 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2001
timestamp 1712078602
transform 1 0 92598 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2013
timestamp 1712078602
transform 1 0 93150 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2025
timestamp 1712078602
transform 1 0 93702 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2037
timestamp 1712078602
transform 1 0 94254 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2043
timestamp 1712078602
transform 1 0 94530 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2045
timestamp 1712078602
transform 1 0 94622 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2057
timestamp 1712078602
transform 1 0 95174 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_14_2069
timestamp 1712078602
transform 1 0 95726 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_2076
timestamp 1712078602
transform 1 0 96048 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_2083
timestamp 1712078602
transform 1 0 96370 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_14_2090
timestamp 1712078602
transform 1 0 96692 0 1 4896
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_14_2098
timestamp 1712078602
transform 1 0 97060 0 1 4896
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2101
timestamp 1712078602
transform 1 0 97198 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2113
timestamp 1712078602
transform 1 0 97750 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2125
timestamp 1712078602
transform 1 0 98302 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2137
timestamp 1712078602
transform 1 0 98854 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2149
timestamp 1712078602
transform 1 0 99406 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2155
timestamp 1712078602
transform 1 0 99682 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2157
timestamp 1712078602
transform 1 0 99774 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2169
timestamp 1712078602
transform 1 0 100326 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2181
timestamp 1712078602
transform 1 0 100878 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2193
timestamp 1712078602
transform 1 0 101430 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2205
timestamp 1712078602
transform 1 0 101982 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2211
timestamp 1712078602
transform 1 0 102258 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2213
timestamp 1712078602
transform 1 0 102350 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2225
timestamp 1712078602
transform 1 0 102902 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2237
timestamp 1712078602
transform 1 0 103454 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2249
timestamp 1712078602
transform 1 0 104006 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2261
timestamp 1712078602
transform 1 0 104558 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2267
timestamp 1712078602
transform 1 0 104834 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2269
timestamp 1712078602
transform 1 0 104926 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2281
timestamp 1712078602
transform 1 0 105478 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2293
timestamp 1712078602
transform 1 0 106030 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2305
timestamp 1712078602
transform 1 0 106582 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2317
timestamp 1712078602
transform 1 0 107134 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2323
timestamp 1712078602
transform 1 0 107410 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2325
timestamp 1712078602
transform 1 0 107502 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2337
timestamp 1712078602
transform 1 0 108054 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2349
timestamp 1712078602
transform 1 0 108606 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2361
timestamp 1712078602
transform 1 0 109158 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2373
timestamp 1712078602
transform 1 0 109710 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2379
timestamp 1712078602
transform 1 0 109986 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2381
timestamp 1712078602
transform 1 0 110078 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2393
timestamp 1712078602
transform 1 0 110630 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2405
timestamp 1712078602
transform 1 0 111182 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2417
timestamp 1712078602
transform 1 0 111734 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2429
timestamp 1712078602
transform 1 0 112286 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2435
timestamp 1712078602
transform 1 0 112562 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2437
timestamp 1712078602
transform 1 0 112654 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2449
timestamp 1712078602
transform 1 0 113206 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2461
timestamp 1712078602
transform 1 0 113758 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2473
timestamp 1712078602
transform 1 0 114310 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2485
timestamp 1712078602
transform 1 0 114862 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2491
timestamp 1712078602
transform 1 0 115138 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2493
timestamp 1712078602
transform 1 0 115230 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2505
timestamp 1712078602
transform 1 0 115782 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2517
timestamp 1712078602
transform 1 0 116334 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2529
timestamp 1712078602
transform 1 0 116886 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2541
timestamp 1712078602
transform 1 0 117438 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2547
timestamp 1712078602
transform 1 0 117714 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2549
timestamp 1712078602
transform 1 0 117806 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2561
timestamp 1712078602
transform 1 0 118358 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2573
timestamp 1712078602
transform 1 0 118910 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2585
timestamp 1712078602
transform 1 0 119462 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2597
timestamp 1712078602
transform 1 0 120014 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2603
timestamp 1712078602
transform 1 0 120290 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2605
timestamp 1712078602
transform 1 0 120382 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2617
timestamp 1712078602
transform 1 0 120934 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2629
timestamp 1712078602
transform 1 0 121486 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2641
timestamp 1712078602
transform 1 0 122038 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2653
timestamp 1712078602
transform 1 0 122590 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2659
timestamp 1712078602
transform 1 0 122866 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2661
timestamp 1712078602
transform 1 0 122958 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2673
timestamp 1712078602
transform 1 0 123510 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2685
timestamp 1712078602
transform 1 0 124062 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2697
timestamp 1712078602
transform 1 0 124614 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2709
timestamp 1712078602
transform 1 0 125166 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2715
timestamp 1712078602
transform 1 0 125442 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2717
timestamp 1712078602
transform 1 0 125534 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2729
timestamp 1712078602
transform 1 0 126086 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2741
timestamp 1712078602
transform 1 0 126638 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2753
timestamp 1712078602
transform 1 0 127190 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2765
timestamp 1712078602
transform 1 0 127742 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2771
timestamp 1712078602
transform 1 0 128018 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2773
timestamp 1712078602
transform 1 0 128110 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2785
timestamp 1712078602
transform 1 0 128662 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2797
timestamp 1712078602
transform 1 0 129214 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2809
timestamp 1712078602
transform 1 0 129766 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2821
timestamp 1712078602
transform 1 0 130318 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2827
timestamp 1712078602
transform 1 0 130594 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2829
timestamp 1712078602
transform 1 0 130686 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2841
timestamp 1712078602
transform 1 0 131238 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2853
timestamp 1712078602
transform 1 0 131790 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2865
timestamp 1712078602
transform 1 0 132342 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2877
timestamp 1712078602
transform 1 0 132894 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2883
timestamp 1712078602
transform 1 0 133170 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2885
timestamp 1712078602
transform 1 0 133262 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_14_2894
timestamp 1712078602
transform 1 0 133676 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_2901
timestamp 1712078602
transform 1 0 133998 0 1 4896
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_14_2908
timestamp 1712078602
transform 1 0 134320 0 1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2915
timestamp 1712078602
transform 1 0 134642 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2927
timestamp 1712078602
transform 1 0 135194 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2939
timestamp 1712078602
transform 1 0 135746 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2941
timestamp 1712078602
transform 1 0 135838 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2953
timestamp 1712078602
transform 1 0 136390 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2965
timestamp 1712078602
transform 1 0 136942 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2977
timestamp 1712078602
transform 1 0 137494 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_2989
timestamp 1712078602
transform 1 0 138046 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_2995
timestamp 1712078602
transform 1 0 138322 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_2997
timestamp 1712078602
transform 1 0 138414 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3009
timestamp 1712078602
transform 1 0 138966 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3021
timestamp 1712078602
transform 1 0 139518 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3033
timestamp 1712078602
transform 1 0 140070 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_3045
timestamp 1712078602
transform 1 0 140622 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_3051
timestamp 1712078602
transform 1 0 140898 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3053
timestamp 1712078602
transform 1 0 140990 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3065
timestamp 1712078602
transform 1 0 141542 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3077
timestamp 1712078602
transform 1 0 142094 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3089
timestamp 1712078602
transform 1 0 142646 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_3101
timestamp 1712078602
transform 1 0 143198 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_3107
timestamp 1712078602
transform 1 0 143474 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3109
timestamp 1712078602
transform 1 0 143566 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3121
timestamp 1712078602
transform 1 0 144118 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3133
timestamp 1712078602
transform 1 0 144670 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3145
timestamp 1712078602
transform 1 0 145222 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_3157
timestamp 1712078602
transform 1 0 145774 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_3163
timestamp 1712078602
transform 1 0 146050 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3165
timestamp 1712078602
transform 1 0 146142 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3177
timestamp 1712078602
transform 1 0 146694 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3189
timestamp 1712078602
transform 1 0 147246 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3201
timestamp 1712078602
transform 1 0 147798 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_3213
timestamp 1712078602
transform 1 0 148350 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_3219
timestamp 1712078602
transform 1 0 148626 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3221
timestamp 1712078602
transform 1 0 148718 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3233
timestamp 1712078602
transform 1 0 149270 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3245
timestamp 1712078602
transform 1 0 149822 0 1 4896
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3257
timestamp 1712078602
transform 1 0 150374 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_3269
timestamp 1712078602
transform 1 0 150926 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_3275
timestamp 1712078602
transform 1 0 151202 0 1 4896
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_14_3277
timestamp 1712078602
transform 1 0 151294 0 1 4896
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_14_3289
timestamp 1712078602
transform 1 0 151846 0 1 4896
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_14_3295
timestamp 1712078602
transform 1 0 152122 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_14_3305
timestamp 1712078602
transform 1 0 152582 0 1 4896
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1712078602
transform 1 0 690 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1712078602
transform 1 0 1242 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1712078602
transform 1 0 1794 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1712078602
transform 1 0 2346 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1712078602
transform 1 0 2898 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1712078602
transform 1 0 3082 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1712078602
transform 1 0 3174 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1712078602
transform 1 0 3726 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1712078602
transform 1 0 4278 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1712078602
transform 1 0 4830 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1712078602
transform 1 0 5382 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1712078602
transform 1 0 5658 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1712078602
transform 1 0 5750 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1712078602
transform 1 0 6302 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1712078602
transform 1 0 6854 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1712078602
transform 1 0 7406 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1712078602
transform 1 0 7958 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1712078602
transform 1 0 8234 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1712078602
transform 1 0 8326 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1712078602
transform 1 0 8878 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1712078602
transform 1 0 9430 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1712078602
transform 1 0 9982 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1712078602
transform 1 0 10534 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1712078602
transform 1 0 10810 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1712078602
transform 1 0 10902 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1712078602
transform 1 0 11454 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1712078602
transform 1 0 12006 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1712078602
transform 1 0 12558 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1712078602
transform 1 0 13110 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1712078602
transform 1 0 13386 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1712078602
transform 1 0 13478 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1712078602
transform 1 0 14030 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1712078602
transform 1 0 14582 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_15_309
timestamp 1712078602
transform 1 0 14766 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_15_313
timestamp 1712078602
transform 1 0 14950 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1712078602
transform 1 0 15548 0 -1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1712078602
transform 1 0 15916 0 -1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_15_340
timestamp 1712078602
transform 1 0 16192 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_15_347
timestamp 1712078602
transform 1 0 16514 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_354
timestamp 1712078602
transform 1 0 16836 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_366
timestamp 1712078602
transform 1 0 17388 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_378
timestamp 1712078602
transform 1 0 17940 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1712078602
transform 1 0 18492 0 -1 5440
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1712078602
transform 1 0 18630 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1712078602
transform 1 0 19182 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1712078602
transform 1 0 19734 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1712078602
transform 1 0 20286 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1712078602
transform 1 0 20838 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1712078602
transform 1 0 21114 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1712078602
transform 1 0 21206 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1712078602
transform 1 0 21758 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1712078602
transform 1 0 22310 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1712078602
transform 1 0 22862 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1712078602
transform 1 0 23414 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1712078602
transform 1 0 23690 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1712078602
transform 1 0 23782 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1712078602
transform 1 0 24334 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1712078602
transform 1 0 24886 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1712078602
transform 1 0 25438 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1712078602
transform 1 0 25990 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1712078602
transform 1 0 26266 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1712078602
transform 1 0 26358 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1712078602
transform 1 0 26910 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1712078602
transform 1 0 27462 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1712078602
transform 1 0 28014 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1712078602
transform 1 0 28566 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1712078602
transform 1 0 28842 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1712078602
transform 1 0 28934 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1712078602
transform 1 0 29486 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1712078602
transform 1 0 30038 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1712078602
transform 1 0 30590 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1712078602
transform 1 0 31142 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1712078602
transform 1 0 31418 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1712078602
transform 1 0 31510 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1712078602
transform 1 0 32062 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1712078602
transform 1 0 32614 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1712078602
transform 1 0 33166 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1712078602
transform 1 0 33718 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1712078602
transform 1 0 33994 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1712078602
transform 1 0 34086 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1712078602
transform 1 0 34638 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1712078602
transform 1 0 35190 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1712078602
transform 1 0 35742 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1712078602
transform 1 0 36294 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1712078602
transform 1 0 36570 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1712078602
transform 1 0 36662 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1712078602
transform 1 0 37214 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1712078602
transform 1 0 37766 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_821
timestamp 1712078602
transform 1 0 38318 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1712078602
transform 1 0 38870 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1712078602
transform 1 0 39146 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_841
timestamp 1712078602
transform 1 0 39238 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_853
timestamp 1712078602
transform 1 0 39790 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_865
timestamp 1712078602
transform 1 0 40342 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_877
timestamp 1712078602
transform 1 0 40894 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1712078602
transform 1 0 41446 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1712078602
transform 1 0 41722 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1712078602
transform 1 0 41814 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_909
timestamp 1712078602
transform 1 0 42366 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_921
timestamp 1712078602
transform 1 0 42918 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_933
timestamp 1712078602
transform 1 0 43470 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_945
timestamp 1712078602
transform 1 0 44022 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_951
timestamp 1712078602
transform 1 0 44298 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_953
timestamp 1712078602
transform 1 0 44390 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_965
timestamp 1712078602
transform 1 0 44942 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_977
timestamp 1712078602
transform 1 0 45494 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_989
timestamp 1712078602
transform 1 0 46046 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1001
timestamp 1712078602
transform 1 0 46598 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1712078602
transform 1 0 46874 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1009
timestamp 1712078602
transform 1 0 46966 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1021
timestamp 1712078602
transform 1 0 47518 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1033
timestamp 1712078602
transform 1 0 48070 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1045
timestamp 1712078602
transform 1 0 48622 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1057
timestamp 1712078602
transform 1 0 49174 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1063
timestamp 1712078602
transform 1 0 49450 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1065
timestamp 1712078602
transform 1 0 49542 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1077
timestamp 1712078602
transform 1 0 50094 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_15_1089
timestamp 1712078602
transform 1 0 50646 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1096
timestamp 1712078602
transform 1 0 50968 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1108
timestamp 1712078602
transform 1 0 51520 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1121
timestamp 1712078602
transform 1 0 52118 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1133
timestamp 1712078602
transform 1 0 52670 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1145
timestamp 1712078602
transform 1 0 53222 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1157
timestamp 1712078602
transform 1 0 53774 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1169
timestamp 1712078602
transform 1 0 54326 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1175
timestamp 1712078602
transform 1 0 54602 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1177
timestamp 1712078602
transform 1 0 54694 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1189
timestamp 1712078602
transform 1 0 55246 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1201
timestamp 1712078602
transform 1 0 55798 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1213
timestamp 1712078602
transform 1 0 56350 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1225
timestamp 1712078602
transform 1 0 56902 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1231
timestamp 1712078602
transform 1 0 57178 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1233
timestamp 1712078602
transform 1 0 57270 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1245
timestamp 1712078602
transform 1 0 57822 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1257
timestamp 1712078602
transform 1 0 58374 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1269
timestamp 1712078602
transform 1 0 58926 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1281
timestamp 1712078602
transform 1 0 59478 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1287
timestamp 1712078602
transform 1 0 59754 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1289
timestamp 1712078602
transform 1 0 59846 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1301
timestamp 1712078602
transform 1 0 60398 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1313
timestamp 1712078602
transform 1 0 60950 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1325
timestamp 1712078602
transform 1 0 61502 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1337
timestamp 1712078602
transform 1 0 62054 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1343
timestamp 1712078602
transform 1 0 62330 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1345
timestamp 1712078602
transform 1 0 62422 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1357
timestamp 1712078602
transform 1 0 62974 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1369
timestamp 1712078602
transform 1 0 63526 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1381
timestamp 1712078602
transform 1 0 64078 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1393
timestamp 1712078602
transform 1 0 64630 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1399
timestamp 1712078602
transform 1 0 64906 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_15_1401
timestamp 1712078602
transform 1 0 64998 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1408
timestamp 1712078602
transform 1 0 65320 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1420
timestamp 1712078602
transform 1 0 65872 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1432
timestamp 1712078602
transform 1 0 66424 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1444
timestamp 1712078602
transform 1 0 66976 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1457
timestamp 1712078602
transform 1 0 67574 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1469
timestamp 1712078602
transform 1 0 68126 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1481
timestamp 1712078602
transform 1 0 68678 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1493
timestamp 1712078602
transform 1 0 69230 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1505
timestamp 1712078602
transform 1 0 69782 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1511
timestamp 1712078602
transform 1 0 70058 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_15_1513
timestamp 1712078602
transform 1 0 70150 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1537
timestamp 1712078602
transform 1 0 71254 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1549
timestamp 1712078602
transform 1 0 71806 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1561
timestamp 1712078602
transform 1 0 72358 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1567
timestamp 1712078602
transform 1 0 72634 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1569
timestamp 1712078602
transform 1 0 72726 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1581
timestamp 1712078602
transform 1 0 73278 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1593
timestamp 1712078602
transform 1 0 73830 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1605
timestamp 1712078602
transform 1 0 74382 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1609
timestamp 1712078602
transform 1 0 74566 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_15_1621
timestamp 1712078602
transform 1 0 75118 0 -1 5440
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1628
timestamp 1712078602
transform 1 0 75440 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1640
timestamp 1712078602
transform 1 0 75992 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1652
timestamp 1712078602
transform 1 0 76544 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1664
timestamp 1712078602
transform 1 0 77096 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_15_1676
timestamp 1712078602
transform 1 0 77648 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_15_1681
timestamp 1712078602
transform 1 0 77878 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1705
timestamp 1712078602
transform 1 0 78982 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1717
timestamp 1712078602
transform 1 0 79534 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1729
timestamp 1712078602
transform 1 0 80086 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1735
timestamp 1712078602
transform 1 0 80362 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1737
timestamp 1712078602
transform 1 0 80454 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1749
timestamp 1712078602
transform 1 0 81006 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1761
timestamp 1712078602
transform 1 0 81558 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1773
timestamp 1712078602
transform 1 0 82110 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1785
timestamp 1712078602
transform 1 0 82662 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1791
timestamp 1712078602
transform 1 0 82938 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1793
timestamp 1712078602
transform 1 0 83030 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1805
timestamp 1712078602
transform 1 0 83582 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1817
timestamp 1712078602
transform 1 0 84134 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1829
timestamp 1712078602
transform 1 0 84686 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1841
timestamp 1712078602
transform 1 0 85238 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1847
timestamp 1712078602
transform 1 0 85514 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1849
timestamp 1712078602
transform 1 0 85606 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1861
timestamp 1712078602
transform 1 0 86158 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1873
timestamp 1712078602
transform 1 0 86710 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1885
timestamp 1712078602
transform 1 0 87262 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1897
timestamp 1712078602
transform 1 0 87814 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1903
timestamp 1712078602
transform 1 0 88090 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1905
timestamp 1712078602
transform 1 0 88182 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1917
timestamp 1712078602
transform 1 0 88734 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1929
timestamp 1712078602
transform 1 0 89286 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1941
timestamp 1712078602
transform 1 0 89838 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_1953
timestamp 1712078602
transform 1 0 90390 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_1959
timestamp 1712078602
transform 1 0 90666 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1961
timestamp 1712078602
transform 1 0 90758 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1973
timestamp 1712078602
transform 1 0 91310 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1985
timestamp 1712078602
transform 1 0 91862 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_1997
timestamp 1712078602
transform 1 0 92414 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2009
timestamp 1712078602
transform 1 0 92966 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2015
timestamp 1712078602
transform 1 0 93242 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2017
timestamp 1712078602
transform 1 0 93334 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2021
timestamp 1712078602
transform 1 0 93518 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2031
timestamp 1712078602
transform 1 0 93978 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2043
timestamp 1712078602
transform 1 0 94530 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_15_2055
timestamp 1712078602
transform 1 0 95082 0 -1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_15_2063
timestamp 1712078602
transform 1 0 95450 0 -1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2068
timestamp 1712078602
transform 1 0 95680 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2076
timestamp 1712078602
transform 1 0 96048 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2086
timestamp 1712078602
transform 1 0 96508 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2094
timestamp 1712078602
transform 1 0 96876 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2101
timestamp 1712078602
transform 1 0 97198 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2113
timestamp 1712078602
transform 1 0 97750 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_15_2125
timestamp 1712078602
transform 1 0 98302 0 -1 5440
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2129
timestamp 1712078602
transform 1 0 98486 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2141
timestamp 1712078602
transform 1 0 99038 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2153
timestamp 1712078602
transform 1 0 99590 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2165
timestamp 1712078602
transform 1 0 100142 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2177
timestamp 1712078602
transform 1 0 100694 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2183
timestamp 1712078602
transform 1 0 100970 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_15_2185
timestamp 1712078602
transform 1 0 101062 0 -1 5440
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2196
timestamp 1712078602
transform 1 0 101568 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2208
timestamp 1712078602
transform 1 0 102120 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2220
timestamp 1712078602
transform 1 0 102672 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_15_2232
timestamp 1712078602
transform 1 0 103224 0 -1 5440
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2241
timestamp 1712078602
transform 1 0 103638 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2253
timestamp 1712078602
transform 1 0 104190 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2265
timestamp 1712078602
transform 1 0 104742 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2277
timestamp 1712078602
transform 1 0 105294 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2289
timestamp 1712078602
transform 1 0 105846 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2295
timestamp 1712078602
transform 1 0 106122 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2297
timestamp 1712078602
transform 1 0 106214 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2309
timestamp 1712078602
transform 1 0 106766 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2321
timestamp 1712078602
transform 1 0 107318 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2333
timestamp 1712078602
transform 1 0 107870 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2345
timestamp 1712078602
transform 1 0 108422 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2351
timestamp 1712078602
transform 1 0 108698 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2353
timestamp 1712078602
transform 1 0 108790 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2365
timestamp 1712078602
transform 1 0 109342 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2377
timestamp 1712078602
transform 1 0 109894 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2389
timestamp 1712078602
transform 1 0 110446 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2401
timestamp 1712078602
transform 1 0 110998 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2407
timestamp 1712078602
transform 1 0 111274 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2409
timestamp 1712078602
transform 1 0 111366 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2421
timestamp 1712078602
transform 1 0 111918 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2433
timestamp 1712078602
transform 1 0 112470 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2445
timestamp 1712078602
transform 1 0 113022 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2457
timestamp 1712078602
transform 1 0 113574 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2463
timestamp 1712078602
transform 1 0 113850 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2465
timestamp 1712078602
transform 1 0 113942 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2477
timestamp 1712078602
transform 1 0 114494 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2489
timestamp 1712078602
transform 1 0 115046 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2501
timestamp 1712078602
transform 1 0 115598 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2513
timestamp 1712078602
transform 1 0 116150 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2519
timestamp 1712078602
transform 1 0 116426 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2521
timestamp 1712078602
transform 1 0 116518 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2533
timestamp 1712078602
transform 1 0 117070 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2545
timestamp 1712078602
transform 1 0 117622 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2557
timestamp 1712078602
transform 1 0 118174 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2569
timestamp 1712078602
transform 1 0 118726 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2575
timestamp 1712078602
transform 1 0 119002 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2577
timestamp 1712078602
transform 1 0 119094 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2589
timestamp 1712078602
transform 1 0 119646 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2601
timestamp 1712078602
transform 1 0 120198 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2613
timestamp 1712078602
transform 1 0 120750 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2625
timestamp 1712078602
transform 1 0 121302 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2631
timestamp 1712078602
transform 1 0 121578 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2633
timestamp 1712078602
transform 1 0 121670 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2645
timestamp 1712078602
transform 1 0 122222 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2657
timestamp 1712078602
transform 1 0 122774 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2669
timestamp 1712078602
transform 1 0 123326 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2681
timestamp 1712078602
transform 1 0 123878 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2687
timestamp 1712078602
transform 1 0 124154 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2689
timestamp 1712078602
transform 1 0 124246 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2701
timestamp 1712078602
transform 1 0 124798 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2713
timestamp 1712078602
transform 1 0 125350 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2725
timestamp 1712078602
transform 1 0 125902 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2737
timestamp 1712078602
transform 1 0 126454 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2743
timestamp 1712078602
transform 1 0 126730 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2748
timestamp 1712078602
transform 1 0 126960 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2760
timestamp 1712078602
transform 1 0 127512 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2772
timestamp 1712078602
transform 1 0 128064 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2784
timestamp 1712078602
transform 1 0 128616 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2796
timestamp 1712078602
transform 1 0 129168 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2801
timestamp 1712078602
transform 1 0 129398 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2813
timestamp 1712078602
transform 1 0 129950 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2825
timestamp 1712078602
transform 1 0 130502 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2837
timestamp 1712078602
transform 1 0 131054 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_2849
timestamp 1712078602
transform 1 0 131606 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_2855
timestamp 1712078602
transform 1 0 131882 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2857
timestamp 1712078602
transform 1 0 131974 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_15_2869
timestamp 1712078602
transform 1 0 132526 0 -1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2880
timestamp 1712078602
transform 1 0 133032 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2887
timestamp 1712078602
transform 1 0 133354 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2894
timestamp 1712078602
transform 1 0 133676 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2901
timestamp 1712078602
transform 1 0 133998 0 -1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2908
timestamp 1712078602
transform 1 0 134320 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2916
timestamp 1712078602
transform 1 0 134688 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2928
timestamp 1712078602
transform 1 0 135240 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2940
timestamp 1712078602
transform 1 0 135792 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2952
timestamp 1712078602
transform 1 0 136344 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_15_2964
timestamp 1712078602
transform 1 0 136896 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2969
timestamp 1712078602
transform 1 0 137126 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2981
timestamp 1712078602
transform 1 0 137678 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_2993
timestamp 1712078602
transform 1 0 138230 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3005
timestamp 1712078602
transform 1 0 138782 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_3017
timestamp 1712078602
transform 1 0 139334 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_3023
timestamp 1712078602
transform 1 0 139610 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3025
timestamp 1712078602
transform 1 0 139702 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3037
timestamp 1712078602
transform 1 0 140254 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3049
timestamp 1712078602
transform 1 0 140806 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3061
timestamp 1712078602
transform 1 0 141358 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_3073
timestamp 1712078602
transform 1 0 141910 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_3079
timestamp 1712078602
transform 1 0 142186 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3081
timestamp 1712078602
transform 1 0 142278 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3093
timestamp 1712078602
transform 1 0 142830 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3105
timestamp 1712078602
transform 1 0 143382 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3117
timestamp 1712078602
transform 1 0 143934 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_3129
timestamp 1712078602
transform 1 0 144486 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_3135
timestamp 1712078602
transform 1 0 144762 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3137
timestamp 1712078602
transform 1 0 144854 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3149
timestamp 1712078602
transform 1 0 145406 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3161
timestamp 1712078602
transform 1 0 145958 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3173
timestamp 1712078602
transform 1 0 146510 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_3185
timestamp 1712078602
transform 1 0 147062 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_3191
timestamp 1712078602
transform 1 0 147338 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3193
timestamp 1712078602
transform 1 0 147430 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3205
timestamp 1712078602
transform 1 0 147982 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3217
timestamp 1712078602
transform 1 0 148534 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3229
timestamp 1712078602
transform 1 0 149086 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_3241
timestamp 1712078602
transform 1 0 149638 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_3247
timestamp 1712078602
transform 1 0 149914 0 -1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3249
timestamp 1712078602
transform 1 0 150006 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3261
timestamp 1712078602
transform 1 0 150558 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3273
timestamp 1712078602
transform 1 0 151110 0 -1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_15_3285
timestamp 1712078602
transform 1 0 151662 0 -1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_15_3297
timestamp 1712078602
transform 1 0 152214 0 -1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_15_3303
timestamp 1712078602
transform 1 0 152490 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_15_3305
timestamp 1712078602
transform 1 0 152582 0 -1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1712078602
transform 1 0 690 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1712078602
transform 1 0 1242 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1712078602
transform 1 0 1794 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1712078602
transform 1 0 1886 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1712078602
transform 1 0 2438 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1712078602
transform 1 0 2990 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1712078602
transform 1 0 3542 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1712078602
transform 1 0 4094 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1712078602
transform 1 0 4370 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1712078602
transform 1 0 4462 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1712078602
transform 1 0 5014 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1712078602
transform 1 0 5566 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1712078602
transform 1 0 6118 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1712078602
transform 1 0 6670 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1712078602
transform 1 0 6946 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1712078602
transform 1 0 7038 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1712078602
transform 1 0 7590 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1712078602
transform 1 0 8142 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1712078602
transform 1 0 8694 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1712078602
transform 1 0 9246 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1712078602
transform 1 0 9522 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1712078602
transform 1 0 9614 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1712078602
transform 1 0 10166 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1712078602
transform 1 0 10718 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1712078602
transform 1 0 11270 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1712078602
transform 1 0 11822 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1712078602
transform 1 0 12098 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1712078602
transform 1 0 12190 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1712078602
transform 1 0 12742 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1712078602
transform 1 0 13294 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1712078602
transform 1 0 13846 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1712078602
transform 1 0 14536 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_309
timestamp 1712078602
transform 1 0 14766 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_330
timestamp 1712078602
transform 1 0 15732 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_16_343
timestamp 1712078602
transform 1 0 16330 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_16_351
timestamp 1712078602
transform 1 0 16698 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 1712078602
transform 1 0 16882 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1712078602
transform 1 0 17250 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1712078602
transform 1 0 17342 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1712078602
transform 1 0 17894 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1712078602
transform 1 0 18446 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1712078602
transform 1 0 18998 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1712078602
transform 1 0 19550 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1712078602
transform 1 0 19826 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_421
timestamp 1712078602
transform 1 0 19918 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_425
timestamp 1712078602
transform 1 0 20102 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1712078602
transform 1 0 20286 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_436
timestamp 1712078602
transform 1 0 20608 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_443
timestamp 1712078602
transform 1 0 20930 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_450
timestamp 1712078602
transform 1 0 21252 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_462
timestamp 1712078602
transform 1 0 21804 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1712078602
transform 1 0 22356 0 1 5440
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1712078602
transform 1 0 22494 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1712078602
transform 1 0 23046 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1712078602
transform 1 0 23598 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1712078602
transform 1 0 24150 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1712078602
transform 1 0 24702 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1712078602
transform 1 0 24978 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1712078602
transform 1 0 25070 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1712078602
transform 1 0 25622 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1712078602
transform 1 0 26174 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1712078602
transform 1 0 26726 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1712078602
transform 1 0 27278 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1712078602
transform 1 0 27554 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_16_592
timestamp 1712078602
transform 1 0 27784 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_598
timestamp 1712078602
transform 1 0 28060 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_602
timestamp 1712078602
transform 1 0 28244 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_614
timestamp 1712078602
transform 1 0 28796 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_626
timestamp 1712078602
transform 1 0 29348 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_638
timestamp 1712078602
transform 1 0 29900 0 1 5440
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1712078602
transform 1 0 30222 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1712078602
transform 1 0 30774 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1712078602
transform 1 0 31326 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1712078602
transform 1 0 31878 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1712078602
transform 1 0 32430 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1712078602
transform 1 0 32706 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1712078602
transform 1 0 32798 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1712078602
transform 1 0 33350 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1712078602
transform 1 0 33902 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1712078602
transform 1 0 34454 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1712078602
transform 1 0 35006 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1712078602
transform 1 0 35282 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1712078602
transform 1 0 35374 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1712078602
transform 1 0 35926 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1712078602
transform 1 0 36478 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1712078602
transform 1 0 37030 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1712078602
transform 1 0 37582 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1712078602
transform 1 0 37858 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_16_813
timestamp 1712078602
transform 1 0 37950 0 1 5440
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_16_822
timestamp 1712078602
transform 1 0 38364 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_834
timestamp 1712078602
transform 1 0 38916 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_841
timestamp 1712078602
transform 1 0 39238 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_853
timestamp 1712078602
transform 1 0 39790 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_16_865
timestamp 1712078602
transform 1 0 40342 0 1 5440
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_16_869
timestamp 1712078602
transform 1 0 40526 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_881
timestamp 1712078602
transform 1 0 41078 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_893
timestamp 1712078602
transform 1 0 41630 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_905
timestamp 1712078602
transform 1 0 42182 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1712078602
transform 1 0 42734 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1712078602
transform 1 0 43010 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_928
timestamp 1712078602
transform 1 0 43240 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_935
timestamp 1712078602
transform 1 0 43562 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_939
timestamp 1712078602
transform 1 0 43746 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_943
timestamp 1712078602
transform 1 0 43930 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_950
timestamp 1712078602
transform 1 0 44252 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_962
timestamp 1712078602
transform 1 0 44804 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_974
timestamp 1712078602
transform 1 0 45356 0 1 5440
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_16_981
timestamp 1712078602
transform 1 0 45678 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_993
timestamp 1712078602
transform 1 0 46230 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1005
timestamp 1712078602
transform 1 0 46782 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1017
timestamp 1712078602
transform 1 0 47334 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1029
timestamp 1712078602
transform 1 0 47886 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1035
timestamp 1712078602
transform 1 0 48162 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1037
timestamp 1712078602
transform 1 0 48254 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1049
timestamp 1712078602
transform 1 0 48806 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1061
timestamp 1712078602
transform 1 0 49358 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1073
timestamp 1712078602
transform 1 0 49910 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1085
timestamp 1712078602
transform 1 0 50462 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1712078602
transform 1 0 50738 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1093
timestamp 1712078602
transform 1 0 50830 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1101
timestamp 1712078602
transform 1 0 51198 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1105
timestamp 1712078602
transform 1 0 51382 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1109
timestamp 1712078602
transform 1 0 51566 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1116
timestamp 1712078602
transform 1 0 51888 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1128
timestamp 1712078602
transform 1 0 52440 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_16_1140
timestamp 1712078602
transform 1 0 52992 0 1 5440
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1149
timestamp 1712078602
transform 1 0 53406 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1161
timestamp 1712078602
transform 1 0 53958 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1173
timestamp 1712078602
transform 1 0 54510 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1185
timestamp 1712078602
transform 1 0 55062 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1197
timestamp 1712078602
transform 1 0 55614 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1203
timestamp 1712078602
transform 1 0 55890 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1205
timestamp 1712078602
transform 1 0 55982 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1217
timestamp 1712078602
transform 1 0 56534 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1229
timestamp 1712078602
transform 1 0 57086 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1244
timestamp 1712078602
transform 1 0 57776 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1248
timestamp 1712078602
transform 1 0 57960 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_16_1252
timestamp 1712078602
transform 1 0 58144 0 1 5440
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1264
timestamp 1712078602
transform 1 0 58696 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1276
timestamp 1712078602
transform 1 0 59248 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1288
timestamp 1712078602
transform 1 0 59800 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1300
timestamp 1712078602
transform 1 0 60352 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1312
timestamp 1712078602
transform 1 0 60904 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1317
timestamp 1712078602
transform 1 0 61134 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1329
timestamp 1712078602
transform 1 0 61686 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1341
timestamp 1712078602
transform 1 0 62238 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1353
timestamp 1712078602
transform 1 0 62790 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1365
timestamp 1712078602
transform 1 0 63342 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1371
timestamp 1712078602
transform 1 0 63618 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1373
timestamp 1712078602
transform 1 0 63710 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1385
timestamp 1712078602
transform 1 0 64262 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_16_1397
timestamp 1712078602
transform 1 0 64814 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1405
timestamp 1712078602
transform 1 0 65182 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1409
timestamp 1712078602
transform 1 0 65366 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1416
timestamp 1712078602
transform 1 0 65688 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1423
timestamp 1712078602
transform 1 0 66010 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1427
timestamp 1712078602
transform 1 0 66194 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1429
timestamp 1712078602
transform 1 0 66286 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1441
timestamp 1712078602
transform 1 0 66838 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1453
timestamp 1712078602
transform 1 0 67390 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1465
timestamp 1712078602
transform 1 0 67942 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1477
timestamp 1712078602
transform 1 0 68494 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1483
timestamp 1712078602
transform 1 0 68770 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1485
timestamp 1712078602
transform 1 0 68862 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1497
timestamp 1712078602
transform 1 0 69414 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1509
timestamp 1712078602
transform 1 0 69966 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1513
timestamp 1712078602
transform 1 0 70150 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1534
timestamp 1712078602
transform 1 0 71116 0 1 5440
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1541
timestamp 1712078602
transform 1 0 71438 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1553
timestamp 1712078602
transform 1 0 71990 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1565
timestamp 1712078602
transform 1 0 72542 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1577
timestamp 1712078602
transform 1 0 73094 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1589
timestamp 1712078602
transform 1 0 73646 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1595
timestamp 1712078602
transform 1 0 73922 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1606
timestamp 1712078602
transform 1 0 74428 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1612
timestamp 1712078602
transform 1 0 74704 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_16_1619
timestamp 1712078602
transform 1 0 75026 0 1 5440
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1630
timestamp 1712078602
transform 1 0 75532 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_16_1642
timestamp 1712078602
transform 1 0 76084 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_16_1650
timestamp 1712078602
transform 1 0 76452 0 1 5440
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1653
timestamp 1712078602
transform 1 0 76590 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1665
timestamp 1712078602
transform 1 0 77142 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1677
timestamp 1712078602
transform 1 0 77694 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1683
timestamp 1712078602
transform 1 0 77970 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1704
timestamp 1712078602
transform 1 0 78936 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1709
timestamp 1712078602
transform 1 0 79166 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1721
timestamp 1712078602
transform 1 0 79718 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1733
timestamp 1712078602
transform 1 0 80270 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1745
timestamp 1712078602
transform 1 0 80822 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1752
timestamp 1712078602
transform 1 0 81144 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1759
timestamp 1712078602
transform 1 0 81466 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1763
timestamp 1712078602
transform 1 0 81650 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1768
timestamp 1712078602
transform 1 0 81880 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1780
timestamp 1712078602
transform 1 0 82432 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1792
timestamp 1712078602
transform 1 0 82984 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1804
timestamp 1712078602
transform 1 0 83536 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1816
timestamp 1712078602
transform 1 0 84088 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1821
timestamp 1712078602
transform 1 0 84318 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1833
timestamp 1712078602
transform 1 0 84870 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1845
timestamp 1712078602
transform 1 0 85422 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1857
timestamp 1712078602
transform 1 0 85974 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_1869
timestamp 1712078602
transform 1 0 86526 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1875
timestamp 1712078602
transform 1 0 86802 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1877
timestamp 1712078602
transform 1 0 86894 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1889
timestamp 1712078602
transform 1 0 87446 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1901
timestamp 1712078602
transform 1 0 87998 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1913
timestamp 1712078602
transform 1 0 88550 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1920
timestamp 1712078602
transform 1 0 88872 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1927
timestamp 1712078602
transform 1 0 89194 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_1931
timestamp 1712078602
transform 1 0 89378 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1936
timestamp 1712078602
transform 1 0 89608 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1948
timestamp 1712078602
transform 1 0 90160 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1960
timestamp 1712078602
transform 1 0 90712 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1972
timestamp 1712078602
transform 1 0 91264 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_1984
timestamp 1712078602
transform 1 0 91816 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_1989
timestamp 1712078602
transform 1 0 92046 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2001
timestamp 1712078602
transform 1 0 92598 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2013
timestamp 1712078602
transform 1 0 93150 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2025
timestamp 1712078602
transform 1 0 93702 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2037
timestamp 1712078602
transform 1 0 94254 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2043
timestamp 1712078602
transform 1 0 94530 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_16_2045
timestamp 1712078602
transform 1 0 94622 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2053
timestamp 1712078602
transform 1 0 94990 0 1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2058
timestamp 1712078602
transform 1 0 95220 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_16_2065
timestamp 1712078602
transform 1 0 95542 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2073
timestamp 1712078602
transform 1 0 95910 0 1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2095
timestamp 1712078602
transform 1 0 96922 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2099
timestamp 1712078602
transform 1 0 97106 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2110
timestamp 1712078602
transform 1 0 97612 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2117
timestamp 1712078602
transform 1 0 97934 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2129
timestamp 1712078602
transform 1 0 98486 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2141
timestamp 1712078602
transform 1 0 99038 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_16_2153
timestamp 1712078602
transform 1 0 99590 0 1 5440
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2157
timestamp 1712078602
transform 1 0 99774 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2169
timestamp 1712078602
transform 1 0 100326 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2181
timestamp 1712078602
transform 1 0 100878 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2188
timestamp 1712078602
transform 1 0 101200 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2195
timestamp 1712078602
transform 1 0 101522 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_16_2202
timestamp 1712078602
transform 1 0 101844 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2210
timestamp 1712078602
transform 1 0 102212 0 1 5440
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2216
timestamp 1712078602
transform 1 0 102488 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2228
timestamp 1712078602
transform 1 0 103040 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2240
timestamp 1712078602
transform 1 0 103592 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2252
timestamp 1712078602
transform 1 0 104144 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2264
timestamp 1712078602
transform 1 0 104696 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2269
timestamp 1712078602
transform 1 0 104926 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2281
timestamp 1712078602
transform 1 0 105478 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2293
timestamp 1712078602
transform 1 0 106030 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2305
timestamp 1712078602
transform 1 0 106582 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2317
timestamp 1712078602
transform 1 0 107134 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2323
timestamp 1712078602
transform 1 0 107410 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2325
timestamp 1712078602
transform 1 0 107502 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2337
timestamp 1712078602
transform 1 0 108054 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2349
timestamp 1712078602
transform 1 0 108606 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2361
timestamp 1712078602
transform 1 0 109158 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2373
timestamp 1712078602
transform 1 0 109710 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2379
timestamp 1712078602
transform 1 0 109986 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2381
timestamp 1712078602
transform 1 0 110078 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2393
timestamp 1712078602
transform 1 0 110630 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2405
timestamp 1712078602
transform 1 0 111182 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2417
timestamp 1712078602
transform 1 0 111734 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2429
timestamp 1712078602
transform 1 0 112286 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2435
timestamp 1712078602
transform 1 0 112562 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2437
timestamp 1712078602
transform 1 0 112654 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2449
timestamp 1712078602
transform 1 0 113206 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2461
timestamp 1712078602
transform 1 0 113758 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2473
timestamp 1712078602
transform 1 0 114310 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__decap_8  FILLER_16_2482
timestamp 1712078602
transform 1 0 114724 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2490
timestamp 1712078602
transform 1 0 115092 0 1 5440
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2493
timestamp 1712078602
transform 1 0 115230 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2505
timestamp 1712078602
transform 1 0 115782 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2517
timestamp 1712078602
transform 1 0 116334 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2529
timestamp 1712078602
transform 1 0 116886 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2541
timestamp 1712078602
transform 1 0 117438 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2547
timestamp 1712078602
transform 1 0 117714 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2549
timestamp 1712078602
transform 1 0 117806 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2561
timestamp 1712078602
transform 1 0 118358 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2573
timestamp 1712078602
transform 1 0 118910 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_16_2585
timestamp 1712078602
transform 1 0 119462 0 1 5440
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2593
timestamp 1712078602
transform 1 0 119830 0 1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2598
timestamp 1712078602
transform 1 0 120060 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2608
timestamp 1712078602
transform 1 0 120520 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2615
timestamp 1712078602
transform 1 0 120842 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2622
timestamp 1712078602
transform 1 0 121164 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2634
timestamp 1712078602
transform 1 0 121716 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2646
timestamp 1712078602
transform 1 0 122268 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2658
timestamp 1712078602
transform 1 0 122820 0 1 5440
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2661
timestamp 1712078602
transform 1 0 122958 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2673
timestamp 1712078602
transform 1 0 123510 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2685
timestamp 1712078602
transform 1 0 124062 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2697
timestamp 1712078602
transform 1 0 124614 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2709
timestamp 1712078602
transform 1 0 125166 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2715
timestamp 1712078602
transform 1 0 125442 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2717
timestamp 1712078602
transform 1 0 125534 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_16_2729
timestamp 1712078602
transform 1 0 126086 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2735
timestamp 1712078602
transform 1 0 126362 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2742
timestamp 1712078602
transform 1 0 126684 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2749
timestamp 1712078602
transform 1 0 127006 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2756
timestamp 1712078602
transform 1 0 127328 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2768
timestamp 1712078602
transform 1 0 127880 0 1 5440
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2773
timestamp 1712078602
transform 1 0 128110 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2785
timestamp 1712078602
transform 1 0 128662 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2797
timestamp 1712078602
transform 1 0 129214 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2809
timestamp 1712078602
transform 1 0 129766 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2821
timestamp 1712078602
transform 1 0 130318 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2827
timestamp 1712078602
transform 1 0 130594 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2829
timestamp 1712078602
transform 1 0 130686 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2841
timestamp 1712078602
transform 1 0 131238 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2853
timestamp 1712078602
transform 1 0 131790 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2865
timestamp 1712078602
transform 1 0 132342 0 1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2870
timestamp 1712078602
transform 1 0 132572 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2877
timestamp 1712078602
transform 1 0 132894 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2883
timestamp 1712078602
transform 1 0 133170 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_16_2885
timestamp 1712078602
transform 1 0 133262 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2897
timestamp 1712078602
transform 1 0 133814 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2904
timestamp 1712078602
transform 1 0 134136 0 1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_16_2908
timestamp 1712078602
transform 1 0 134320 0 1 5440
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_16_2919
timestamp 1712078602
transform 1 0 134826 0 1 5440
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_16_2932
timestamp 1712078602
transform 1 0 135424 0 1 5440
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2941
timestamp 1712078602
transform 1 0 135838 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2953
timestamp 1712078602
transform 1 0 136390 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2965
timestamp 1712078602
transform 1 0 136942 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2977
timestamp 1712078602
transform 1 0 137494 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_2989
timestamp 1712078602
transform 1 0 138046 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_2995
timestamp 1712078602
transform 1 0 138322 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_2997
timestamp 1712078602
transform 1 0 138414 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3009
timestamp 1712078602
transform 1 0 138966 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3021
timestamp 1712078602
transform 1 0 139518 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3033
timestamp 1712078602
transform 1 0 140070 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_3045
timestamp 1712078602
transform 1 0 140622 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_3051
timestamp 1712078602
transform 1 0 140898 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3053
timestamp 1712078602
transform 1 0 140990 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3065
timestamp 1712078602
transform 1 0 141542 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3077
timestamp 1712078602
transform 1 0 142094 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3089
timestamp 1712078602
transform 1 0 142646 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_3101
timestamp 1712078602
transform 1 0 143198 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_3107
timestamp 1712078602
transform 1 0 143474 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3109
timestamp 1712078602
transform 1 0 143566 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3121
timestamp 1712078602
transform 1 0 144118 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3133
timestamp 1712078602
transform 1 0 144670 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3145
timestamp 1712078602
transform 1 0 145222 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_3157
timestamp 1712078602
transform 1 0 145774 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_3163
timestamp 1712078602
transform 1 0 146050 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3165
timestamp 1712078602
transform 1 0 146142 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3177
timestamp 1712078602
transform 1 0 146694 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3189
timestamp 1712078602
transform 1 0 147246 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3201
timestamp 1712078602
transform 1 0 147798 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_3213
timestamp 1712078602
transform 1 0 148350 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_3219
timestamp 1712078602
transform 1 0 148626 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3221
timestamp 1712078602
transform 1 0 148718 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3233
timestamp 1712078602
transform 1 0 149270 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3245
timestamp 1712078602
transform 1 0 149822 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3257
timestamp 1712078602
transform 1 0 150374 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_16_3269
timestamp 1712078602
transform 1 0 150926 0 1 5440
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_16_3275
timestamp 1712078602
transform 1 0 151202 0 1 5440
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3277
timestamp 1712078602
transform 1 0 151294 0 1 5440
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_16_3289
timestamp 1712078602
transform 1 0 151846 0 1 5440
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_16_3301
timestamp 1712078602
transform 1 0 152398 0 1 5440
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1712078602
transform 1 0 690 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1712078602
transform 1 0 1242 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1712078602
transform 1 0 1794 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1712078602
transform 1 0 2346 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1712078602
transform 1 0 2898 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1712078602
transform 1 0 3082 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1712078602
transform 1 0 3174 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1712078602
transform 1 0 3726 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1712078602
transform 1 0 4278 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1712078602
transform 1 0 4830 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1712078602
transform 1 0 5382 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1712078602
transform 1 0 5658 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1712078602
transform 1 0 5750 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1712078602
transform 1 0 6302 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1712078602
transform 1 0 6854 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1712078602
transform 1 0 7406 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1712078602
transform 1 0 7958 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1712078602
transform 1 0 8234 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1712078602
transform 1 0 8326 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1712078602
transform 1 0 8878 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1712078602
transform 1 0 9430 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1712078602
transform 1 0 9982 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1712078602
transform 1 0 10534 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1712078602
transform 1 0 10810 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1712078602
transform 1 0 10902 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1712078602
transform 1 0 11454 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1712078602
transform 1 0 12006 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1712078602
transform 1 0 12558 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1712078602
transform 1 0 13110 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1712078602
transform 1 0 13386 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_17_281
timestamp 1712078602
transform 1 0 13478 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_17_289
timestamp 1712078602
transform 1 0 13846 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1712078602
transform 1 0 14030 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1712078602
transform 1 0 14628 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_17_330
timestamp 1712078602
transform 1 0 15732 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_8  FILLER_17_346
timestamp 1712078602
transform 1 0 16468 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1712078602
transform 1 0 16974 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_364
timestamp 1712078602
transform 1 0 17296 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_371
timestamp 1712078602
transform 1 0 17618 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_17_383
timestamp 1712078602
transform 1 0 18170 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1712078602
transform 1 0 18538 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1712078602
transform 1 0 18630 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_408
timestamp 1712078602
transform 1 0 19320 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_415
timestamp 1712078602
transform 1 0 19642 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_17_428
timestamp 1712078602
transform 1 0 20240 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_17_437
timestamp 1712078602
transform 1 0 20654 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_444
timestamp 1712078602
transform 1 0 20976 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_449
timestamp 1712078602
transform 1 0 21206 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_17_457
timestamp 1712078602
transform 1 0 21574 0 -1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1712078602
transform 1 0 21758 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1712078602
transform 1 0 22310 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1712078602
transform 1 0 22862 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1712078602
transform 1 0 23414 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1712078602
transform 1 0 23690 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1712078602
transform 1 0 23782 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1712078602
transform 1 0 24334 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1712078602
transform 1 0 24886 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1712078602
transform 1 0 25438 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1712078602
transform 1 0 25990 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1712078602
transform 1 0 26266 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_17_561
timestamp 1712078602
transform 1 0 26358 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_17_565
timestamp 1712078602
transform 1 0 26542 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_17_574
timestamp 1712078602
transform 1 0 26956 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_581
timestamp 1712078602
transform 1 0 27278 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_17_594
timestamp 1712078602
transform 1 0 27876 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_600
timestamp 1712078602
transform 1 0 28152 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_604
timestamp 1712078602
transform 1 0 28336 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_611
timestamp 1712078602
transform 1 0 28658 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1712078602
transform 1 0 28842 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1712078602
transform 1 0 28934 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1712078602
transform 1 0 29486 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1712078602
transform 1 0 30038 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1712078602
transform 1 0 30590 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1712078602
transform 1 0 31142 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1712078602
transform 1 0 31418 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1712078602
transform 1 0 31510 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1712078602
transform 1 0 32062 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1712078602
transform 1 0 32614 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1712078602
transform 1 0 33166 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1712078602
transform 1 0 33718 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1712078602
transform 1 0 33994 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1712078602
transform 1 0 34086 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1712078602
transform 1 0 34638 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1712078602
transform 1 0 35190 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1712078602
transform 1 0 35742 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1712078602
transform 1 0 36294 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1712078602
transform 1 0 36570 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1712078602
transform 1 0 36662 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1712078602
transform 1 0 37214 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_818
timestamp 1712078602
transform 1 0 38180 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_6  FILLER_17_827
timestamp 1712078602
transform 1 0 38594 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_17_836
timestamp 1712078602
transform 1 0 39008 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_844
timestamp 1712078602
transform 1 0 39376 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_856
timestamp 1712078602
transform 1 0 39928 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_868
timestamp 1712078602
transform 1 0 40480 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_880
timestamp 1712078602
transform 1 0 41032 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_892
timestamp 1712078602
transform 1 0 41584 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_17_897
timestamp 1712078602
transform 1 0 41814 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_17_908
timestamp 1712078602
transform 1 0 42320 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_915
timestamp 1712078602
transform 1 0 42642 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_928
timestamp 1712078602
transform 1 0 43240 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_932
timestamp 1712078602
transform 1 0 43424 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_937
timestamp 1712078602
transform 1 0 43654 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1712078602
transform 1 0 44022 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1712078602
transform 1 0 44298 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_956
timestamp 1712078602
transform 1 0 44528 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_968
timestamp 1712078602
transform 1 0 45080 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_980
timestamp 1712078602
transform 1 0 45632 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_992
timestamp 1712078602
transform 1 0 46184 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1004
timestamp 1712078602
transform 1 0 46736 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1009
timestamp 1712078602
transform 1 0 46966 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1021
timestamp 1712078602
transform 1 0 47518 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1033
timestamp 1712078602
transform 1 0 48070 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1045
timestamp 1712078602
transform 1 0 48622 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1057
timestamp 1712078602
transform 1 0 49174 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1712078602
transform 1 0 49450 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1065
timestamp 1712078602
transform 1 0 49542 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1080
timestamp 1712078602
transform 1 0 50232 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1087
timestamp 1712078602
transform 1 0 50554 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1100
timestamp 1712078602
transform 1 0 51152 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1106
timestamp 1712078602
transform 1 0 51428 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_17_1110
timestamp 1712078602
transform 1 0 51612 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_17_1118
timestamp 1712078602
transform 1 0 51980 0 -1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1121
timestamp 1712078602
transform 1 0 52118 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1133
timestamp 1712078602
transform 1 0 52670 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1145
timestamp 1712078602
transform 1 0 53222 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1157
timestamp 1712078602
transform 1 0 53774 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1169
timestamp 1712078602
transform 1 0 54326 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1175
timestamp 1712078602
transform 1 0 54602 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1177
timestamp 1712078602
transform 1 0 54694 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1189
timestamp 1712078602
transform 1 0 55246 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1201
timestamp 1712078602
transform 1 0 55798 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1213
timestamp 1712078602
transform 1 0 56350 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1228
timestamp 1712078602
transform 1 0 57040 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1233
timestamp 1712078602
transform 1 0 57270 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_17_1243
timestamp 1712078602
transform 1 0 57730 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1254
timestamp 1712078602
transform 1 0 58236 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1261
timestamp 1712078602
transform 1 0 58558 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1268
timestamp 1712078602
transform 1 0 58880 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_17_1280
timestamp 1712078602
transform 1 0 59432 0 -1 5984
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1289
timestamp 1712078602
transform 1 0 59846 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1301
timestamp 1712078602
transform 1 0 60398 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1313
timestamp 1712078602
transform 1 0 60950 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1325
timestamp 1712078602
transform 1 0 61502 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1337
timestamp 1712078602
transform 1 0 62054 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1343
timestamp 1712078602
transform 1 0 62330 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1345
timestamp 1712078602
transform 1 0 62422 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1357
timestamp 1712078602
transform 1 0 62974 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1369
timestamp 1712078602
transform 1 0 63526 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1381
timestamp 1712078602
transform 1 0 64078 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1396
timestamp 1712078602
transform 1 0 64768 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1401
timestamp 1712078602
transform 1 0 64998 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1405
timestamp 1712078602
transform 1 0 65182 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1415
timestamp 1712078602
transform 1 0 65642 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1423
timestamp 1712078602
transform 1 0 66010 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1430
timestamp 1712078602
transform 1 0 66332 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1442
timestamp 1712078602
transform 1 0 66884 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_17_1454
timestamp 1712078602
transform 1 0 67436 0 -1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1457
timestamp 1712078602
transform 1 0 67574 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1469
timestamp 1712078602
transform 1 0 68126 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1481
timestamp 1712078602
transform 1 0 68678 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1493
timestamp 1712078602
transform 1 0 69230 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1505
timestamp 1712078602
transform 1 0 69782 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1511
timestamp 1712078602
transform 1 0 70058 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1513
timestamp 1712078602
transform 1 0 70150 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1525
timestamp 1712078602
transform 1 0 70702 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1537
timestamp 1712078602
transform 1 0 71254 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1549
timestamp 1712078602
transform 1 0 71806 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1561
timestamp 1712078602
transform 1 0 72358 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1567
timestamp 1712078602
transform 1 0 72634 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1569
timestamp 1712078602
transform 1 0 72726 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_17_1581
timestamp 1712078602
transform 1 0 73278 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_17_1589
timestamp 1712078602
transform 1 0 73646 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1595
timestamp 1712078602
transform 1 0 73922 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1599
timestamp 1712078602
transform 1 0 74106 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1620
timestamp 1712078602
transform 1 0 75072 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1625
timestamp 1712078602
transform 1 0 75302 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1629
timestamp 1712078602
transform 1 0 75486 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1633
timestamp 1712078602
transform 1 0 75670 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1639
timestamp 1712078602
transform 1 0 75946 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1643
timestamp 1712078602
transform 1 0 76130 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1650
timestamp 1712078602
transform 1 0 76452 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1662
timestamp 1712078602
transform 1 0 77004 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1674
timestamp 1712078602
transform 1 0 77556 0 -1 5984
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1681
timestamp 1712078602
transform 1 0 77878 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1693
timestamp 1712078602
transform 1 0 78430 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1705
timestamp 1712078602
transform 1 0 78982 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1717
timestamp 1712078602
transform 1 0 79534 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1729
timestamp 1712078602
transform 1 0 80086 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1735
timestamp 1712078602
transform 1 0 80362 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1740
timestamp 1712078602
transform 1 0 80592 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1747
timestamp 1712078602
transform 1 0 80914 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1754
timestamp 1712078602
transform 1 0 81236 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1761
timestamp 1712078602
transform 1 0 81558 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1768
timestamp 1712078602
transform 1 0 81880 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1775
timestamp 1712078602
transform 1 0 82202 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_17_1782
timestamp 1712078602
transform 1 0 82524 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_17_1790
timestamp 1712078602
transform 1 0 82892 0 -1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1793
timestamp 1712078602
transform 1 0 83030 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1805
timestamp 1712078602
transform 1 0 83582 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1817
timestamp 1712078602
transform 1 0 84134 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1829
timestamp 1712078602
transform 1 0 84686 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1841
timestamp 1712078602
transform 1 0 85238 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1847
timestamp 1712078602
transform 1 0 85514 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1849
timestamp 1712078602
transform 1 0 85606 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1861
timestamp 1712078602
transform 1 0 86158 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1873
timestamp 1712078602
transform 1 0 86710 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1885
timestamp 1712078602
transform 1 0 87262 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_1897
timestamp 1712078602
transform 1 0 87814 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1903
timestamp 1712078602
transform 1 0 88090 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1905
timestamp 1712078602
transform 1 0 88182 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_17_1909
timestamp 1712078602
transform 1 0 88366 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1917
timestamp 1712078602
transform 1 0 88734 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1927
timestamp 1712078602
transform 1 0 89194 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_1940
timestamp 1712078602
transform 1 0 89792 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1947
timestamp 1712078602
transform 1 0 90114 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_17_1959
timestamp 1712078602
transform 1 0 90666 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1961
timestamp 1712078602
transform 1 0 90758 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1973
timestamp 1712078602
transform 1 0 91310 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1985
timestamp 1712078602
transform 1 0 91862 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_1997
timestamp 1712078602
transform 1 0 92414 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2009
timestamp 1712078602
transform 1 0 92966 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2015
timestamp 1712078602
transform 1 0 93242 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2017
timestamp 1712078602
transform 1 0 93334 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2029
timestamp 1712078602
transform 1 0 93886 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2041
timestamp 1712078602
transform 1 0 94438 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2050
timestamp 1712078602
transform 1 0 94852 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2057
timestamp 1712078602
transform 1 0 95174 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_17_2064
timestamp 1712078602
transform 1 0 95496 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2093
timestamp 1712078602
transform 1 0 96830 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2117
timestamp 1712078602
transform 1 0 97934 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2124
timestamp 1712078602
transform 1 0 98256 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2129
timestamp 1712078602
transform 1 0 98486 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2141
timestamp 1712078602
transform 1 0 99038 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2153
timestamp 1712078602
transform 1 0 99590 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2165
timestamp 1712078602
transform 1 0 100142 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2177
timestamp 1712078602
transform 1 0 100694 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2183
timestamp 1712078602
transform 1 0 100970 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2185
timestamp 1712078602
transform 1 0 101062 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2189
timestamp 1712078602
transform 1 0 101246 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2196
timestamp 1712078602
transform 1 0 101568 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2200
timestamp 1712078602
transform 1 0 101752 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2210
timestamp 1712078602
transform 1 0 102212 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2223
timestamp 1712078602
transform 1 0 102810 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2235
timestamp 1712078602
transform 1 0 103362 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2239
timestamp 1712078602
transform 1 0 103546 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2241
timestamp 1712078602
transform 1 0 103638 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2253
timestamp 1712078602
transform 1 0 104190 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2265
timestamp 1712078602
transform 1 0 104742 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2277
timestamp 1712078602
transform 1 0 105294 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2289
timestamp 1712078602
transform 1 0 105846 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2295
timestamp 1712078602
transform 1 0 106122 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2297
timestamp 1712078602
transform 1 0 106214 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2309
timestamp 1712078602
transform 1 0 106766 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2321
timestamp 1712078602
transform 1 0 107318 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2333
timestamp 1712078602
transform 1 0 107870 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2345
timestamp 1712078602
transform 1 0 108422 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2351
timestamp 1712078602
transform 1 0 108698 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2353
timestamp 1712078602
transform 1 0 108790 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2365
timestamp 1712078602
transform 1 0 109342 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2377
timestamp 1712078602
transform 1 0 109894 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2389
timestamp 1712078602
transform 1 0 110446 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2401
timestamp 1712078602
transform 1 0 110998 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2407
timestamp 1712078602
transform 1 0 111274 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2409
timestamp 1712078602
transform 1 0 111366 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2421
timestamp 1712078602
transform 1 0 111918 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2433
timestamp 1712078602
transform 1 0 112470 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2445
timestamp 1712078602
transform 1 0 113022 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2457
timestamp 1712078602
transform 1 0 113574 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2463
timestamp 1712078602
transform 1 0 113850 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2474
timestamp 1712078602
transform 1 0 114356 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2487
timestamp 1712078602
transform 1 0 114954 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2494
timestamp 1712078602
transform 1 0 115276 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2501
timestamp 1712078602
transform 1 0 115598 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2508
timestamp 1712078602
transform 1 0 115920 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2521
timestamp 1712078602
transform 1 0 116518 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2533
timestamp 1712078602
transform 1 0 117070 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2545
timestamp 1712078602
transform 1 0 117622 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2557
timestamp 1712078602
transform 1 0 118174 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2569
timestamp 1712078602
transform 1 0 118726 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2575
timestamp 1712078602
transform 1 0 119002 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2577
timestamp 1712078602
transform 1 0 119094 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_17_2585
timestamp 1712078602
transform 1 0 119462 0 -1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_17_2593
timestamp 1712078602
transform 1 0 119830 0 -1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2604
timestamp 1712078602
transform 1 0 120336 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2611
timestamp 1712078602
transform 1 0 120658 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2618
timestamp 1712078602
transform 1 0 120980 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2625
timestamp 1712078602
transform 1 0 121302 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2631
timestamp 1712078602
transform 1 0 121578 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2633
timestamp 1712078602
transform 1 0 121670 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2645
timestamp 1712078602
transform 1 0 122222 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2657
timestamp 1712078602
transform 1 0 122774 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2669
timestamp 1712078602
transform 1 0 123326 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2681
timestamp 1712078602
transform 1 0 123878 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2687
timestamp 1712078602
transform 1 0 124154 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2689
timestamp 1712078602
transform 1 0 124246 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2701
timestamp 1712078602
transform 1 0 124798 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2713
timestamp 1712078602
transform 1 0 125350 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_17_2728
timestamp 1712078602
transform 1 0 126040 0 -1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_17_2732
timestamp 1712078602
transform 1 0 126224 0 -1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2738
timestamp 1712078602
transform 1 0 126500 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2754
timestamp 1712078602
transform 1 0 127236 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2761
timestamp 1712078602
transform 1 0 127558 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2768
timestamp 1712078602
transform 1 0 127880 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2780
timestamp 1712078602
transform 1 0 128432 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_17_2792
timestamp 1712078602
transform 1 0 128984 0 -1 5984
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2801
timestamp 1712078602
transform 1 0 129398 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2813
timestamp 1712078602
transform 1 0 129950 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2825
timestamp 1712078602
transform 1 0 130502 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2837
timestamp 1712078602
transform 1 0 131054 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_2849
timestamp 1712078602
transform 1 0 131606 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_2855
timestamp 1712078602
transform 1 0 131882 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2857
timestamp 1712078602
transform 1 0 131974 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2864
timestamp 1712078602
transform 1 0 132296 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2871
timestamp 1712078602
transform 1 0 132618 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2895
timestamp 1712078602
transform 1 0 133722 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2908
timestamp 1712078602
transform 1 0 134320 0 -1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2933
timestamp 1712078602
transform 1 0 135470 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2940
timestamp 1712078602
transform 1 0 135792 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2952
timestamp 1712078602
transform 1 0 136344 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_17_2964
timestamp 1712078602
transform 1 0 136896 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2969
timestamp 1712078602
transform 1 0 137126 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2981
timestamp 1712078602
transform 1 0 137678 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_2993
timestamp 1712078602
transform 1 0 138230 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3005
timestamp 1712078602
transform 1 0 138782 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_3017
timestamp 1712078602
transform 1 0 139334 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_3023
timestamp 1712078602
transform 1 0 139610 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3025
timestamp 1712078602
transform 1 0 139702 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3037
timestamp 1712078602
transform 1 0 140254 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3049
timestamp 1712078602
transform 1 0 140806 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3061
timestamp 1712078602
transform 1 0 141358 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_3073
timestamp 1712078602
transform 1 0 141910 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_3079
timestamp 1712078602
transform 1 0 142186 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3081
timestamp 1712078602
transform 1 0 142278 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3093
timestamp 1712078602
transform 1 0 142830 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3105
timestamp 1712078602
transform 1 0 143382 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3117
timestamp 1712078602
transform 1 0 143934 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_3129
timestamp 1712078602
transform 1 0 144486 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_3135
timestamp 1712078602
transform 1 0 144762 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3137
timestamp 1712078602
transform 1 0 144854 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3149
timestamp 1712078602
transform 1 0 145406 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3161
timestamp 1712078602
transform 1 0 145958 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3173
timestamp 1712078602
transform 1 0 146510 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_3185
timestamp 1712078602
transform 1 0 147062 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_3191
timestamp 1712078602
transform 1 0 147338 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3193
timestamp 1712078602
transform 1 0 147430 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3205
timestamp 1712078602
transform 1 0 147982 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3217
timestamp 1712078602
transform 1 0 148534 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3229
timestamp 1712078602
transform 1 0 149086 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_3241
timestamp 1712078602
transform 1 0 149638 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_3247
timestamp 1712078602
transform 1 0 149914 0 -1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3249
timestamp 1712078602
transform 1 0 150006 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3261
timestamp 1712078602
transform 1 0 150558 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3273
timestamp 1712078602
transform 1 0 151110 0 -1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_17_3285
timestamp 1712078602
transform 1 0 151662 0 -1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_17_3297
timestamp 1712078602
transform 1 0 152214 0 -1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_17_3303
timestamp 1712078602
transform 1 0 152490 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_17_3305
timestamp 1712078602
transform 1 0 152582 0 -1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1712078602
transform 1 0 690 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1712078602
transform 1 0 1242 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1712078602
transform 1 0 1794 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1712078602
transform 1 0 1886 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1712078602
transform 1 0 2438 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1712078602
transform 1 0 2990 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1712078602
transform 1 0 3542 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1712078602
transform 1 0 4094 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1712078602
transform 1 0 4370 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1712078602
transform 1 0 4462 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1712078602
transform 1 0 5014 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1712078602
transform 1 0 5566 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1712078602
transform 1 0 6118 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1712078602
transform 1 0 6670 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1712078602
transform 1 0 6946 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1712078602
transform 1 0 7038 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1712078602
transform 1 0 7590 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1712078602
transform 1 0 8142 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1712078602
transform 1 0 8694 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1712078602
transform 1 0 9246 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1712078602
transform 1 0 9522 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1712078602
transform 1 0 9614 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1712078602
transform 1 0 10166 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1712078602
transform 1 0 10718 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1712078602
transform 1 0 11270 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1712078602
transform 1 0 11822 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1712078602
transform 1 0 12098 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1712078602
transform 1 0 12190 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1712078602
transform 1 0 12742 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_277
timestamp 1712078602
transform 1 0 13294 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_281
timestamp 1712078602
transform 1 0 13478 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1712078602
transform 1 0 13938 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1712078602
transform 1 0 14536 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_329
timestamp 1712078602
transform 1 0 15686 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_353
timestamp 1712078602
transform 1 0 16790 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1712078602
transform 1 0 17112 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_368
timestamp 1712078602
transform 1 0 17480 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_18_375
timestamp 1712078602
transform 1 0 17802 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_381
timestamp 1712078602
transform 1 0 18078 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1712078602
transform 1 0 18308 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_394
timestamp 1712078602
transform 1 0 18676 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_409
timestamp 1712078602
transform 1 0 19366 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1712078602
transform 1 0 19688 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1712078602
transform 1 0 19918 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1712078602
transform 1 0 20516 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_458
timestamp 1712078602
transform 1 0 21620 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_18_466
timestamp 1712078602
transform 1 0 21988 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1712078602
transform 1 0 22356 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1712078602
transform 1 0 22494 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1712078602
transform 1 0 23046 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1712078602
transform 1 0 23598 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1712078602
transform 1 0 24150 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1712078602
transform 1 0 24702 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1712078602
transform 1 0 24978 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1712078602
transform 1 0 25070 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1712078602
transform 1 0 25622 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_577
timestamp 1712078602
transform 1 0 27094 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_584
timestamp 1712078602
transform 1 0 27416 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_589
timestamp 1712078602
transform 1 0 27646 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_18_594
timestamp 1712078602
transform 1 0 27876 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_18_607
timestamp 1712078602
transform 1 0 28474 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_614
timestamp 1712078602
transform 1 0 28796 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_621
timestamp 1712078602
transform 1 0 29118 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_633
timestamp 1712078602
transform 1 0 29670 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_18_641
timestamp 1712078602
transform 1 0 30038 0 1 5984
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1712078602
transform 1 0 30222 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1712078602
transform 1 0 30774 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1712078602
transform 1 0 31326 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1712078602
transform 1 0 31878 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1712078602
transform 1 0 32430 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1712078602
transform 1 0 32706 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1712078602
transform 1 0 32798 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1712078602
transform 1 0 33350 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1712078602
transform 1 0 33902 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1712078602
transform 1 0 34454 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1712078602
transform 1 0 35006 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1712078602
transform 1 0 35282 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1712078602
transform 1 0 35374 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1712078602
transform 1 0 35926 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1712078602
transform 1 0 36478 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1712078602
transform 1 0 37030 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_808
timestamp 1712078602
transform 1 0 37720 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_813
timestamp 1712078602
transform 1 0 37950 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_826
timestamp 1712078602
transform 1 0 38548 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_18_839
timestamp 1712078602
transform 1 0 39146 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_18_847
timestamp 1712078602
transform 1 0 39514 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_18_852
timestamp 1712078602
transform 1 0 39744 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_858
timestamp 1712078602
transform 1 0 40020 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_18_862
timestamp 1712078602
transform 1 0 40204 0 1 5984
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_18_869
timestamp 1712078602
transform 1 0 40526 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_881
timestamp 1712078602
transform 1 0 41078 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_893
timestamp 1712078602
transform 1 0 41630 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_6  FILLER_18_910
timestamp 1712078602
transform 1 0 42412 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_916
timestamp 1712078602
transform 1 0 42688 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_920
timestamp 1712078602
transform 1 0 42872 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_18_925
timestamp 1712078602
transform 1 0 43102 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_18_936
timestamp 1712078602
transform 1 0 43608 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_949
timestamp 1712078602
transform 1 0 44206 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_956
timestamp 1712078602
transform 1 0 44528 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_963
timestamp 1712078602
transform 1 0 44850 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_18_970
timestamp 1712078602
transform 1 0 45172 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_18_978
timestamp 1712078602
transform 1 0 45540 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_981
timestamp 1712078602
transform 1 0 45678 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_993
timestamp 1712078602
transform 1 0 46230 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1005
timestamp 1712078602
transform 1 0 46782 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1017
timestamp 1712078602
transform 1 0 47334 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1029
timestamp 1712078602
transform 1 0 47886 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1035
timestamp 1712078602
transform 1 0 48162 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1037
timestamp 1712078602
transform 1 0 48254 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1049
timestamp 1712078602
transform 1 0 48806 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1061
timestamp 1712078602
transform 1 0 49358 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1068
timestamp 1712078602
transform 1 0 49680 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1075
timestamp 1712078602
transform 1 0 50002 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1088
timestamp 1712078602
transform 1 0 50600 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_18_1093
timestamp 1712078602
transform 1 0 50830 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1099
timestamp 1712078602
transform 1 0 51106 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1112
timestamp 1712078602
transform 1 0 51704 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1119
timestamp 1712078602
transform 1 0 52026 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1126
timestamp 1712078602
transform 1 0 52348 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1133
timestamp 1712078602
transform 1 0 52670 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_18_1145
timestamp 1712078602
transform 1 0 53222 0 1 5984
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1149
timestamp 1712078602
transform 1 0 53406 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1161
timestamp 1712078602
transform 1 0 53958 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1173
timestamp 1712078602
transform 1 0 54510 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1185
timestamp 1712078602
transform 1 0 55062 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1197
timestamp 1712078602
transform 1 0 55614 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1203
timestamp 1712078602
transform 1 0 55890 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1205
timestamp 1712078602
transform 1 0 55982 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1220
timestamp 1712078602
transform 1 0 56672 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1227
timestamp 1712078602
transform 1 0 56994 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_18_1251
timestamp 1712078602
transform 1 0 58098 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1712078602
transform 1 0 58466 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1270
timestamp 1712078602
transform 1 0 58972 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1277
timestamp 1712078602
transform 1 0 59294 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1289
timestamp 1712078602
transform 1 0 59846 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1301
timestamp 1712078602
transform 1 0 60398 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_18_1313
timestamp 1712078602
transform 1 0 60950 0 1 5984
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1317
timestamp 1712078602
transform 1 0 61134 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1329
timestamp 1712078602
transform 1 0 61686 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1341
timestamp 1712078602
transform 1 0 62238 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1353
timestamp 1712078602
transform 1 0 62790 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1365
timestamp 1712078602
transform 1 0 63342 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1371
timestamp 1712078602
transform 1 0 63618 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_18_1373
timestamp 1712078602
transform 1 0 63710 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1379
timestamp 1712078602
transform 1 0 63986 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1383
timestamp 1712078602
transform 1 0 64170 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1387
timestamp 1712078602
transform 1 0 64354 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1411
timestamp 1712078602
transform 1 0 65458 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1424
timestamp 1712078602
transform 1 0 66056 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1432
timestamp 1712078602
transform 1 0 66424 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1444
timestamp 1712078602
transform 1 0 66976 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1456
timestamp 1712078602
transform 1 0 67528 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1468
timestamp 1712078602
transform 1 0 68080 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1480
timestamp 1712078602
transform 1 0 68632 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1491
timestamp 1712078602
transform 1 0 69138 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1503
timestamp 1712078602
transform 1 0 69690 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1515
timestamp 1712078602
transform 1 0 70242 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1527
timestamp 1712078602
transform 1 0 70794 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1539
timestamp 1712078602
transform 1 0 71346 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1541
timestamp 1712078602
transform 1 0 71438 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1553
timestamp 1712078602
transform 1 0 71990 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1565
timestamp 1712078602
transform 1 0 72542 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1571
timestamp 1712078602
transform 1 0 72818 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_18_1578
timestamp 1712078602
transform 1 0 73140 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_18_1586
timestamp 1712078602
transform 1 0 73508 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1592
timestamp 1712078602
transform 1 0 73784 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_18_1597
timestamp 1712078602
transform 1 0 74014 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_8  FILLER_18_1603
timestamp 1712078602
transform 1 0 74290 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1611
timestamp 1712078602
transform 1 0 74658 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1632
timestamp 1712078602
transform 1 0 75624 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1648
timestamp 1712078602
transform 1 0 76360 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1653
timestamp 1712078602
transform 1 0 76590 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1666
timestamp 1712078602
transform 1 0 77188 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1678
timestamp 1712078602
transform 1 0 77740 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1690
timestamp 1712078602
transform 1 0 78292 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1702
timestamp 1712078602
transform 1 0 78844 0 1 5984
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1709
timestamp 1712078602
transform 1 0 79166 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1721
timestamp 1712078602
transform 1 0 79718 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1730
timestamp 1712078602
transform 1 0 80132 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1745
timestamp 1712078602
transform 1 0 80822 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1758
timestamp 1712078602
transform 1 0 81420 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1765
timestamp 1712078602
transform 1 0 81742 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1786
timestamp 1712078602
transform 1 0 82708 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1794
timestamp 1712078602
transform 1 0 83076 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1806
timestamp 1712078602
transform 1 0 83628 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_18_1818
timestamp 1712078602
transform 1 0 84180 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1821
timestamp 1712078602
transform 1 0 84318 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1833
timestamp 1712078602
transform 1 0 84870 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1845
timestamp 1712078602
transform 1 0 85422 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1857
timestamp 1712078602
transform 1 0 85974 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1869
timestamp 1712078602
transform 1 0 86526 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1875
timestamp 1712078602
transform 1 0 86802 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1877
timestamp 1712078602
transform 1 0 86894 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_1889
timestamp 1712078602
transform 1 0 87446 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_18_1897
timestamp 1712078602
transform 1 0 87814 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1903
timestamp 1712078602
transform 1 0 88090 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1916
timestamp 1712078602
transform 1 0 88688 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1920
timestamp 1712078602
transform 1 0 88872 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_18_1925
timestamp 1712078602
transform 1 0 89102 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_1931
timestamp 1712078602
transform 1 0 89378 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_18_1933
timestamp 1712078602
transform 1 0 89470 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_18_1955
timestamp 1712078602
transform 1 0 90482 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1962
timestamp 1712078602
transform 1 0 90804 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1974
timestamp 1712078602
transform 1 0 91356 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_18_1986
timestamp 1712078602
transform 1 0 91908 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_1989
timestamp 1712078602
transform 1 0 92046 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2001
timestamp 1712078602
transform 1 0 92598 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2013
timestamp 1712078602
transform 1 0 93150 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2025
timestamp 1712078602
transform 1 0 93702 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2040
timestamp 1712078602
transform 1 0 94392 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_18_2045
timestamp 1712078602
transform 1 0 94622 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2051
timestamp 1712078602
transform 1 0 94898 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2058
timestamp 1712078602
transform 1 0 95220 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2082
timestamp 1712078602
transform 1 0 96324 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2095
timestamp 1712078602
transform 1 0 96922 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2099
timestamp 1712078602
transform 1 0 97106 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_18_2124
timestamp 1712078602
transform 1 0 98256 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2138
timestamp 1712078602
transform 1 0 98900 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_2150
timestamp 1712078602
transform 1 0 99452 0 1 5984
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2157
timestamp 1712078602
transform 1 0 99774 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2169
timestamp 1712078602
transform 1 0 100326 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2176
timestamp 1712078602
transform 1 0 100648 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_18_2183
timestamp 1712078602
transform 1 0 100970 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_18_2191
timestamp 1712078602
transform 1 0 101338 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_8  FILLER_18_2202
timestamp 1712078602
transform 1 0 101844 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_18_2210
timestamp 1712078602
transform 1 0 102212 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2233
timestamp 1712078602
transform 1 0 103270 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2245
timestamp 1712078602
transform 1 0 103822 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_2257
timestamp 1712078602
transform 1 0 104374 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_18_2265
timestamp 1712078602
transform 1 0 104742 0 1 5984
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2269
timestamp 1712078602
transform 1 0 104926 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2281
timestamp 1712078602
transform 1 0 105478 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2293
timestamp 1712078602
transform 1 0 106030 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2305
timestamp 1712078602
transform 1 0 106582 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_2317
timestamp 1712078602
transform 1 0 107134 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2323
timestamp 1712078602
transform 1 0 107410 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2325
timestamp 1712078602
transform 1 0 107502 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2337
timestamp 1712078602
transform 1 0 108054 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2349
timestamp 1712078602
transform 1 0 108606 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2361
timestamp 1712078602
transform 1 0 109158 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_2373
timestamp 1712078602
transform 1 0 109710 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2379
timestamp 1712078602
transform 1 0 109986 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2381
timestamp 1712078602
transform 1 0 110078 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2393
timestamp 1712078602
transform 1 0 110630 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2405
timestamp 1712078602
transform 1 0 111182 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2417
timestamp 1712078602
transform 1 0 111734 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_2429
timestamp 1712078602
transform 1 0 112286 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2435
timestamp 1712078602
transform 1 0 112562 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2437
timestamp 1712078602
transform 1 0 112654 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2449
timestamp 1712078602
transform 1 0 113206 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2481
timestamp 1712078602
transform 1 0 114678 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2488
timestamp 1712078602
transform 1 0 115000 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2493
timestamp 1712078602
transform 1 0 115230 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2497
timestamp 1712078602
transform 1 0 115414 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2507
timestamp 1712078602
transform 1 0 115874 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2514
timestamp 1712078602
transform 1 0 116196 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2526
timestamp 1712078602
transform 1 0 116748 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_2538
timestamp 1712078602
transform 1 0 117300 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_18_2546
timestamp 1712078602
transform 1 0 117668 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2549
timestamp 1712078602
transform 1 0 117806 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2561
timestamp 1712078602
transform 1 0 118358 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_18_2573
timestamp 1712078602
transform 1 0 118910 0 1 5984
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2579
timestamp 1712078602
transform 1 0 119186 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2592
timestamp 1712078602
transform 1 0 119784 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2599
timestamp 1712078602
transform 1 0 120106 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2603
timestamp 1712078602
transform 1 0 120290 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2605
timestamp 1712078602
transform 1 0 120382 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_18_2615
timestamp 1712078602
transform 1 0 120842 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2621
timestamp 1712078602
transform 1 0 121118 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2631
timestamp 1712078602
transform 1 0 121578 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2638
timestamp 1712078602
transform 1 0 121900 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2645
timestamp 1712078602
transform 1 0 122222 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_18_2657
timestamp 1712078602
transform 1 0 122774 0 1 5984
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2661
timestamp 1712078602
transform 1 0 122958 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2673
timestamp 1712078602
transform 1 0 123510 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_2685
timestamp 1712078602
transform 1 0 124062 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2693
timestamp 1712078602
transform 1 0 124430 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2698
timestamp 1712078602
transform 1 0 124660 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_2710
timestamp 1712078602
transform 1 0 125212 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2720
timestamp 1712078602
transform 1 0 125672 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2724
timestamp 1712078602
transform 1 0 125856 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2729
timestamp 1712078602
transform 1 0 126086 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2753
timestamp 1712078602
transform 1 0 127190 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_18_2766
timestamp 1712078602
transform 1 0 127788 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2776
timestamp 1712078602
transform 1 0 128248 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2783
timestamp 1712078602
transform 1 0 128570 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2795
timestamp 1712078602
transform 1 0 129122 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2807
timestamp 1712078602
transform 1 0 129674 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_2819
timestamp 1712078602
transform 1 0 130226 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2827
timestamp 1712078602
transform 1 0 130594 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2829
timestamp 1712078602
transform 1 0 130686 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2844
timestamp 1712078602
transform 1 0 131376 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_18_2856
timestamp 1712078602
transform 1 0 131928 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2860
timestamp 1712078602
transform 1 0 132112 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2867
timestamp 1712078602
transform 1 0 132434 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2880
timestamp 1712078602
transform 1 0 133032 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2905
timestamp 1712078602
transform 1 0 134182 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2929
timestamp 1712078602
transform 1 0 135286 0 1 5984
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_18_2936
timestamp 1712078602
transform 1 0 135608 0 1 5984
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2950
timestamp 1712078602
transform 1 0 136252 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2962
timestamp 1712078602
transform 1 0 136804 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2974
timestamp 1712078602
transform 1 0 137356 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_18_2986
timestamp 1712078602
transform 1 0 137908 0 1 5984
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_18_2994
timestamp 1712078602
transform 1 0 138276 0 1 5984
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_18_2997
timestamp 1712078602
transform 1 0 138414 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3009
timestamp 1712078602
transform 1 0 138966 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3021
timestamp 1712078602
transform 1 0 139518 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3033
timestamp 1712078602
transform 1 0 140070 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_3045
timestamp 1712078602
transform 1 0 140622 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_3051
timestamp 1712078602
transform 1 0 140898 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3053
timestamp 1712078602
transform 1 0 140990 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3065
timestamp 1712078602
transform 1 0 141542 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3077
timestamp 1712078602
transform 1 0 142094 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3089
timestamp 1712078602
transform 1 0 142646 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_3101
timestamp 1712078602
transform 1 0 143198 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_3107
timestamp 1712078602
transform 1 0 143474 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3109
timestamp 1712078602
transform 1 0 143566 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3121
timestamp 1712078602
transform 1 0 144118 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3133
timestamp 1712078602
transform 1 0 144670 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3145
timestamp 1712078602
transform 1 0 145222 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_3157
timestamp 1712078602
transform 1 0 145774 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_3163
timestamp 1712078602
transform 1 0 146050 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3165
timestamp 1712078602
transform 1 0 146142 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3177
timestamp 1712078602
transform 1 0 146694 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3189
timestamp 1712078602
transform 1 0 147246 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3201
timestamp 1712078602
transform 1 0 147798 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_3213
timestamp 1712078602
transform 1 0 148350 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_3219
timestamp 1712078602
transform 1 0 148626 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3221
timestamp 1712078602
transform 1 0 148718 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3233
timestamp 1712078602
transform 1 0 149270 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3245
timestamp 1712078602
transform 1 0 149822 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3257
timestamp 1712078602
transform 1 0 150374 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_3269
timestamp 1712078602
transform 1 0 150926 0 1 5984
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_18_3275
timestamp 1712078602
transform 1 0 151202 0 1 5984
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3277
timestamp 1712078602
transform 1 0 151294 0 1 5984
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_18_3289
timestamp 1712078602
transform 1 0 151846 0 1 5984
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_18_3301
timestamp 1712078602
transform 1 0 152398 0 1 5984
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1712078602
transform 1 0 690 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1712078602
transform 1 0 1242 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1712078602
transform 1 0 1794 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1712078602
transform 1 0 2346 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1712078602
transform 1 0 2898 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1712078602
transform 1 0 3082 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1712078602
transform 1 0 3174 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1712078602
transform 1 0 3726 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1712078602
transform 1 0 4278 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1712078602
transform 1 0 4830 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1712078602
transform 1 0 5382 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1712078602
transform 1 0 5658 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1712078602
transform 1 0 5750 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1712078602
transform 1 0 6302 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1712078602
transform 1 0 6854 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1712078602
transform 1 0 7406 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1712078602
transform 1 0 7958 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1712078602
transform 1 0 8234 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1712078602
transform 1 0 8326 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1712078602
transform 1 0 8878 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1712078602
transform 1 0 9430 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1712078602
transform 1 0 9982 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1712078602
transform 1 0 10534 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1712078602
transform 1 0 10810 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1712078602
transform 1 0 10902 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1712078602
transform 1 0 11454 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1712078602
transform 1 0 12006 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_261
timestamp 1712078602
transform 1 0 12558 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_19_269
timestamp 1712078602
transform 1 0 12926 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1712078602
transform 1 0 13156 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1712078602
transform 1 0 13478 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1712078602
transform 1 0 13662 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1712078602
transform 1 0 14122 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_308
timestamp 1712078602
transform 1 0 14720 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1712078602
transform 1 0 15824 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_357
timestamp 1712078602
transform 1 0 16974 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1712078602
transform 1 0 17572 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_377
timestamp 1712078602
transform 1 0 17894 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_383
timestamp 1712078602
transform 1 0 18170 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1712078602
transform 1 0 18400 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_397
timestamp 1712078602
transform 1 0 18814 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_410
timestamp 1712078602
transform 1 0 19412 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_416
timestamp 1712078602
transform 1 0 19688 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_437
timestamp 1712078602
transform 1 0 20654 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1712078602
transform 1 0 20976 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_452
timestamp 1712078602
transform 1 0 21344 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_465
timestamp 1712078602
transform 1 0 21942 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_471
timestamp 1712078602
transform 1 0 22218 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_475
timestamp 1712078602
transform 1 0 22402 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_487
timestamp 1712078602
transform 1 0 22954 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_499
timestamp 1712078602
transform 1 0 23506 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1712078602
transform 1 0 23690 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1712078602
transform 1 0 23782 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1712078602
transform 1 0 24334 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1712078602
transform 1 0 24886 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1712078602
transform 1 0 25438 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_556
timestamp 1712078602
transform 1 0 26128 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_19_561
timestamp 1712078602
transform 1 0 26358 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_19_566
timestamp 1712078602
transform 1 0 26588 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_579
timestamp 1712078602
transform 1 0 27186 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_603
timestamp 1712078602
transform 1 0 28290 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_611
timestamp 1712078602
transform 1 0 28658 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1712078602
transform 1 0 28842 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_19_617
timestamp 1712078602
transform 1 0 28934 0 -1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1712078602
transform 1 0 29486 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1712078602
transform 1 0 30038 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1712078602
transform 1 0 30590 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1712078602
transform 1 0 31142 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1712078602
transform 1 0 31418 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1712078602
transform 1 0 31510 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1712078602
transform 1 0 32062 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1712078602
transform 1 0 32614 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1712078602
transform 1 0 33166 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1712078602
transform 1 0 33718 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1712078602
transform 1 0 33994 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1712078602
transform 1 0 34086 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1712078602
transform 1 0 34638 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1712078602
transform 1 0 35190 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_765
timestamp 1712078602
transform 1 0 35742 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_771
timestamp 1712078602
transform 1 0 36018 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_19_775
timestamp 1712078602
transform 1 0 36202 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1712078602
transform 1 0 36570 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1712078602
transform 1 0 36662 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_797
timestamp 1712078602
transform 1 0 37214 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_801
timestamp 1712078602
transform 1 0 37398 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_805
timestamp 1712078602
transform 1 0 37582 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_829
timestamp 1712078602
transform 1 0 38686 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_836
timestamp 1712078602
transform 1 0 39008 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_844
timestamp 1712078602
transform 1 0 39376 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_851
timestamp 1712078602
transform 1 0 39698 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_875
timestamp 1712078602
transform 1 0 40802 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_887
timestamp 1712078602
transform 1 0 41354 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1712078602
transform 1 0 41722 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_897
timestamp 1712078602
transform 1 0 41814 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_921
timestamp 1712078602
transform 1 0 42918 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_945
timestamp 1712078602
transform 1 0 44022 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1712078602
transform 1 0 44298 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_953
timestamp 1712078602
transform 1 0 44390 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_966
timestamp 1712078602
transform 1 0 44988 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_974
timestamp 1712078602
transform 1 0 45356 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_981
timestamp 1712078602
transform 1 0 45678 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_993
timestamp 1712078602
transform 1 0 46230 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_19_1005
timestamp 1712078602
transform 1 0 46782 0 -1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1009
timestamp 1712078602
transform 1 0 46966 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1021
timestamp 1712078602
transform 1 0 47518 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1033
timestamp 1712078602
transform 1 0 48070 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1045
timestamp 1712078602
transform 1 0 48622 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1060
timestamp 1712078602
transform 1 0 49312 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1065
timestamp 1712078602
transform 1 0 49542 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1086
timestamp 1712078602
transform 1 0 50508 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_19_1110
timestamp 1712078602
transform 1 0 51612 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1118
timestamp 1712078602
transform 1 0 51980 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_8  FILLER_19_1130
timestamp 1712078602
transform 1 0 52532 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1138
timestamp 1712078602
transform 1 0 52900 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1142
timestamp 1712078602
transform 1 0 53084 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1154
timestamp 1712078602
transform 1 0 53636 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_1166
timestamp 1712078602
transform 1 0 54188 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1174
timestamp 1712078602
transform 1 0 54556 0 -1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1177
timestamp 1712078602
transform 1 0 54694 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1189
timestamp 1712078602
transform 1 0 55246 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_19_1201
timestamp 1712078602
transform 1 0 55798 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1213
timestamp 1712078602
transform 1 0 56350 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1220
timestamp 1712078602
transform 1 0 56672 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1228
timestamp 1712078602
transform 1 0 57040 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1237
timestamp 1712078602
transform 1 0 57454 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1250
timestamp 1712078602
transform 1 0 58052 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1274
timestamp 1712078602
transform 1 0 59156 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_1281
timestamp 1712078602
transform 1 0 59478 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1287
timestamp 1712078602
transform 1 0 59754 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1289
timestamp 1712078602
transform 1 0 59846 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1301
timestamp 1712078602
transform 1 0 60398 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1313
timestamp 1712078602
transform 1 0 60950 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1325
timestamp 1712078602
transform 1 0 61502 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_1337
timestamp 1712078602
transform 1 0 62054 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1343
timestamp 1712078602
transform 1 0 62330 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1345
timestamp 1712078602
transform 1 0 62422 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_1357
timestamp 1712078602
transform 1 0 62974 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1368
timestamp 1712078602
transform 1 0 63480 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1376
timestamp 1712078602
transform 1 0 63848 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1383
timestamp 1712078602
transform 1 0 64170 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1396
timestamp 1712078602
transform 1 0 64768 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1401
timestamp 1712078602
transform 1 0 64998 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1406
timestamp 1712078602
transform 1 0 65228 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1430
timestamp 1712078602
transform 1 0 66332 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1434
timestamp 1712078602
transform 1 0 66516 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1444
timestamp 1712078602
transform 1 0 66976 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1451
timestamp 1712078602
transform 1 0 67298 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1455
timestamp 1712078602
transform 1 0 67482 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1457
timestamp 1712078602
transform 1 0 67574 0 -1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1463
timestamp 1712078602
transform 1 0 67850 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1475
timestamp 1712078602
transform 1 0 68402 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1487
timestamp 1712078602
transform 1 0 68954 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1499
timestamp 1712078602
transform 1 0 69506 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1511
timestamp 1712078602
transform 1 0 70058 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1513
timestamp 1712078602
transform 1 0 70150 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1525
timestamp 1712078602
transform 1 0 70702 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1537
timestamp 1712078602
transform 1 0 71254 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1541
timestamp 1712078602
transform 1 0 71438 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1548
timestamp 1712078602
transform 1 0 71760 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_1560
timestamp 1712078602
transform 1 0 72312 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_6  FILLER_19_1578
timestamp 1712078602
transform 1 0 73140 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1587
timestamp 1712078602
transform 1 0 73554 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_1611
timestamp 1712078602
transform 1 0 74658 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1620
timestamp 1712078602
transform 1 0 75072 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1625
timestamp 1712078602
transform 1 0 75302 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1629
timestamp 1712078602
transform 1 0 75486 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1639
timestamp 1712078602
transform 1 0 75946 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1645
timestamp 1712078602
transform 1 0 76222 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1649
timestamp 1712078602
transform 1 0 76406 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1653
timestamp 1712078602
transform 1 0 76590 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1657
timestamp 1712078602
transform 1 0 76774 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1661
timestamp 1712078602
transform 1 0 76958 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1665
timestamp 1712078602
transform 1 0 77142 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1676
timestamp 1712078602
transform 1 0 77648 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1681
timestamp 1712078602
transform 1 0 77878 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1685
timestamp 1712078602
transform 1 0 78062 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1689
timestamp 1712078602
transform 1 0 78246 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1693
timestamp 1712078602
transform 1 0 78430 0 -1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1697
timestamp 1712078602
transform 1 0 78614 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1709
timestamp 1712078602
transform 1 0 79166 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1713
timestamp 1712078602
transform 1 0 79350 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1723
timestamp 1712078602
transform 1 0 79810 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1731
timestamp 1712078602
transform 1 0 80178 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1735
timestamp 1712078602
transform 1 0 80362 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_19_1737
timestamp 1712078602
transform 1 0 80454 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1743
timestamp 1712078602
transform 1 0 80730 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1767
timestamp 1712078602
transform 1 0 81834 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1780
timestamp 1712078602
transform 1 0 82432 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1788
timestamp 1712078602
transform 1 0 82800 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1793
timestamp 1712078602
transform 1 0 83030 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1801
timestamp 1712078602
transform 1 0 83398 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1808
timestamp 1712078602
transform 1 0 83720 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1815
timestamp 1712078602
transform 1 0 84042 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1827
timestamp 1712078602
transform 1 0 84594 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_1839
timestamp 1712078602
transform 1 0 85146 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1847
timestamp 1712078602
transform 1 0 85514 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1849
timestamp 1712078602
transform 1 0 85606 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1861
timestamp 1712078602
transform 1 0 86158 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1873
timestamp 1712078602
transform 1 0 86710 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1885
timestamp 1712078602
transform 1 0 87262 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_1889
timestamp 1712078602
transform 1 0 87446 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1893
timestamp 1712078602
transform 1 0 87630 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1900
timestamp 1712078602
transform 1 0 87952 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1925
timestamp 1712078602
transform 1 0 89102 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1949
timestamp 1712078602
transform 1 0 90206 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1956
timestamp 1712078602
transform 1 0 90528 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_1964
timestamp 1712078602
transform 1 0 90896 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1971
timestamp 1712078602
transform 1 0 91218 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1983
timestamp 1712078602
transform 1 0 91770 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_1995
timestamp 1712078602
transform 1 0 92322 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2007
timestamp 1712078602
transform 1 0 92874 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2015
timestamp 1712078602
transform 1 0 93242 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2017
timestamp 1712078602
transform 1 0 93334 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2029
timestamp 1712078602
transform 1 0 93886 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2033
timestamp 1712078602
transform 1 0 94070 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2041
timestamp 1712078602
transform 1 0 94438 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2049
timestamp 1712078602
transform 1 0 94806 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_19_2057
timestamp 1712078602
transform 1 0 95174 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2068
timestamp 1712078602
transform 1 0 95680 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2082
timestamp 1712078602
transform 1 0 96324 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2109
timestamp 1712078602
transform 1 0 97566 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_2122
timestamp 1712078602
transform 1 0 98164 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_2  FILLER_19_2138
timestamp 1712078602
transform 1 0 98900 0 -1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2145
timestamp 1712078602
transform 1 0 99222 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2157
timestamp 1712078602
transform 1 0 99774 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_19_2165
timestamp 1712078602
transform 1 0 100142 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2170
timestamp 1712078602
transform 1 0 100372 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_2177
timestamp 1712078602
transform 1 0 100694 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2183
timestamp 1712078602
transform 1 0 100970 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2185
timestamp 1712078602
transform 1 0 101062 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2189
timestamp 1712078602
transform 1 0 101246 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2210
timestamp 1712078602
transform 1 0 102212 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_19_2234
timestamp 1712078602
transform 1 0 103316 0 -1 6528
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2244
timestamp 1712078602
transform 1 0 103776 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2256
timestamp 1712078602
transform 1 0 104328 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2268
timestamp 1712078602
transform 1 0 104880 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2280
timestamp 1712078602
transform 1 0 105432 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2292
timestamp 1712078602
transform 1 0 105984 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2297
timestamp 1712078602
transform 1 0 106214 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2309
timestamp 1712078602
transform 1 0 106766 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2321
timestamp 1712078602
transform 1 0 107318 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2333
timestamp 1712078602
transform 1 0 107870 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_2345
timestamp 1712078602
transform 1 0 108422 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2351
timestamp 1712078602
transform 1 0 108698 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2353
timestamp 1712078602
transform 1 0 108790 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2365
timestamp 1712078602
transform 1 0 109342 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2377
timestamp 1712078602
transform 1 0 109894 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2389
timestamp 1712078602
transform 1 0 110446 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_2401
timestamp 1712078602
transform 1 0 110998 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2407
timestamp 1712078602
transform 1 0 111274 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2409
timestamp 1712078602
transform 1 0 111366 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2421
timestamp 1712078602
transform 1 0 111918 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2433
timestamp 1712078602
transform 1 0 112470 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2445
timestamp 1712078602
transform 1 0 113022 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2449
timestamp 1712078602
transform 1 0 113206 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2453
timestamp 1712078602
transform 1 0 113390 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2460
timestamp 1712078602
transform 1 0 113712 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2485
timestamp 1712078602
transform 1 0 114862 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2492
timestamp 1712078602
transform 1 0 115184 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2516
timestamp 1712078602
transform 1 0 116288 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2524
timestamp 1712078602
transform 1 0 116656 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2536
timestamp 1712078602
transform 1 0 117208 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2548
timestamp 1712078602
transform 1 0 117760 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_19_2560
timestamp 1712078602
transform 1 0 118312 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2565
timestamp 1712078602
transform 1 0 118542 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2572
timestamp 1712078602
transform 1 0 118864 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_19_2577
timestamp 1712078602
transform 1 0 119094 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2600
timestamp 1712078602
transform 1 0 120152 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2624
timestamp 1712078602
transform 1 0 121256 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2633
timestamp 1712078602
transform 1 0 121670 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2641
timestamp 1712078602
transform 1 0 122038 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2649
timestamp 1712078602
transform 1 0 122406 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2656
timestamp 1712078602
transform 1 0 122728 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2668
timestamp 1712078602
transform 1 0 123280 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2680
timestamp 1712078602
transform 1 0 123832 0 -1 6528
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2689
timestamp 1712078602
transform 1 0 124246 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_2701
timestamp 1712078602
transform 1 0 124798 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2710
timestamp 1712078602
transform 1 0 125212 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2718
timestamp 1712078602
transform 1 0 125580 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2723
timestamp 1712078602
transform 1 0 125810 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2736
timestamp 1712078602
transform 1 0 126408 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2765
timestamp 1712078602
transform 1 0 127742 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2778
timestamp 1712078602
transform 1 0 128340 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2785
timestamp 1712078602
transform 1 0 128662 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_19_2797
timestamp 1712078602
transform 1 0 129214 0 -1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2801
timestamp 1712078602
transform 1 0 129398 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2813
timestamp 1712078602
transform 1 0 129950 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_2825
timestamp 1712078602
transform 1 0 130502 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2831
timestamp 1712078602
transform 1 0 130778 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2836
timestamp 1712078602
transform 1 0 131008 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2844
timestamp 1712078602
transform 1 0 131376 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2852
timestamp 1712078602
transform 1 0 131744 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2860
timestamp 1712078602
transform 1 0 132112 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2867
timestamp 1712078602
transform 1 0 132434 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2891
timestamp 1712078602
transform 1 0 133538 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2904
timestamp 1712078602
transform 1 0 134136 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2933
timestamp 1712078602
transform 1 0 135470 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_19_2946
timestamp 1712078602
transform 1 0 136068 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_19_2959
timestamp 1712078602
transform 1 0 136666 0 -1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_19_2967
timestamp 1712078602
transform 1 0 137034 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2969
timestamp 1712078602
transform 1 0 137126 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2981
timestamp 1712078602
transform 1 0 137678 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_2993
timestamp 1712078602
transform 1 0 138230 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3005
timestamp 1712078602
transform 1 0 138782 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_3017
timestamp 1712078602
transform 1 0 139334 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_3023
timestamp 1712078602
transform 1 0 139610 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3025
timestamp 1712078602
transform 1 0 139702 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3037
timestamp 1712078602
transform 1 0 140254 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3049
timestamp 1712078602
transform 1 0 140806 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3061
timestamp 1712078602
transform 1 0 141358 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_3073
timestamp 1712078602
transform 1 0 141910 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_3079
timestamp 1712078602
transform 1 0 142186 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3081
timestamp 1712078602
transform 1 0 142278 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3093
timestamp 1712078602
transform 1 0 142830 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3105
timestamp 1712078602
transform 1 0 143382 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3117
timestamp 1712078602
transform 1 0 143934 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_3129
timestamp 1712078602
transform 1 0 144486 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_3135
timestamp 1712078602
transform 1 0 144762 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3137
timestamp 1712078602
transform 1 0 144854 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3149
timestamp 1712078602
transform 1 0 145406 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3161
timestamp 1712078602
transform 1 0 145958 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3173
timestamp 1712078602
transform 1 0 146510 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_3185
timestamp 1712078602
transform 1 0 147062 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_3191
timestamp 1712078602
transform 1 0 147338 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3193
timestamp 1712078602
transform 1 0 147430 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3205
timestamp 1712078602
transform 1 0 147982 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3217
timestamp 1712078602
transform 1 0 148534 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3229
timestamp 1712078602
transform 1 0 149086 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_19_3241
timestamp 1712078602
transform 1 0 149638 0 -1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_19_3247
timestamp 1712078602
transform 1 0 149914 0 -1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3249
timestamp 1712078602
transform 1 0 150006 0 -1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3261
timestamp 1712078602
transform 1 0 150558 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_3273
timestamp 1712078602
transform 1 0 151110 0 -1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_19_3280
timestamp 1712078602
transform 1 0 151432 0 -1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_19_3292
timestamp 1712078602
transform 1 0 151984 0 -1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_19_3296
timestamp 1712078602
transform 1 0 152168 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_19_3300
timestamp 1712078602
transform 1 0 152352 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_19_3305
timestamp 1712078602
transform 1 0 152582 0 -1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1712078602
transform 1 0 690 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1712078602
transform 1 0 920 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1712078602
transform 1 0 1472 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1712078602
transform 1 0 1886 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_20_37
timestamp 1712078602
transform 1 0 2254 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1712078602
transform 1 0 2438 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1712078602
transform 1 0 2990 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_57
timestamp 1712078602
transform 1 0 3174 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1712078602
transform 1 0 3726 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_8  FILLER_20_74
timestamp 1712078602
transform 1 0 3956 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1712078602
transform 1 0 4324 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1712078602
transform 1 0 4462 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1712078602
transform 1 0 5014 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1712078602
transform 1 0 5520 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_113
timestamp 1712078602
transform 1 0 5750 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_125
timestamp 1712078602
transform 1 0 6302 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1712078602
transform 1 0 6854 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_144
timestamp 1712078602
transform 1 0 7176 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_156
timestamp 1712078602
transform 1 0 7728 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_169
timestamp 1712078602
transform 1 0 8326 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_174
timestamp 1712078602
transform 1 0 8556 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1712078602
transform 1 0 9108 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1712078602
transform 1 0 9476 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1712078602
transform 1 0 9614 0 1 6528
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_20_208
timestamp 1712078602
transform 1 0 10120 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1712078602
transform 1 0 10672 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_225
timestamp 1712078602
transform 1 0 10902 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_20_237
timestamp 1712078602
transform 1 0 11454 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_20_241
timestamp 1712078602
transform 1 0 11638 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1712078602
transform 1 0 12006 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1712078602
transform 1 0 12190 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_265
timestamp 1712078602
transform 1 0 12742 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1712078602
transform 1 0 13248 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_281
timestamp 1712078602
transform 1 0 13478 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1712078602
transform 1 0 14536 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1712078602
transform 1 0 14766 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1712078602
transform 1 0 15824 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_337
timestamp 1712078602
transform 1 0 16054 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1712078602
transform 1 0 17112 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_385
timestamp 1712078602
transform 1 0 18262 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_391
timestamp 1712078602
transform 1 0 18538 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_20_393
timestamp 1712078602
transform 1 0 18630 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1712078602
transform 1 0 19688 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_421
timestamp 1712078602
transform 1 0 19918 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_444
timestamp 1712078602
transform 1 0 20976 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_449
timestamp 1712078602
transform 1 0 21206 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_470
timestamp 1712078602
transform 1 0 22172 0 1 6528
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_20_486
timestamp 1712078602
transform 1 0 22908 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_498
timestamp 1712078602
transform 1 0 23460 0 1 6528
box -19 -24 295 296
use sky130_ef_sc_hd__decap_12  FILLER_20_508
timestamp 1712078602
transform 1 0 23920 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_520
timestamp 1712078602
transform 1 0 24472 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_533
timestamp 1712078602
transform 1 0 25070 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_538
timestamp 1712078602
transform 1 0 25300 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_551
timestamp 1712078602
transform 1 0 25898 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_20_559
timestamp 1712078602
transform 1 0 26266 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_20_561
timestamp 1712078602
transform 1 0 26358 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_584
timestamp 1712078602
transform 1 0 27416 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_589
timestamp 1712078602
transform 1 0 27646 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_612
timestamp 1712078602
transform 1 0 28704 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1712078602
transform 1 0 29854 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1712078602
transform 1 0 30130 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_648
timestamp 1712078602
transform 1 0 30360 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_660
timestamp 1712078602
transform 1 0 30912 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_676
timestamp 1712078602
transform 1 0 31648 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_688
timestamp 1712078602
transform 1 0 32200 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_701
timestamp 1712078602
transform 1 0 32798 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_708
timestamp 1712078602
transform 1 0 33120 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_720
timestamp 1712078602
transform 1 0 33672 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_8  FILLER_20_729
timestamp 1712078602
transform 1 0 34086 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_737
timestamp 1712078602
transform 1 0 34454 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_742
timestamp 1712078602
transform 1 0 34684 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_754
timestamp 1712078602
transform 1 0 35236 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1712078602
transform 1 0 35374 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_769
timestamp 1712078602
transform 1 0 35926 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_780
timestamp 1712078602
transform 1 0 36432 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_785
timestamp 1712078602
transform 1 0 36662 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_808
timestamp 1712078602
transform 1 0 37720 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_813
timestamp 1712078602
transform 1 0 37950 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_836
timestamp 1712078602
transform 1 0 39008 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1712078602
transform 1 0 40158 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1712078602
transform 1 0 40434 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_878
timestamp 1712078602
transform 1 0 40940 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_885
timestamp 1712078602
transform 1 0 41262 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_892
timestamp 1712078602
transform 1 0 41584 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_897
timestamp 1712078602
transform 1 0 41814 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_920
timestamp 1712078602
transform 1 0 42872 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_925
timestamp 1712078602
transform 1 0 43102 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_948
timestamp 1712078602
transform 1 0 44160 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_973
timestamp 1712078602
transform 1 0 45310 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_979
timestamp 1712078602
transform 1 0 45586 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_981
timestamp 1712078602
transform 1 0 45678 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_989
timestamp 1712078602
transform 1 0 46046 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1001
timestamp 1712078602
transform 1 0 46598 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1007
timestamp 1712078602
transform 1 0 46874 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1012
timestamp 1712078602
transform 1 0 47104 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1024
timestamp 1712078602
transform 1 0 47656 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_1037
timestamp 1712078602
transform 1 0 48254 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1042
timestamp 1712078602
transform 1 0 48484 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1057
timestamp 1712078602
transform 1 0 49174 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1063
timestamp 1712078602
transform 1 0 49450 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1065
timestamp 1712078602
transform 1 0 49542 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1088
timestamp 1712078602
transform 1 0 50600 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1093
timestamp 1712078602
transform 1 0 50830 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1116
timestamp 1712078602
transform 1 0 51888 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1141
timestamp 1712078602
transform 1 0 53038 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1712078602
transform 1 0 53314 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1149
timestamp 1712078602
transform 1 0 53406 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1161
timestamp 1712078602
transform 1 0 53958 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1173
timestamp 1712078602
transform 1 0 54510 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1180
timestamp 1712078602
transform 1 0 54832 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1192
timestamp 1712078602
transform 1 0 55384 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1196
timestamp 1712078602
transform 1 0 55568 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1200
timestamp 1712078602
transform 1 0 55752 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1205
timestamp 1712078602
transform 1 0 55982 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1228
timestamp 1712078602
transform 1 0 57040 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1233
timestamp 1712078602
transform 1 0 57270 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1256
timestamp 1712078602
transform 1 0 58328 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1261
timestamp 1712078602
transform 1 0 58558 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1284
timestamp 1712078602
transform 1 0 59616 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1298
timestamp 1712078602
transform 1 0 60260 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1309
timestamp 1712078602
transform 1 0 60766 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1315
timestamp 1712078602
transform 1 0 61042 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1317
timestamp 1712078602
transform 1 0 61134 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1329
timestamp 1712078602
transform 1 0 61686 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1340
timestamp 1712078602
transform 1 0 62192 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1345
timestamp 1712078602
transform 1 0 62422 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1355
timestamp 1712078602
transform 1 0 62882 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1368
timestamp 1712078602
transform 1 0 63480 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1373
timestamp 1712078602
transform 1 0 63710 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1394
timestamp 1712078602
transform 1 0 64676 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1401
timestamp 1712078602
transform 1 0 64998 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1424
timestamp 1712078602
transform 1 0 66056 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1449
timestamp 1712078602
transform 1 0 67206 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1455
timestamp 1712078602
transform 1 0 67482 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1457
timestamp 1712078602
transform 1 0 67574 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1469
timestamp 1712078602
transform 1 0 68126 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1476
timestamp 1712078602
transform 1 0 68448 0 1 6528
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1485
timestamp 1712078602
transform 1 0 68862 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1497
timestamp 1712078602
transform 1 0 69414 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1509
timestamp 1712078602
transform 1 0 69966 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1516
timestamp 1712078602
transform 1 0 70288 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1528
timestamp 1712078602
transform 1 0 70840 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1544
timestamp 1712078602
transform 1 0 71576 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1556
timestamp 1712078602
transform 1 0 72128 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1560
timestamp 1712078602
transform 1 0 72312 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1564
timestamp 1712078602
transform 1 0 72496 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1569
timestamp 1712078602
transform 1 0 72726 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1592
timestamp 1712078602
transform 1 0 73784 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1620
timestamp 1712078602
transform 1 0 75072 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1625
timestamp 1712078602
transform 1 0 75302 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1648
timestamp 1712078602
transform 1 0 76360 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1653
timestamp 1712078602
transform 1 0 76590 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1676
timestamp 1712078602
transform 1 0 77648 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1684
timestamp 1712078602
transform 1 0 78016 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1691
timestamp 1712078602
transform 1 0 78338 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_1699
timestamp 1712078602
transform 1 0 78706 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1704
timestamp 1712078602
transform 1 0 78936 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1709
timestamp 1712078602
transform 1 0 79166 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1732
timestamp 1712078602
transform 1 0 80224 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1757
timestamp 1712078602
transform 1 0 81374 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1763
timestamp 1712078602
transform 1 0 81650 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1785
timestamp 1712078602
transform 1 0 82662 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1791
timestamp 1712078602
transform 1 0 82938 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1802
timestamp 1712078602
transform 1 0 83444 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1810
timestamp 1712078602
transform 1 0 83812 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_1818
timestamp 1712078602
transform 1 0 84180 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1821
timestamp 1712078602
transform 1 0 84318 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1833
timestamp 1712078602
transform 1 0 84870 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1839
timestamp 1712078602
transform 1 0 85146 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1843
timestamp 1712078602
transform 1 0 85330 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1847
timestamp 1712078602
transform 1 0 85514 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1849
timestamp 1712078602
transform 1 0 85606 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1861
timestamp 1712078602
transform 1 0 86158 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1872
timestamp 1712078602
transform 1 0 86664 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1886
timestamp 1712078602
transform 1 0 87308 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_1894
timestamp 1712078602
transform 1 0 87676 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1900
timestamp 1712078602
transform 1 0 87952 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1925
timestamp 1712078602
transform 1 0 89102 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1931
timestamp 1712078602
transform 1 0 89378 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_1953
timestamp 1712078602
transform 1 0 90390 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_1959
timestamp 1712078602
transform 1 0 90666 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_1970
timestamp 1712078602
transform 1 0 91172 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_1977
timestamp 1712078602
transform 1 0 91494 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_20_1985
timestamp 1712078602
transform 1 0 91862 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_1989
timestamp 1712078602
transform 1 0 92046 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2001
timestamp 1712078602
transform 1 0 92598 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2010
timestamp 1712078602
transform 1 0 93012 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2017
timestamp 1712078602
transform 1 0 93334 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2023
timestamp 1712078602
transform 1 0 93610 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2027
timestamp 1712078602
transform 1 0 93794 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2040
timestamp 1712078602
transform 1 0 94392 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_2045
timestamp 1712078602
transform 1 0 94622 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2068
timestamp 1712078602
transform 1 0 95680 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2096
timestamp 1712078602
transform 1 0 96968 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2124
timestamp 1712078602
transform 1 0 98256 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2129
timestamp 1712078602
transform 1 0 98486 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2137
timestamp 1712078602
transform 1 0 98854 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_20_2140
timestamp 1712078602
transform 1 0 98992 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2151
timestamp 1712078602
transform 1 0 99498 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2155
timestamp 1712078602
transform 1 0 99682 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_20_2157
timestamp 1712078602
transform 1 0 99774 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2163
timestamp 1712078602
transform 1 0 100050 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2176
timestamp 1712078602
transform 1 0 100648 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2205
timestamp 1712078602
transform 1 0 101982 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2211
timestamp 1712078602
transform 1 0 102258 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2233
timestamp 1712078602
transform 1 0 103270 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2239
timestamp 1712078602
transform 1 0 103546 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2250
timestamp 1712078602
transform 1 0 104052 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2262
timestamp 1712078602
transform 1 0 104604 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2269
timestamp 1712078602
transform 1 0 104926 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2273
timestamp 1712078602
transform 1 0 105110 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2277
timestamp 1712078602
transform 1 0 105294 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2289
timestamp 1712078602
transform 1 0 105846 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2295
timestamp 1712078602
transform 1 0 106122 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2297
timestamp 1712078602
transform 1 0 106214 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_2305
timestamp 1712078602
transform 1 0 106582 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2310
timestamp 1712078602
transform 1 0 106812 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_2322
timestamp 1712078602
transform 1 0 107364 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2325
timestamp 1712078602
transform 1 0 107502 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_2337
timestamp 1712078602
transform 1 0 108054 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2343
timestamp 1712078602
transform 1 0 108330 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2351
timestamp 1712078602
transform 1 0 108698 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2353
timestamp 1712078602
transform 1 0 108790 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2365
timestamp 1712078602
transform 1 0 109342 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_2377
timestamp 1712078602
transform 1 0 109894 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2384
timestamp 1712078602
transform 1 0 110216 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2396
timestamp 1712078602
transform 1 0 110768 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2412
timestamp 1712078602
transform 1 0 111504 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2418
timestamp 1712078602
transform 1 0 111780 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2428
timestamp 1712078602
transform 1 0 112240 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2437
timestamp 1712078602
transform 1 0 112654 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2444
timestamp 1712078602
transform 1 0 112976 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2450
timestamp 1712078602
transform 1 0 113252 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2460
timestamp 1712078602
transform 1 0 113712 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2485
timestamp 1712078602
transform 1 0 114862 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2491
timestamp 1712078602
transform 1 0 115138 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2513
timestamp 1712078602
transform 1 0 116150 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2519
timestamp 1712078602
transform 1 0 116426 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2524
timestamp 1712078602
transform 1 0 116656 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2531
timestamp 1712078602
transform 1 0 116978 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_2539
timestamp 1712078602
transform 1 0 117346 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2544
timestamp 1712078602
transform 1 0 117576 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2549
timestamp 1712078602
transform 1 0 117806 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2570
timestamp 1712078602
transform 1 0 118772 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2597
timestamp 1712078602
transform 1 0 120014 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2603
timestamp 1712078602
transform 1 0 120290 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2625
timestamp 1712078602
transform 1 0 121302 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2631
timestamp 1712078602
transform 1 0 121578 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2653
timestamp 1712078602
transform 1 0 122590 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2659
timestamp 1712078602
transform 1 0 122866 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2661
timestamp 1712078602
transform 1 0 122958 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2673
timestamp 1712078602
transform 1 0 123510 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2677
timestamp 1712078602
transform 1 0 123694 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_20_2685
timestamp 1712078602
transform 1 0 124062 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2689
timestamp 1712078602
transform 1 0 124246 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_20_2697
timestamp 1712078602
transform 1 0 124614 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2709
timestamp 1712078602
transform 1 0 125166 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2715
timestamp 1712078602
transform 1 0 125442 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2737
timestamp 1712078602
transform 1 0 126454 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2743
timestamp 1712078602
transform 1 0 126730 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2765
timestamp 1712078602
transform 1 0 127742 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2771
timestamp 1712078602
transform 1 0 128018 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2793
timestamp 1712078602
transform 1 0 129030 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2799
timestamp 1712078602
transform 1 0 129306 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2801
timestamp 1712078602
transform 1 0 129398 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2807
timestamp 1712078602
transform 1 0 129674 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2811
timestamp 1712078602
transform 1 0 129858 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2823
timestamp 1712078602
transform 1 0 130410 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2827
timestamp 1712078602
transform 1 0 130594 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2829
timestamp 1712078602
transform 1 0 130686 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2837
timestamp 1712078602
transform 1 0 131054 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2852
timestamp 1712078602
transform 1 0 131744 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_3  FILLER_20_2857
timestamp 1712078602
transform 1 0 131974 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2880
timestamp 1712078602
transform 1 0 133032 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2908
timestamp 1712078602
transform 1 0 134320 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2933
timestamp 1712078602
transform 1 0 135470 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2939
timestamp 1712078602
transform 1 0 135746 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_20_2961
timestamp 1712078602
transform 1 0 136758 0 1 6528
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2967
timestamp 1712078602
transform 1 0 137034 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2972
timestamp 1712078602
transform 1 0 137264 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_2979
timestamp 1712078602
transform 1 0 137586 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_2991
timestamp 1712078602
transform 1 0 138138 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_20_2995
timestamp 1712078602
transform 1 0 138322 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_20_2997
timestamp 1712078602
transform 1 0 138414 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_20_3005
timestamp 1712078602
transform 1 0 138782 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3011
timestamp 1712078602
transform 1 0 139058 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_20_3023
timestamp 1712078602
transform 1 0 139610 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3025
timestamp 1712078602
transform 1 0 139702 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_3037
timestamp 1712078602
transform 1 0 140254 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__decap_8  FILLER_20_3044
timestamp 1712078602
transform 1 0 140576 0 1 6528
box -19 -24 387 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3053
timestamp 1712078602
transform 1 0 140990 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3065
timestamp 1712078602
transform 1 0 141542 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_3077
timestamp 1712078602
transform 1 0 142094 0 1 6528
box -19 -24 157 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3084
timestamp 1712078602
transform 1 0 142416 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3096
timestamp 1712078602
transform 1 0 142968 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3112
timestamp 1712078602
transform 1 0 143704 0 1 6528
box -19 -24 571 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3124
timestamp 1712078602
transform 1 0 144256 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_4  FILLER_20_3137
timestamp 1712078602
transform 1 0 144854 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3144
timestamp 1712078602
transform 1 0 145176 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_3156
timestamp 1712078602
transform 1 0 145728 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_8  FILLER_20_3165
timestamp 1712078602
transform 1 0 146142 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3173
timestamp 1712078602
transform 1 0 146510 0 1 6528
box -19 -24 111 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3178
timestamp 1712078602
transform 1 0 146740 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3190
timestamp 1712078602
transform 1 0 147292 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_8  FILLER_20_3193
timestamp 1712078602
transform 1 0 147430 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  FILLER_20_3201
timestamp 1712078602
transform 1 0 147798 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3206
timestamp 1712078602
transform 1 0 148028 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_8  FILLER_20_3211
timestamp 1712078602
transform 1 0 148258 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__fill_1  FILLER_20_3219
timestamp 1712078602
transform 1 0 148626 0 1 6528
box -19 -24 65 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3221
timestamp 1712078602
transform 1 0 148718 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_20_3233
timestamp 1712078602
transform 1 0 149270 0 1 6528
box -19 -24 387 296
use sky130_fd_sc_hd__decap_4  FILLER_20_3244
timestamp 1712078602
transform 1 0 149776 0 1 6528
box -19 -24 203 296
use sky130_ef_sc_hd__decap_12  FILLER_20_3249
timestamp 1712078602
transform 1 0 150006 0 1 6528
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_20_3261
timestamp 1712078602
transform 1 0 150558 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3266
timestamp 1712078602
transform 1 0 150788 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3270
timestamp 1712078602
transform 1 0 150972 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3274
timestamp 1712078602
transform 1 0 151156 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__decap_4  FILLER_20_3277
timestamp 1712078602
transform 1 0 151294 0 1 6528
box -19 -24 203 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3283
timestamp 1712078602
transform 1 0 151570 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3287
timestamp 1712078602
transform 1 0 151754 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3300
timestamp 1712078602
transform 1 0 152352 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_20_3305
timestamp 1712078602
transform 1 0 152582 0 1 6528
box -19 -24 111 296
use sky130_fd_sc_hd__clkbuf_8  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 151846 0 1 6528
box -19 -24 525 296
use sky130_fd_sc_hd__buf_6  input2
timestamp 1712078602
transform 1 0 151938 0 -1 3264
box -19 -24 433 296
use sky130_fd_sc_hd__buf_6  input3
timestamp 1712078602
transform 1 0 152168 0 1 4896
box -19 -24 433 296
use sky130_fd_sc_hd__clkbuf_1  output4
timestamp 1712078602
transform 1 0 782 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output5
timestamp 1712078602
transform 1 0 16422 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1712078602
transform 1 0 17756 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output7
timestamp 1712078602
transform 1 0 19182 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output8
timestamp 1712078602
transform 1 0 21114 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output9
timestamp 1712078602
transform 1 0 22264 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1712078602
transform 1 0 23782 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1712078602
transform 1 0 25162 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1712078602
transform 1 0 26818 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1712078602
transform 1 0 28658 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output14
timestamp 1712078602
transform 1 0 30222 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output15
timestamp 1712078602
transform 1 0 2300 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output16
timestamp 1712078602
transform 1 0 31510 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1712078602
transform 1 0 32982 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output18
timestamp 1712078602
transform 1 0 34546 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output19
timestamp 1712078602
transform 1 0 36064 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1712078602
transform 1 0 37582 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1712078602
transform 1 0 39238 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output22
timestamp 1712078602
transform 1 0 41124 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1712078602
transform 1 0 42182 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output24
timestamp 1712078602
transform 1 0 44712 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output25
timestamp 1712078602
transform 1 0 45540 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output26
timestamp 1712078602
transform 1 0 3818 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output27
timestamp 1712078602
transform 1 0 46966 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output28
timestamp 1712078602
transform 1 0 48346 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output29
timestamp 1712078602
transform 1 0 49174 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output30
timestamp 1712078602
transform 1 0 51428 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output31
timestamp 1712078602
transform 1 0 52946 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output32
timestamp 1712078602
transform 1 0 54694 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output33
timestamp 1712078602
transform 1 0 55614 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output34
timestamp 1712078602
transform 1 0 56856 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output35
timestamp 1712078602
transform 1 0 59340 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output36
timestamp 1712078602
transform 1 0 60628 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1712078602
transform 1 0 5382 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1712078602
transform 1 0 62054 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output39
timestamp 1712078602
transform 1 0 63342 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output40
timestamp 1712078602
transform 1 0 65228 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output41
timestamp 1712078602
transform 1 0 67160 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output42
timestamp 1712078602
transform 1 0 68310 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output43
timestamp 1712078602
transform 1 0 70150 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1712078602
transform 1 0 71438 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1712078602
transform 1 0 72358 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1712078602
transform 1 0 73416 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1712078602
transform 1 0 75992 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output48
timestamp 1712078602
transform 1 0 7038 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output49
timestamp 1712078602
transform 1 0 77878 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output50
timestamp 1712078602
transform 1 0 78798 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output51
timestamp 1712078602
transform 1 0 80776 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output52
timestamp 1712078602
transform 1 0 83582 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output53
timestamp 1712078602
transform 1 0 83904 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output54
timestamp 1712078602
transform 1 0 85192 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output55
timestamp 1712078602
transform 1 0 86526 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output56
timestamp 1712078602
transform 1 0 87952 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output57
timestamp 1712078602
transform 1 0 90666 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output58
timestamp 1712078602
transform 1 0 91356 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output59
timestamp 1712078602
transform 1 0 8418 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output60
timestamp 1712078602
transform 1 0 92874 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output61
timestamp 1712078602
transform 1 0 93932 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output62
timestamp 1712078602
transform 1 0 95910 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output63
timestamp 1712078602
transform 1 0 97796 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output64
timestamp 1712078602
transform 1 0 99084 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output65
timestamp 1712078602
transform 1 0 100556 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output66
timestamp 1712078602
transform 1 0 102350 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output67
timestamp 1712078602
transform 1 0 103638 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output68
timestamp 1712078602
transform 1 0 105156 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output69
timestamp 1712078602
transform 1 0 106674 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output70
timestamp 1712078602
transform 1 0 9982 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output71
timestamp 1712078602
transform 1 0 108192 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output72
timestamp 1712078602
transform 1 0 110078 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output73
timestamp 1712078602
transform 1 0 111366 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output74
timestamp 1712078602
transform 1 0 112838 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output75
timestamp 1712078602
transform 1 0 114862 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output76
timestamp 1712078602
transform 1 0 116840 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output77
timestamp 1712078602
transform 1 0 117438 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output78
timestamp 1712078602
transform 1 0 118726 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output79
timestamp 1712078602
transform 1 0 121164 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output80
timestamp 1712078602
transform 1 0 122084 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output81
timestamp 1712078602
transform 1 0 11500 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output82
timestamp 1712078602
transform 1 0 123556 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output83
timestamp 1712078602
transform 1 0 125074 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output84
timestamp 1712078602
transform 1 0 127190 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output85
timestamp 1712078602
transform 1 0 128432 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output86
timestamp 1712078602
transform 1 0 129720 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output87
timestamp 1712078602
transform 1 0 131238 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output88
timestamp 1712078602
transform 1 0 132756 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output89
timestamp 1712078602
transform 1 0 134504 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output90
timestamp 1712078602
transform 1 0 137126 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output91
timestamp 1712078602
transform 1 0 137448 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output92
timestamp 1712078602
transform 1 0 13018 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output93
timestamp 1712078602
transform 1 0 138920 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output94
timestamp 1712078602
transform 1 0 140438 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output95
timestamp 1712078602
transform 1 0 142278 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output96
timestamp 1712078602
transform 1 0 143566 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output97
timestamp 1712078602
transform 1 0 145038 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output98
timestamp 1712078602
transform 1 0 146602 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output99
timestamp 1712078602
transform 1 0 148120 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output100
timestamp 1712078602
transform 1 0 149638 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output101
timestamp 1712078602
transform 1 0 151294 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output102
timestamp 1712078602
transform 1 0 152214 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output103
timestamp 1712078602
transform 1 0 13892 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__clkbuf_1  output104
timestamp 1712078602
transform 1 0 690 0 -1 4352
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1712078602
transform 1 0 552 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1712078602
transform -1 0 152904 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1712078602
transform 1 0 552 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1712078602
transform -1 0 152904 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1712078602
transform 1 0 552 0 1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1712078602
transform -1 0 152904 0 1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1712078602
transform 1 0 552 0 -1 2176
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1712078602
transform -1 0 152904 0 -1 2176
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1712078602
transform 1 0 552 0 1 2176
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1712078602
transform -1 0 152904 0 1 2176
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1712078602
transform 1 0 552 0 -1 2720
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1712078602
transform -1 0 152904 0 -1 2720
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1712078602
transform 1 0 552 0 1 2720
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1712078602
transform -1 0 152904 0 1 2720
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1712078602
transform 1 0 552 0 -1 3264
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1712078602
transform -1 0 152904 0 -1 3264
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1712078602
transform 1 0 552 0 1 3264
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1712078602
transform -1 0 152904 0 1 3264
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1712078602
transform 1 0 552 0 -1 3808
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1712078602
transform -1 0 152904 0 -1 3808
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1712078602
transform 1 0 552 0 1 3808
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1712078602
transform -1 0 152904 0 1 3808
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1712078602
transform 1 0 552 0 -1 4352
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1712078602
transform -1 0 152904 0 -1 4352
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1712078602
transform 1 0 552 0 1 4352
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1712078602
transform -1 0 152904 0 1 4352
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1712078602
transform 1 0 552 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1712078602
transform -1 0 152904 0 -1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1712078602
transform 1 0 552 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1712078602
transform -1 0 152904 0 1 4896
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1712078602
transform 1 0 552 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1712078602
transform -1 0 152904 0 -1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1712078602
transform 1 0 552 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1712078602
transform -1 0 152904 0 1 5440
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1712078602
transform 1 0 552 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1712078602
transform -1 0 152904 0 -1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1712078602
transform 1 0 552 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1712078602
transform -1 0 152904 0 1 5984
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1712078602
transform 1 0 552 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1712078602
transform -1 0 152904 0 -1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1712078602
transform 1 0 552 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1712078602
transform -1 0 152904 0 1 6528
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 1840 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1712078602
transform 1 0 3128 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1712078602
transform 1 0 4416 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1712078602
transform 1 0 5704 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1712078602
transform 1 0 6992 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1712078602
transform 1 0 8280 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1712078602
transform 1 0 9568 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1712078602
transform 1 0 10856 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1712078602
transform 1 0 12144 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1712078602
transform 1 0 13432 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1712078602
transform 1 0 14720 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1712078602
transform 1 0 16008 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1712078602
transform 1 0 17296 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1712078602
transform 1 0 18584 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1712078602
transform 1 0 19872 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1712078602
transform 1 0 21160 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1712078602
transform 1 0 22448 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1712078602
transform 1 0 23736 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1712078602
transform 1 0 25024 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1712078602
transform 1 0 26312 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1712078602
transform 1 0 27600 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1712078602
transform 1 0 28888 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1712078602
transform 1 0 30176 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1712078602
transform 1 0 31464 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1712078602
transform 1 0 32752 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1712078602
transform 1 0 34040 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1712078602
transform 1 0 35328 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1712078602
transform 1 0 36616 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1712078602
transform 1 0 37904 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1712078602
transform 1 0 39192 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1712078602
transform 1 0 40480 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1712078602
transform 1 0 41768 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1712078602
transform 1 0 43056 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1712078602
transform 1 0 44344 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1712078602
transform 1 0 45632 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1712078602
transform 1 0 46920 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1712078602
transform 1 0 48208 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1712078602
transform 1 0 49496 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1712078602
transform 1 0 50784 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1712078602
transform 1 0 52072 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1712078602
transform 1 0 53360 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1712078602
transform 1 0 54648 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1712078602
transform 1 0 55936 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1712078602
transform 1 0 57224 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1712078602
transform 1 0 58512 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1712078602
transform 1 0 59800 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1712078602
transform 1 0 61088 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1712078602
transform 1 0 62376 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1712078602
transform 1 0 63664 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1712078602
transform 1 0 64952 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1712078602
transform 1 0 66240 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1712078602
transform 1 0 67528 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1712078602
transform 1 0 68816 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1712078602
transform 1 0 70104 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1712078602
transform 1 0 71392 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1712078602
transform 1 0 72680 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1712078602
transform 1 0 73968 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1712078602
transform 1 0 75256 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1712078602
transform 1 0 76544 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1712078602
transform 1 0 77832 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1712078602
transform 1 0 79120 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1712078602
transform 1 0 80408 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1712078602
transform 1 0 81696 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1712078602
transform 1 0 82984 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1712078602
transform 1 0 84272 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1712078602
transform 1 0 85560 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1712078602
transform 1 0 86848 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1712078602
transform 1 0 88136 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1712078602
transform 1 0 89424 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1712078602
transform 1 0 90712 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1712078602
transform 1 0 92000 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1712078602
transform 1 0 93288 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1712078602
transform 1 0 94576 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1712078602
transform 1 0 95864 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1712078602
transform 1 0 97152 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1712078602
transform 1 0 98440 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1712078602
transform 1 0 99728 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1712078602
transform 1 0 101016 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1712078602
transform 1 0 102304 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1712078602
transform 1 0 103592 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1712078602
transform 1 0 104880 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1712078602
transform 1 0 106168 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1712078602
transform 1 0 107456 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1712078602
transform 1 0 108744 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1712078602
transform 1 0 110032 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1712078602
transform 1 0 111320 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1712078602
transform 1 0 112608 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1712078602
transform 1 0 113896 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1712078602
transform 1 0 115184 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1712078602
transform 1 0 116472 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1712078602
transform 1 0 117760 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1712078602
transform 1 0 119048 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1712078602
transform 1 0 120336 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1712078602
transform 1 0 121624 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1712078602
transform 1 0 122912 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1712078602
transform 1 0 124200 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1712078602
transform 1 0 125488 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1712078602
transform 1 0 126776 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1712078602
transform 1 0 128064 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1712078602
transform 1 0 129352 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1712078602
transform 1 0 130640 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1712078602
transform 1 0 131928 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1712078602
transform 1 0 133216 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1712078602
transform 1 0 134504 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1712078602
transform 1 0 135792 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1712078602
transform 1 0 137080 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1712078602
transform 1 0 138368 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1712078602
transform 1 0 139656 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1712078602
transform 1 0 140944 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1712078602
transform 1 0 142232 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1712078602
transform 1 0 143520 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1712078602
transform 1 0 144808 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1712078602
transform 1 0 146096 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1712078602
transform 1 0 147384 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1712078602
transform 1 0 148672 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1712078602
transform 1 0 149960 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1712078602
transform 1 0 151248 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1712078602
transform 1 0 152536 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1712078602
transform 1 0 3128 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1712078602
transform 1 0 5704 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1712078602
transform 1 0 8280 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1712078602
transform 1 0 10856 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1712078602
transform 1 0 13432 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1712078602
transform 1 0 16008 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1712078602
transform 1 0 18584 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1712078602
transform 1 0 21160 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1712078602
transform 1 0 23736 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1712078602
transform 1 0 26312 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1712078602
transform 1 0 28888 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1712078602
transform 1 0 31464 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1712078602
transform 1 0 34040 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1712078602
transform 1 0 36616 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1712078602
transform 1 0 39192 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1712078602
transform 1 0 41768 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1712078602
transform 1 0 44344 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1712078602
transform 1 0 46920 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1712078602
transform 1 0 49496 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1712078602
transform 1 0 52072 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1712078602
transform 1 0 54648 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1712078602
transform 1 0 57224 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1712078602
transform 1 0 59800 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1712078602
transform 1 0 62376 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1712078602
transform 1 0 64952 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1712078602
transform 1 0 67528 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1712078602
transform 1 0 70104 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1712078602
transform 1 0 72680 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1712078602
transform 1 0 75256 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1712078602
transform 1 0 77832 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1712078602
transform 1 0 80408 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1712078602
transform 1 0 82984 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1712078602
transform 1 0 85560 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1712078602
transform 1 0 88136 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1712078602
transform 1 0 90712 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1712078602
transform 1 0 93288 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1712078602
transform 1 0 95864 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1712078602
transform 1 0 98440 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1712078602
transform 1 0 101016 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1712078602
transform 1 0 103592 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1712078602
transform 1 0 106168 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1712078602
transform 1 0 108744 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1712078602
transform 1 0 111320 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1712078602
transform 1 0 113896 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1712078602
transform 1 0 116472 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1712078602
transform 1 0 119048 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1712078602
transform 1 0 121624 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1712078602
transform 1 0 124200 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1712078602
transform 1 0 126776 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1712078602
transform 1 0 129352 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1712078602
transform 1 0 131928 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1712078602
transform 1 0 134504 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1712078602
transform 1 0 137080 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1712078602
transform 1 0 139656 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1712078602
transform 1 0 142232 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1712078602
transform 1 0 144808 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1712078602
transform 1 0 147384 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1712078602
transform 1 0 149960 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1712078602
transform 1 0 152536 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1712078602
transform 1 0 1840 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1712078602
transform 1 0 4416 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1712078602
transform 1 0 6992 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1712078602
transform 1 0 9568 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1712078602
transform 1 0 12144 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1712078602
transform 1 0 14720 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1712078602
transform 1 0 17296 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1712078602
transform 1 0 19872 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1712078602
transform 1 0 22448 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1712078602
transform 1 0 25024 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1712078602
transform 1 0 27600 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1712078602
transform 1 0 30176 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1712078602
transform 1 0 32752 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1712078602
transform 1 0 35328 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1712078602
transform 1 0 37904 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1712078602
transform 1 0 40480 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1712078602
transform 1 0 43056 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1712078602
transform 1 0 45632 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1712078602
transform 1 0 48208 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1712078602
transform 1 0 50784 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1712078602
transform 1 0 53360 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1712078602
transform 1 0 55936 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1712078602
transform 1 0 58512 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1712078602
transform 1 0 61088 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1712078602
transform 1 0 63664 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1712078602
transform 1 0 66240 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1712078602
transform 1 0 68816 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1712078602
transform 1 0 71392 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1712078602
transform 1 0 73968 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1712078602
transform 1 0 76544 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1712078602
transform 1 0 79120 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1712078602
transform 1 0 81696 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1712078602
transform 1 0 84272 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1712078602
transform 1 0 86848 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1712078602
transform 1 0 89424 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1712078602
transform 1 0 92000 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1712078602
transform 1 0 94576 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1712078602
transform 1 0 97152 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1712078602
transform 1 0 99728 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1712078602
transform 1 0 102304 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1712078602
transform 1 0 104880 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1712078602
transform 1 0 107456 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1712078602
transform 1 0 110032 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1712078602
transform 1 0 112608 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1712078602
transform 1 0 115184 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1712078602
transform 1 0 117760 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1712078602
transform 1 0 120336 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1712078602
transform 1 0 122912 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1712078602
transform 1 0 125488 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1712078602
transform 1 0 128064 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1712078602
transform 1 0 130640 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1712078602
transform 1 0 133216 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1712078602
transform 1 0 135792 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1712078602
transform 1 0 138368 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1712078602
transform 1 0 140944 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1712078602
transform 1 0 143520 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1712078602
transform 1 0 146096 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1712078602
transform 1 0 148672 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1712078602
transform 1 0 151248 0 1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1712078602
transform 1 0 3128 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1712078602
transform 1 0 5704 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1712078602
transform 1 0 8280 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1712078602
transform 1 0 10856 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1712078602
transform 1 0 13432 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1712078602
transform 1 0 16008 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1712078602
transform 1 0 18584 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1712078602
transform 1 0 21160 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1712078602
transform 1 0 23736 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1712078602
transform 1 0 26312 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1712078602
transform 1 0 28888 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1712078602
transform 1 0 31464 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1712078602
transform 1 0 34040 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1712078602
transform 1 0 36616 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1712078602
transform 1 0 39192 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1712078602
transform 1 0 41768 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1712078602
transform 1 0 44344 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1712078602
transform 1 0 46920 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1712078602
transform 1 0 49496 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1712078602
transform 1 0 52072 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1712078602
transform 1 0 54648 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1712078602
transform 1 0 57224 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1712078602
transform 1 0 59800 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1712078602
transform 1 0 62376 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1712078602
transform 1 0 64952 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1712078602
transform 1 0 67528 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1712078602
transform 1 0 70104 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1712078602
transform 1 0 72680 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1712078602
transform 1 0 75256 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1712078602
transform 1 0 77832 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1712078602
transform 1 0 80408 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1712078602
transform 1 0 82984 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1712078602
transform 1 0 85560 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1712078602
transform 1 0 88136 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1712078602
transform 1 0 90712 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1712078602
transform 1 0 93288 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1712078602
transform 1 0 95864 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1712078602
transform 1 0 98440 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1712078602
transform 1 0 101016 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1712078602
transform 1 0 103592 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1712078602
transform 1 0 106168 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1712078602
transform 1 0 108744 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1712078602
transform 1 0 111320 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1712078602
transform 1 0 113896 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1712078602
transform 1 0 116472 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1712078602
transform 1 0 119048 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1712078602
transform 1 0 121624 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1712078602
transform 1 0 124200 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1712078602
transform 1 0 126776 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1712078602
transform 1 0 129352 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1712078602
transform 1 0 131928 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1712078602
transform 1 0 134504 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1712078602
transform 1 0 137080 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1712078602
transform 1 0 139656 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1712078602
transform 1 0 142232 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1712078602
transform 1 0 144808 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1712078602
transform 1 0 147384 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1712078602
transform 1 0 149960 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1712078602
transform 1 0 152536 0 -1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1712078602
transform 1 0 1840 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1712078602
transform 1 0 4416 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1712078602
transform 1 0 6992 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1712078602
transform 1 0 9568 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1712078602
transform 1 0 12144 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1712078602
transform 1 0 14720 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1712078602
transform 1 0 17296 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1712078602
transform 1 0 19872 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1712078602
transform 1 0 22448 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1712078602
transform 1 0 25024 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1712078602
transform 1 0 27600 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1712078602
transform 1 0 30176 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1712078602
transform 1 0 32752 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1712078602
transform 1 0 35328 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1712078602
transform 1 0 37904 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1712078602
transform 1 0 40480 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1712078602
transform 1 0 43056 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1712078602
transform 1 0 45632 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1712078602
transform 1 0 48208 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1712078602
transform 1 0 50784 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1712078602
transform 1 0 53360 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1712078602
transform 1 0 55936 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1712078602
transform 1 0 58512 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1712078602
transform 1 0 61088 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1712078602
transform 1 0 63664 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1712078602
transform 1 0 66240 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1712078602
transform 1 0 68816 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1712078602
transform 1 0 71392 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1712078602
transform 1 0 73968 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1712078602
transform 1 0 76544 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1712078602
transform 1 0 79120 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1712078602
transform 1 0 81696 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1712078602
transform 1 0 84272 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1712078602
transform 1 0 86848 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1712078602
transform 1 0 89424 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1712078602
transform 1 0 92000 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1712078602
transform 1 0 94576 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1712078602
transform 1 0 97152 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1712078602
transform 1 0 99728 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1712078602
transform 1 0 102304 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1712078602
transform 1 0 104880 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1712078602
transform 1 0 107456 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1712078602
transform 1 0 110032 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1712078602
transform 1 0 112608 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1712078602
transform 1 0 115184 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1712078602
transform 1 0 117760 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1712078602
transform 1 0 120336 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1712078602
transform 1 0 122912 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1712078602
transform 1 0 125488 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1712078602
transform 1 0 128064 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1712078602
transform 1 0 130640 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1712078602
transform 1 0 133216 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1712078602
transform 1 0 135792 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1712078602
transform 1 0 138368 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1712078602
transform 1 0 140944 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1712078602
transform 1 0 143520 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1712078602
transform 1 0 146096 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1712078602
transform 1 0 148672 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1712078602
transform 1 0 151248 0 1 2176
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1712078602
transform 1 0 3128 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1712078602
transform 1 0 5704 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1712078602
transform 1 0 8280 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1712078602
transform 1 0 10856 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1712078602
transform 1 0 13432 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1712078602
transform 1 0 16008 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1712078602
transform 1 0 18584 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1712078602
transform 1 0 21160 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1712078602
transform 1 0 23736 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1712078602
transform 1 0 26312 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1712078602
transform 1 0 28888 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1712078602
transform 1 0 31464 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1712078602
transform 1 0 34040 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1712078602
transform 1 0 36616 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1712078602
transform 1 0 39192 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1712078602
transform 1 0 41768 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1712078602
transform 1 0 44344 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1712078602
transform 1 0 46920 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1712078602
transform 1 0 49496 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1712078602
transform 1 0 52072 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1712078602
transform 1 0 54648 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1712078602
transform 1 0 57224 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1712078602
transform 1 0 59800 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1712078602
transform 1 0 62376 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1712078602
transform 1 0 64952 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1712078602
transform 1 0 67528 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1712078602
transform 1 0 70104 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1712078602
transform 1 0 72680 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1712078602
transform 1 0 75256 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1712078602
transform 1 0 77832 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1712078602
transform 1 0 80408 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1712078602
transform 1 0 82984 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1712078602
transform 1 0 85560 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1712078602
transform 1 0 88136 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1712078602
transform 1 0 90712 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1712078602
transform 1 0 93288 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1712078602
transform 1 0 95864 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1712078602
transform 1 0 98440 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1712078602
transform 1 0 101016 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1712078602
transform 1 0 103592 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1712078602
transform 1 0 106168 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1712078602
transform 1 0 108744 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1712078602
transform 1 0 111320 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1712078602
transform 1 0 113896 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1712078602
transform 1 0 116472 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1712078602
transform 1 0 119048 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1712078602
transform 1 0 121624 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1712078602
transform 1 0 124200 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1712078602
transform 1 0 126776 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1712078602
transform 1 0 129352 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1712078602
transform 1 0 131928 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1712078602
transform 1 0 134504 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1712078602
transform 1 0 137080 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1712078602
transform 1 0 139656 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1712078602
transform 1 0 142232 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1712078602
transform 1 0 144808 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1712078602
transform 1 0 147384 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1712078602
transform 1 0 149960 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1712078602
transform 1 0 152536 0 -1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1712078602
transform 1 0 1840 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1712078602
transform 1 0 4416 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1712078602
transform 1 0 6992 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1712078602
transform 1 0 9568 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1712078602
transform 1 0 12144 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1712078602
transform 1 0 14720 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1712078602
transform 1 0 17296 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1712078602
transform 1 0 19872 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1712078602
transform 1 0 22448 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1712078602
transform 1 0 25024 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1712078602
transform 1 0 27600 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1712078602
transform 1 0 30176 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1712078602
transform 1 0 32752 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1712078602
transform 1 0 35328 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1712078602
transform 1 0 37904 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1712078602
transform 1 0 40480 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1712078602
transform 1 0 43056 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1712078602
transform 1 0 45632 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1712078602
transform 1 0 48208 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1712078602
transform 1 0 50784 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1712078602
transform 1 0 53360 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1712078602
transform 1 0 55936 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1712078602
transform 1 0 58512 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1712078602
transform 1 0 61088 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1712078602
transform 1 0 63664 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1712078602
transform 1 0 66240 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1712078602
transform 1 0 68816 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1712078602
transform 1 0 71392 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1712078602
transform 1 0 73968 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1712078602
transform 1 0 76544 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1712078602
transform 1 0 79120 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1712078602
transform 1 0 81696 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1712078602
transform 1 0 84272 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1712078602
transform 1 0 86848 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1712078602
transform 1 0 89424 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1712078602
transform 1 0 92000 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1712078602
transform 1 0 94576 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1712078602
transform 1 0 97152 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1712078602
transform 1 0 99728 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1712078602
transform 1 0 102304 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1712078602
transform 1 0 104880 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1712078602
transform 1 0 107456 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1712078602
transform 1 0 110032 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1712078602
transform 1 0 112608 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1712078602
transform 1 0 115184 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1712078602
transform 1 0 117760 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1712078602
transform 1 0 120336 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1712078602
transform 1 0 122912 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1712078602
transform 1 0 125488 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1712078602
transform 1 0 128064 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1712078602
transform 1 0 130640 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1712078602
transform 1 0 133216 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1712078602
transform 1 0 135792 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1712078602
transform 1 0 138368 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1712078602
transform 1 0 140944 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1712078602
transform 1 0 143520 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1712078602
transform 1 0 146096 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1712078602
transform 1 0 148672 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1712078602
transform 1 0 151248 0 1 2720
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1712078602
transform 1 0 3128 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1712078602
transform 1 0 5704 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1712078602
transform 1 0 8280 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1712078602
transform 1 0 10856 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1712078602
transform 1 0 13432 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1712078602
transform 1 0 16008 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1712078602
transform 1 0 18584 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1712078602
transform 1 0 21160 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1712078602
transform 1 0 23736 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1712078602
transform 1 0 26312 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1712078602
transform 1 0 28888 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1712078602
transform 1 0 31464 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1712078602
transform 1 0 34040 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1712078602
transform 1 0 36616 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1712078602
transform 1 0 39192 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1712078602
transform 1 0 41768 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1712078602
transform 1 0 44344 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1712078602
transform 1 0 46920 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1712078602
transform 1 0 49496 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1712078602
transform 1 0 52072 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1712078602
transform 1 0 54648 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1712078602
transform 1 0 57224 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1712078602
transform 1 0 59800 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1712078602
transform 1 0 62376 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1712078602
transform 1 0 64952 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1712078602
transform 1 0 67528 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1712078602
transform 1 0 70104 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1712078602
transform 1 0 72680 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1712078602
transform 1 0 75256 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1712078602
transform 1 0 77832 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1712078602
transform 1 0 80408 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1712078602
transform 1 0 82984 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1712078602
transform 1 0 85560 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1712078602
transform 1 0 88136 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1712078602
transform 1 0 90712 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1712078602
transform 1 0 93288 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1712078602
transform 1 0 95864 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1712078602
transform 1 0 98440 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1712078602
transform 1 0 101016 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1712078602
transform 1 0 103592 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1712078602
transform 1 0 106168 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1712078602
transform 1 0 108744 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1712078602
transform 1 0 111320 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1712078602
transform 1 0 113896 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1712078602
transform 1 0 116472 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1712078602
transform 1 0 119048 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1712078602
transform 1 0 121624 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1712078602
transform 1 0 124200 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1712078602
transform 1 0 126776 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1712078602
transform 1 0 129352 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1712078602
transform 1 0 131928 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1712078602
transform 1 0 134504 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1712078602
transform 1 0 137080 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1712078602
transform 1 0 139656 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1712078602
transform 1 0 142232 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1712078602
transform 1 0 144808 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1712078602
transform 1 0 147384 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1712078602
transform 1 0 149960 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1712078602
transform 1 0 152536 0 -1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1712078602
transform 1 0 1840 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1712078602
transform 1 0 4416 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1712078602
transform 1 0 6992 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1712078602
transform 1 0 9568 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1712078602
transform 1 0 12144 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1712078602
transform 1 0 14720 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1712078602
transform 1 0 17296 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1712078602
transform 1 0 19872 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1712078602
transform 1 0 22448 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1712078602
transform 1 0 25024 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1712078602
transform 1 0 27600 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1712078602
transform 1 0 30176 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1712078602
transform 1 0 32752 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1712078602
transform 1 0 35328 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1712078602
transform 1 0 37904 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1712078602
transform 1 0 40480 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1712078602
transform 1 0 43056 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1712078602
transform 1 0 45632 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1712078602
transform 1 0 48208 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1712078602
transform 1 0 50784 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1712078602
transform 1 0 53360 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1712078602
transform 1 0 55936 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1712078602
transform 1 0 58512 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1712078602
transform 1 0 61088 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1712078602
transform 1 0 63664 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1712078602
transform 1 0 66240 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1712078602
transform 1 0 68816 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1712078602
transform 1 0 71392 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1712078602
transform 1 0 73968 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1712078602
transform 1 0 76544 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1712078602
transform 1 0 79120 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1712078602
transform 1 0 81696 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1712078602
transform 1 0 84272 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1712078602
transform 1 0 86848 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1712078602
transform 1 0 89424 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1712078602
transform 1 0 92000 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1712078602
transform 1 0 94576 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1712078602
transform 1 0 97152 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1712078602
transform 1 0 99728 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1712078602
transform 1 0 102304 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1712078602
transform 1 0 104880 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1712078602
transform 1 0 107456 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1712078602
transform 1 0 110032 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1712078602
transform 1 0 112608 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1712078602
transform 1 0 115184 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1712078602
transform 1 0 117760 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1712078602
transform 1 0 120336 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1712078602
transform 1 0 122912 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1712078602
transform 1 0 125488 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1712078602
transform 1 0 128064 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1712078602
transform 1 0 130640 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1712078602
transform 1 0 133216 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1712078602
transform 1 0 135792 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1712078602
transform 1 0 138368 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1712078602
transform 1 0 140944 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1712078602
transform 1 0 143520 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1712078602
transform 1 0 146096 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1712078602
transform 1 0 148672 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1712078602
transform 1 0 151248 0 1 3264
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1712078602
transform 1 0 3128 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1712078602
transform 1 0 5704 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1712078602
transform 1 0 8280 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1712078602
transform 1 0 10856 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1712078602
transform 1 0 13432 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1712078602
transform 1 0 16008 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1712078602
transform 1 0 18584 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1712078602
transform 1 0 21160 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1712078602
transform 1 0 23736 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1712078602
transform 1 0 26312 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1712078602
transform 1 0 28888 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1712078602
transform 1 0 31464 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1712078602
transform 1 0 34040 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1712078602
transform 1 0 36616 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1712078602
transform 1 0 39192 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1712078602
transform 1 0 41768 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1712078602
transform 1 0 44344 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1712078602
transform 1 0 46920 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1712078602
transform 1 0 49496 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1712078602
transform 1 0 52072 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1712078602
transform 1 0 54648 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1712078602
transform 1 0 57224 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1712078602
transform 1 0 59800 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1712078602
transform 1 0 62376 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1712078602
transform 1 0 64952 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1712078602
transform 1 0 67528 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1712078602
transform 1 0 70104 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1712078602
transform 1 0 72680 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1712078602
transform 1 0 75256 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1712078602
transform 1 0 77832 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1712078602
transform 1 0 80408 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1712078602
transform 1 0 82984 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1712078602
transform 1 0 85560 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1712078602
transform 1 0 88136 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1712078602
transform 1 0 90712 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1712078602
transform 1 0 93288 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1712078602
transform 1 0 95864 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1712078602
transform 1 0 98440 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1712078602
transform 1 0 101016 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1712078602
transform 1 0 103592 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1712078602
transform 1 0 106168 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1712078602
transform 1 0 108744 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1712078602
transform 1 0 111320 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1712078602
transform 1 0 113896 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1712078602
transform 1 0 116472 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1712078602
transform 1 0 119048 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1712078602
transform 1 0 121624 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1712078602
transform 1 0 124200 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1712078602
transform 1 0 126776 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1712078602
transform 1 0 129352 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1712078602
transform 1 0 131928 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1712078602
transform 1 0 134504 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1712078602
transform 1 0 137080 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1712078602
transform 1 0 139656 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1712078602
transform 1 0 142232 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1712078602
transform 1 0 144808 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1712078602
transform 1 0 147384 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1712078602
transform 1 0 149960 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1712078602
transform 1 0 152536 0 -1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1712078602
transform 1 0 1840 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1712078602
transform 1 0 4416 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1712078602
transform 1 0 6992 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1712078602
transform 1 0 9568 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1712078602
transform 1 0 12144 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1712078602
transform 1 0 14720 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1712078602
transform 1 0 17296 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1712078602
transform 1 0 19872 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1712078602
transform 1 0 22448 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1712078602
transform 1 0 25024 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1712078602
transform 1 0 27600 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1712078602
transform 1 0 30176 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1712078602
transform 1 0 32752 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1712078602
transform 1 0 35328 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1712078602
transform 1 0 37904 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1712078602
transform 1 0 40480 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1712078602
transform 1 0 43056 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1712078602
transform 1 0 45632 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1712078602
transform 1 0 48208 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1712078602
transform 1 0 50784 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1712078602
transform 1 0 53360 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1712078602
transform 1 0 55936 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1712078602
transform 1 0 58512 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1712078602
transform 1 0 61088 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1712078602
transform 1 0 63664 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1712078602
transform 1 0 66240 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1712078602
transform 1 0 68816 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1712078602
transform 1 0 71392 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1712078602
transform 1 0 73968 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1712078602
transform 1 0 76544 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1712078602
transform 1 0 79120 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1712078602
transform 1 0 81696 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1712078602
transform 1 0 84272 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1712078602
transform 1 0 86848 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1712078602
transform 1 0 89424 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1712078602
transform 1 0 92000 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1712078602
transform 1 0 94576 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1712078602
transform 1 0 97152 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1712078602
transform 1 0 99728 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1712078602
transform 1 0 102304 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1712078602
transform 1 0 104880 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1712078602
transform 1 0 107456 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1712078602
transform 1 0 110032 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1712078602
transform 1 0 112608 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1712078602
transform 1 0 115184 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1712078602
transform 1 0 117760 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1712078602
transform 1 0 120336 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1712078602
transform 1 0 122912 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1712078602
transform 1 0 125488 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1712078602
transform 1 0 128064 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1712078602
transform 1 0 130640 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1712078602
transform 1 0 133216 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1712078602
transform 1 0 135792 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1712078602
transform 1 0 138368 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1712078602
transform 1 0 140944 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1712078602
transform 1 0 143520 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1712078602
transform 1 0 146096 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1712078602
transform 1 0 148672 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1712078602
transform 1 0 151248 0 1 3808
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1712078602
transform 1 0 3128 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1712078602
transform 1 0 5704 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1712078602
transform 1 0 8280 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1712078602
transform 1 0 10856 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1712078602
transform 1 0 13432 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1712078602
transform 1 0 16008 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1712078602
transform 1 0 18584 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1712078602
transform 1 0 21160 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1712078602
transform 1 0 23736 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1712078602
transform 1 0 26312 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1712078602
transform 1 0 28888 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1712078602
transform 1 0 31464 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1712078602
transform 1 0 34040 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1712078602
transform 1 0 36616 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1712078602
transform 1 0 39192 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1712078602
transform 1 0 41768 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1712078602
transform 1 0 44344 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1712078602
transform 1 0 46920 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1712078602
transform 1 0 49496 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1712078602
transform 1 0 52072 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1712078602
transform 1 0 54648 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1712078602
transform 1 0 57224 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1712078602
transform 1 0 59800 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1712078602
transform 1 0 62376 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1712078602
transform 1 0 64952 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1712078602
transform 1 0 67528 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1712078602
transform 1 0 70104 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1712078602
transform 1 0 72680 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1712078602
transform 1 0 75256 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1712078602
transform 1 0 77832 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1712078602
transform 1 0 80408 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1712078602
transform 1 0 82984 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1712078602
transform 1 0 85560 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1712078602
transform 1 0 88136 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1712078602
transform 1 0 90712 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1712078602
transform 1 0 93288 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1712078602
transform 1 0 95864 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1712078602
transform 1 0 98440 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1712078602
transform 1 0 101016 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1712078602
transform 1 0 103592 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1712078602
transform 1 0 106168 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1712078602
transform 1 0 108744 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1712078602
transform 1 0 111320 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1712078602
transform 1 0 113896 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1712078602
transform 1 0 116472 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1712078602
transform 1 0 119048 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1712078602
transform 1 0 121624 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1712078602
transform 1 0 124200 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1712078602
transform 1 0 126776 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1712078602
transform 1 0 129352 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1712078602
transform 1 0 131928 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1712078602
transform 1 0 134504 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1712078602
transform 1 0 137080 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1712078602
transform 1 0 139656 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1712078602
transform 1 0 142232 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1712078602
transform 1 0 144808 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1712078602
transform 1 0 147384 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1712078602
transform 1 0 149960 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1712078602
transform 1 0 152536 0 -1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1712078602
transform 1 0 1840 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1712078602
transform 1 0 4416 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1712078602
transform 1 0 6992 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1712078602
transform 1 0 9568 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1712078602
transform 1 0 12144 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1712078602
transform 1 0 14720 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1712078602
transform 1 0 17296 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1712078602
transform 1 0 19872 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1712078602
transform 1 0 22448 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1712078602
transform 1 0 25024 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1712078602
transform 1 0 27600 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1712078602
transform 1 0 30176 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1712078602
transform 1 0 32752 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1712078602
transform 1 0 35328 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1712078602
transform 1 0 37904 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1712078602
transform 1 0 40480 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1712078602
transform 1 0 43056 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1712078602
transform 1 0 45632 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1712078602
transform 1 0 48208 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1712078602
transform 1 0 50784 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1712078602
transform 1 0 53360 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1712078602
transform 1 0 55936 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1712078602
transform 1 0 58512 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1712078602
transform 1 0 61088 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1712078602
transform 1 0 63664 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1712078602
transform 1 0 66240 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1712078602
transform 1 0 68816 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1712078602
transform 1 0 71392 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1712078602
transform 1 0 73968 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1712078602
transform 1 0 76544 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1712078602
transform 1 0 79120 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1712078602
transform 1 0 81696 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1712078602
transform 1 0 84272 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1712078602
transform 1 0 86848 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1712078602
transform 1 0 89424 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1712078602
transform 1 0 92000 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1712078602
transform 1 0 94576 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1712078602
transform 1 0 97152 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1712078602
transform 1 0 99728 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1712078602
transform 1 0 102304 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1712078602
transform 1 0 104880 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1712078602
transform 1 0 107456 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1712078602
transform 1 0 110032 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1712078602
transform 1 0 112608 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1712078602
transform 1 0 115184 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1712078602
transform 1 0 117760 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1712078602
transform 1 0 120336 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1712078602
transform 1 0 122912 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1712078602
transform 1 0 125488 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1712078602
transform 1 0 128064 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1712078602
transform 1 0 130640 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1712078602
transform 1 0 133216 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1712078602
transform 1 0 135792 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1712078602
transform 1 0 138368 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1712078602
transform 1 0 140944 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1712078602
transform 1 0 143520 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1712078602
transform 1 0 146096 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1712078602
transform 1 0 148672 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1712078602
transform 1 0 151248 0 1 4352
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1712078602
transform 1 0 3128 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1712078602
transform 1 0 5704 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1712078602
transform 1 0 8280 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1712078602
transform 1 0 10856 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1712078602
transform 1 0 13432 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1712078602
transform 1 0 16008 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1712078602
transform 1 0 18584 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1712078602
transform 1 0 21160 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1712078602
transform 1 0 23736 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1712078602
transform 1 0 26312 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1712078602
transform 1 0 28888 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1712078602
transform 1 0 31464 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1712078602
transform 1 0 34040 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1712078602
transform 1 0 36616 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1712078602
transform 1 0 39192 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1712078602
transform 1 0 41768 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1712078602
transform 1 0 44344 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1712078602
transform 1 0 46920 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1712078602
transform 1 0 49496 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1712078602
transform 1 0 52072 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1712078602
transform 1 0 54648 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1712078602
transform 1 0 57224 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1712078602
transform 1 0 59800 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1712078602
transform 1 0 62376 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1712078602
transform 1 0 64952 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1712078602
transform 1 0 67528 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1712078602
transform 1 0 70104 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1712078602
transform 1 0 72680 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1712078602
transform 1 0 75256 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1712078602
transform 1 0 77832 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1712078602
transform 1 0 80408 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1712078602
transform 1 0 82984 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1712078602
transform 1 0 85560 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1712078602
transform 1 0 88136 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1712078602
transform 1 0 90712 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1712078602
transform 1 0 93288 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1712078602
transform 1 0 95864 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1712078602
transform 1 0 98440 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1712078602
transform 1 0 101016 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1712078602
transform 1 0 103592 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1712078602
transform 1 0 106168 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1712078602
transform 1 0 108744 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1712078602
transform 1 0 111320 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1712078602
transform 1 0 113896 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1712078602
transform 1 0 116472 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1712078602
transform 1 0 119048 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1712078602
transform 1 0 121624 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1712078602
transform 1 0 124200 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1712078602
transform 1 0 126776 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1712078602
transform 1 0 129352 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1712078602
transform 1 0 131928 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1712078602
transform 1 0 134504 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1712078602
transform 1 0 137080 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1712078602
transform 1 0 139656 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1712078602
transform 1 0 142232 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1712078602
transform 1 0 144808 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1712078602
transform 1 0 147384 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1712078602
transform 1 0 149960 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1712078602
transform 1 0 152536 0 -1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1712078602
transform 1 0 1840 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1712078602
transform 1 0 4416 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1712078602
transform 1 0 6992 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1712078602
transform 1 0 9568 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1712078602
transform 1 0 12144 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1712078602
transform 1 0 14720 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1712078602
transform 1 0 17296 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1712078602
transform 1 0 19872 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1712078602
transform 1 0 22448 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1712078602
transform 1 0 25024 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1712078602
transform 1 0 27600 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1712078602
transform 1 0 30176 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1712078602
transform 1 0 32752 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1712078602
transform 1 0 35328 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1712078602
transform 1 0 37904 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1712078602
transform 1 0 40480 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1712078602
transform 1 0 43056 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1712078602
transform 1 0 45632 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1712078602
transform 1 0 48208 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1712078602
transform 1 0 50784 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1712078602
transform 1 0 53360 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1712078602
transform 1 0 55936 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1712078602
transform 1 0 58512 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1712078602
transform 1 0 61088 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1712078602
transform 1 0 63664 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1712078602
transform 1 0 66240 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1712078602
transform 1 0 68816 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1712078602
transform 1 0 71392 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1712078602
transform 1 0 73968 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1712078602
transform 1 0 76544 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1712078602
transform 1 0 79120 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1712078602
transform 1 0 81696 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1712078602
transform 1 0 84272 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1712078602
transform 1 0 86848 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1712078602
transform 1 0 89424 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1712078602
transform 1 0 92000 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1712078602
transform 1 0 94576 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1712078602
transform 1 0 97152 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1712078602
transform 1 0 99728 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1712078602
transform 1 0 102304 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1712078602
transform 1 0 104880 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1712078602
transform 1 0 107456 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1712078602
transform 1 0 110032 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1712078602
transform 1 0 112608 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1712078602
transform 1 0 115184 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1712078602
transform 1 0 117760 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1712078602
transform 1 0 120336 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1712078602
transform 1 0 122912 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1712078602
transform 1 0 125488 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1712078602
transform 1 0 128064 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1712078602
transform 1 0 130640 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1712078602
transform 1 0 133216 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1712078602
transform 1 0 135792 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1712078602
transform 1 0 138368 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1712078602
transform 1 0 140944 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1712078602
transform 1 0 143520 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1712078602
transform 1 0 146096 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1712078602
transform 1 0 148672 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1712078602
transform 1 0 151248 0 1 4896
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1712078602
transform 1 0 3128 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1712078602
transform 1 0 5704 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1712078602
transform 1 0 8280 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1712078602
transform 1 0 10856 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1712078602
transform 1 0 13432 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1712078602
transform 1 0 16008 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1712078602
transform 1 0 18584 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1712078602
transform 1 0 21160 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1712078602
transform 1 0 23736 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1712078602
transform 1 0 26312 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1712078602
transform 1 0 28888 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1712078602
transform 1 0 31464 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1712078602
transform 1 0 34040 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1712078602
transform 1 0 36616 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1712078602
transform 1 0 39192 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1712078602
transform 1 0 41768 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1712078602
transform 1 0 44344 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1712078602
transform 1 0 46920 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1712078602
transform 1 0 49496 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1712078602
transform 1 0 52072 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1712078602
transform 1 0 54648 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1712078602
transform 1 0 57224 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1712078602
transform 1 0 59800 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1712078602
transform 1 0 62376 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1712078602
transform 1 0 64952 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1712078602
transform 1 0 67528 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1712078602
transform 1 0 70104 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1712078602
transform 1 0 72680 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1712078602
transform 1 0 75256 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1712078602
transform 1 0 77832 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1712078602
transform 1 0 80408 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1712078602
transform 1 0 82984 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1712078602
transform 1 0 85560 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1712078602
transform 1 0 88136 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1712078602
transform 1 0 90712 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1712078602
transform 1 0 93288 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1712078602
transform 1 0 95864 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1712078602
transform 1 0 98440 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1712078602
transform 1 0 101016 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1712078602
transform 1 0 103592 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1712078602
transform 1 0 106168 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1712078602
transform 1 0 108744 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1712078602
transform 1 0 111320 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1712078602
transform 1 0 113896 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1712078602
transform 1 0 116472 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1712078602
transform 1 0 119048 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1712078602
transform 1 0 121624 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1712078602
transform 1 0 124200 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1712078602
transform 1 0 126776 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1712078602
transform 1 0 129352 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1712078602
transform 1 0 131928 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1712078602
transform 1 0 134504 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1712078602
transform 1 0 137080 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1712078602
transform 1 0 139656 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1712078602
transform 1 0 142232 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1712078602
transform 1 0 144808 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1712078602
transform 1 0 147384 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1712078602
transform 1 0 149960 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1712078602
transform 1 0 152536 0 -1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1712078602
transform 1 0 1840 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1712078602
transform 1 0 4416 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1712078602
transform 1 0 6992 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1712078602
transform 1 0 9568 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1712078602
transform 1 0 12144 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1712078602
transform 1 0 14720 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1712078602
transform 1 0 17296 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1712078602
transform 1 0 19872 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1712078602
transform 1 0 22448 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1712078602
transform 1 0 25024 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1712078602
transform 1 0 27600 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1712078602
transform 1 0 30176 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1712078602
transform 1 0 32752 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1712078602
transform 1 0 35328 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1712078602
transform 1 0 37904 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1712078602
transform 1 0 40480 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1712078602
transform 1 0 43056 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1712078602
transform 1 0 45632 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1712078602
transform 1 0 48208 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1712078602
transform 1 0 50784 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1712078602
transform 1 0 53360 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1712078602
transform 1 0 55936 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1712078602
transform 1 0 58512 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1712078602
transform 1 0 61088 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1712078602
transform 1 0 63664 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1712078602
transform 1 0 66240 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1712078602
transform 1 0 68816 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1712078602
transform 1 0 71392 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1712078602
transform 1 0 73968 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1712078602
transform 1 0 76544 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1712078602
transform 1 0 79120 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1712078602
transform 1 0 81696 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1712078602
transform 1 0 84272 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1712078602
transform 1 0 86848 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1712078602
transform 1 0 89424 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1712078602
transform 1 0 92000 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1712078602
transform 1 0 94576 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1712078602
transform 1 0 97152 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1712078602
transform 1 0 99728 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1712078602
transform 1 0 102304 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1712078602
transform 1 0 104880 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1712078602
transform 1 0 107456 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1712078602
transform 1 0 110032 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1712078602
transform 1 0 112608 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1712078602
transform 1 0 115184 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1712078602
transform 1 0 117760 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1712078602
transform 1 0 120336 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1712078602
transform 1 0 122912 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1712078602
transform 1 0 125488 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1712078602
transform 1 0 128064 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1712078602
transform 1 0 130640 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1712078602
transform 1 0 133216 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1712078602
transform 1 0 135792 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1712078602
transform 1 0 138368 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1712078602
transform 1 0 140944 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1712078602
transform 1 0 143520 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1712078602
transform 1 0 146096 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1712078602
transform 1 0 148672 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1712078602
transform 1 0 151248 0 1 5440
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1712078602
transform 1 0 3128 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1712078602
transform 1 0 5704 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1712078602
transform 1 0 8280 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1712078602
transform 1 0 10856 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1712078602
transform 1 0 13432 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1712078602
transform 1 0 16008 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1712078602
transform 1 0 18584 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1712078602
transform 1 0 21160 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1712078602
transform 1 0 23736 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1712078602
transform 1 0 26312 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1712078602
transform 1 0 28888 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1712078602
transform 1 0 31464 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1712078602
transform 1 0 34040 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1712078602
transform 1 0 36616 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1712078602
transform 1 0 39192 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1712078602
transform 1 0 41768 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1712078602
transform 1 0 44344 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1712078602
transform 1 0 46920 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1712078602
transform 1 0 49496 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1712078602
transform 1 0 52072 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1712078602
transform 1 0 54648 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1712078602
transform 1 0 57224 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1712078602
transform 1 0 59800 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1712078602
transform 1 0 62376 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1712078602
transform 1 0 64952 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1712078602
transform 1 0 67528 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1712078602
transform 1 0 70104 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1712078602
transform 1 0 72680 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1712078602
transform 1 0 75256 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1712078602
transform 1 0 77832 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1712078602
transform 1 0 80408 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1712078602
transform 1 0 82984 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1712078602
transform 1 0 85560 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1712078602
transform 1 0 88136 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1712078602
transform 1 0 90712 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1712078602
transform 1 0 93288 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1712078602
transform 1 0 95864 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1712078602
transform 1 0 98440 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1712078602
transform 1 0 101016 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1712078602
transform 1 0 103592 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1712078602
transform 1 0 106168 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1712078602
transform 1 0 108744 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1712078602
transform 1 0 111320 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1712078602
transform 1 0 113896 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1712078602
transform 1 0 116472 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1712078602
transform 1 0 119048 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1712078602
transform 1 0 121624 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1712078602
transform 1 0 124200 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1712078602
transform 1 0 126776 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1712078602
transform 1 0 129352 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1712078602
transform 1 0 131928 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1712078602
transform 1 0 134504 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1712078602
transform 1 0 137080 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1712078602
transform 1 0 139656 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1712078602
transform 1 0 142232 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1712078602
transform 1 0 144808 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1712078602
transform 1 0 147384 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1712078602
transform 1 0 149960 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1712078602
transform 1 0 152536 0 -1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1712078602
transform 1 0 1840 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1712078602
transform 1 0 4416 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1712078602
transform 1 0 6992 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1712078602
transform 1 0 9568 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1712078602
transform 1 0 12144 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1712078602
transform 1 0 14720 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1712078602
transform 1 0 17296 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1712078602
transform 1 0 19872 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1712078602
transform 1 0 22448 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1712078602
transform 1 0 25024 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1712078602
transform 1 0 27600 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1712078602
transform 1 0 30176 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1712078602
transform 1 0 32752 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1712078602
transform 1 0 35328 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1712078602
transform 1 0 37904 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1712078602
transform 1 0 40480 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1712078602
transform 1 0 43056 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1712078602
transform 1 0 45632 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1712078602
transform 1 0 48208 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1712078602
transform 1 0 50784 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1712078602
transform 1 0 53360 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1712078602
transform 1 0 55936 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1712078602
transform 1 0 58512 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1712078602
transform 1 0 61088 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1712078602
transform 1 0 63664 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1712078602
transform 1 0 66240 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1712078602
transform 1 0 68816 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1712078602
transform 1 0 71392 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1712078602
transform 1 0 73968 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1712078602
transform 1 0 76544 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1712078602
transform 1 0 79120 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1712078602
transform 1 0 81696 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1712078602
transform 1 0 84272 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1712078602
transform 1 0 86848 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1712078602
transform 1 0 89424 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1712078602
transform 1 0 92000 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1712078602
transform 1 0 94576 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1712078602
transform 1 0 97152 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1712078602
transform 1 0 99728 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1712078602
transform 1 0 102304 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1712078602
transform 1 0 104880 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1712078602
transform 1 0 107456 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1712078602
transform 1 0 110032 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1712078602
transform 1 0 112608 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1712078602
transform 1 0 115184 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1712078602
transform 1 0 117760 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1712078602
transform 1 0 120336 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1712078602
transform 1 0 122912 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1712078602
transform 1 0 125488 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1712078602
transform 1 0 128064 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1712078602
transform 1 0 130640 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1712078602
transform 1 0 133216 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1712078602
transform 1 0 135792 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1712078602
transform 1 0 138368 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1712078602
transform 1 0 140944 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1712078602
transform 1 0 143520 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1712078602
transform 1 0 146096 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1712078602
transform 1 0 148672 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1712078602
transform 1 0 151248 0 1 5984
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1712078602
transform 1 0 3128 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1712078602
transform 1 0 5704 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1712078602
transform 1 0 8280 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1712078602
transform 1 0 10856 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1712078602
transform 1 0 13432 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1712078602
transform 1 0 16008 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1712078602
transform 1 0 18584 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1712078602
transform 1 0 21160 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1712078602
transform 1 0 23736 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1712078602
transform 1 0 26312 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1712078602
transform 1 0 28888 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1712078602
transform 1 0 31464 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1712078602
transform 1 0 34040 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1712078602
transform 1 0 36616 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1712078602
transform 1 0 39192 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1712078602
transform 1 0 41768 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1712078602
transform 1 0 44344 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1712078602
transform 1 0 46920 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1712078602
transform 1 0 49496 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1712078602
transform 1 0 52072 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1712078602
transform 1 0 54648 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1712078602
transform 1 0 57224 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1712078602
transform 1 0 59800 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1712078602
transform 1 0 62376 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1712078602
transform 1 0 64952 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1712078602
transform 1 0 67528 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1712078602
transform 1 0 70104 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1712078602
transform 1 0 72680 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1712078602
transform 1 0 75256 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1712078602
transform 1 0 77832 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1712078602
transform 1 0 80408 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1712078602
transform 1 0 82984 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1712078602
transform 1 0 85560 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1712078602
transform 1 0 88136 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1712078602
transform 1 0 90712 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1712078602
transform 1 0 93288 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1712078602
transform 1 0 95864 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1712078602
transform 1 0 98440 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1712078602
transform 1 0 101016 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1712078602
transform 1 0 103592 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1712078602
transform 1 0 106168 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1712078602
transform 1 0 108744 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1712078602
transform 1 0 111320 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1712078602
transform 1 0 113896 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1712078602
transform 1 0 116472 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1712078602
transform 1 0 119048 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1712078602
transform 1 0 121624 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1712078602
transform 1 0 124200 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1712078602
transform 1 0 126776 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1712078602
transform 1 0 129352 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1712078602
transform 1 0 131928 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1712078602
transform 1 0 134504 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1712078602
transform 1 0 137080 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1712078602
transform 1 0 139656 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1712078602
transform 1 0 142232 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1712078602
transform 1 0 144808 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1712078602
transform 1 0 147384 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1712078602
transform 1 0 149960 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1712078602
transform 1 0 152536 0 -1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1712078602
transform 1 0 1840 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1712078602
transform 1 0 3128 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1712078602
transform 1 0 4416 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1712078602
transform 1 0 5704 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1712078602
transform 1 0 6992 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1712078602
transform 1 0 8280 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1712078602
transform 1 0 9568 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1712078602
transform 1 0 10856 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1712078602
transform 1 0 12144 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1712078602
transform 1 0 13432 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1712078602
transform 1 0 14720 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1712078602
transform 1 0 16008 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1712078602
transform 1 0 17296 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1712078602
transform 1 0 18584 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1712078602
transform 1 0 19872 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1712078602
transform 1 0 21160 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1712078602
transform 1 0 22448 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1712078602
transform 1 0 23736 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1712078602
transform 1 0 25024 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1712078602
transform 1 0 26312 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1712078602
transform 1 0 27600 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1712078602
transform 1 0 28888 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1712078602
transform 1 0 30176 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1712078602
transform 1 0 31464 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1712078602
transform 1 0 32752 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1712078602
transform 1 0 34040 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1712078602
transform 1 0 35328 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1712078602
transform 1 0 36616 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1712078602
transform 1 0 37904 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1712078602
transform 1 0 39192 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1712078602
transform 1 0 40480 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1712078602
transform 1 0 41768 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1712078602
transform 1 0 43056 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1712078602
transform 1 0 44344 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1712078602
transform 1 0 45632 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1712078602
transform 1 0 46920 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1712078602
transform 1 0 48208 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1712078602
transform 1 0 49496 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1712078602
transform 1 0 50784 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1712078602
transform 1 0 52072 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1712078602
transform 1 0 53360 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1712078602
transform 1 0 54648 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1712078602
transform 1 0 55936 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1712078602
transform 1 0 57224 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1712078602
transform 1 0 58512 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1712078602
transform 1 0 59800 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1712078602
transform 1 0 61088 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1712078602
transform 1 0 62376 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1712078602
transform 1 0 63664 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1712078602
transform 1 0 64952 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1712078602
transform 1 0 66240 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1712078602
transform 1 0 67528 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1712078602
transform 1 0 68816 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1712078602
transform 1 0 70104 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1712078602
transform 1 0 71392 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1712078602
transform 1 0 72680 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1712078602
transform 1 0 73968 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1712078602
transform 1 0 75256 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1712078602
transform 1 0 76544 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1712078602
transform 1 0 77832 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1712078602
transform 1 0 79120 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1712078602
transform 1 0 80408 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1712078602
transform 1 0 81696 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1712078602
transform 1 0 82984 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1712078602
transform 1 0 84272 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1712078602
transform 1 0 85560 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1712078602
transform 1 0 86848 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1712078602
transform 1 0 88136 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1712078602
transform 1 0 89424 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1712078602
transform 1 0 90712 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1712078602
transform 1 0 92000 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1712078602
transform 1 0 93288 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1712078602
transform 1 0 94576 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1712078602
transform 1 0 95864 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1712078602
transform 1 0 97152 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1712078602
transform 1 0 98440 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1712078602
transform 1 0 99728 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1712078602
transform 1 0 101016 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1712078602
transform 1 0 102304 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1712078602
transform 1 0 103592 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1712078602
transform 1 0 104880 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1712078602
transform 1 0 106168 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1712078602
transform 1 0 107456 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1712078602
transform 1 0 108744 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1712078602
transform 1 0 110032 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1712078602
transform 1 0 111320 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1712078602
transform 1 0 112608 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1712078602
transform 1 0 113896 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1712078602
transform 1 0 115184 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1712078602
transform 1 0 116472 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1712078602
transform 1 0 117760 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1712078602
transform 1 0 119048 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1712078602
transform 1 0 120336 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1712078602
transform 1 0 121624 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1712078602
transform 1 0 122912 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1712078602
transform 1 0 124200 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1712078602
transform 1 0 125488 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1712078602
transform 1 0 126776 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1712078602
transform 1 0 128064 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1712078602
transform 1 0 129352 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1712078602
transform 1 0 130640 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1712078602
transform 1 0 131928 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1712078602
transform 1 0 133216 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1712078602
transform 1 0 134504 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1712078602
transform 1 0 135792 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1712078602
transform 1 0 137080 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1712078602
transform 1 0 138368 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1712078602
transform 1 0 139656 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1712078602
transform 1 0 140944 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1712078602
transform 1 0 142232 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1712078602
transform 1 0 143520 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1712078602
transform 1 0 144808 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1712078602
transform 1 0 146096 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1712078602
transform 1 0 147384 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1712078602
transform 1 0 148672 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1712078602
transform 1 0 149960 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1712078602
transform 1 0 151248 0 1 6528
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1712078602
transform 1 0 152536 0 1 6528
box -19 -24 65 296
<< labels >>
rlabel metal4 s -538 -2 -378 7890 4 GND
port 0 nsew ground bidirectional
rlabel metal5 s -538 -2 153994 158 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -538 7730 153994 7890 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 153834 -2 153994 7890 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 38571 -2 38731 7890 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 76670 -2 76830 7890 6 GND
port 0 nsew ground bidirectional
rlabel metal4 s 114769 -2 114929 7890 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -538 2464 153994 2624 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -538 3920 153994 4080 6 GND
port 0 nsew ground bidirectional
rlabel metal5 s -538 5376 153994 5536 6 GND
port 0 nsew ground bidirectional
rlabel metal2 s 745 7600 773 8000 6 ROW_SEL[0]
port 1 nsew signal tristate
rlabel metal2 s 16063 7600 16091 8000 6 ROW_SEL[10]
port 2 nsew signal tristate
rlabel metal2 s 17627 7600 17655 8000 6 ROW_SEL[11]
port 3 nsew signal tristate
rlabel metal2 s 19145 7600 19173 8000 6 ROW_SEL[12]
port 4 nsew signal tristate
rlabel metal2 s 20663 7600 20691 8000 6 ROW_SEL[13]
port 5 nsew signal tristate
rlabel metal2 s 22227 7600 22255 8000 6 ROW_SEL[14]
port 6 nsew signal tristate
rlabel metal2 s 23745 7600 23773 8000 6 ROW_SEL[15]
port 7 nsew signal tristate
rlabel metal2 s 25263 7600 25291 8000 6 ROW_SEL[16]
port 8 nsew signal tristate
rlabel metal2 s 26827 7600 26855 8000 6 ROW_SEL[17]
port 9 nsew signal tristate
rlabel metal2 s 28345 7600 28373 8000 6 ROW_SEL[18]
port 10 nsew signal tristate
rlabel metal2 s 29909 7600 29937 8000 6 ROW_SEL[19]
port 11 nsew signal tristate
rlabel metal2 s 2263 7600 2291 8000 6 ROW_SEL[1]
port 12 nsew signal tristate
rlabel metal2 s 31427 7600 31455 8000 6 ROW_SEL[20]
port 13 nsew signal tristate
rlabel metal2 s 32945 7600 32973 8000 6 ROW_SEL[21]
port 14 nsew signal tristate
rlabel metal2 s 34509 7600 34537 8000 6 ROW_SEL[22]
port 15 nsew signal tristate
rlabel metal2 s 36027 7600 36055 8000 6 ROW_SEL[23]
port 16 nsew signal tristate
rlabel metal2 s 37545 7600 37573 8000 6 ROW_SEL[24]
port 17 nsew signal tristate
rlabel metal2 s 39109 7600 39137 8000 6 ROW_SEL[25]
port 18 nsew signal tristate
rlabel metal2 s 40627 7600 40655 8000 6 ROW_SEL[26]
port 19 nsew signal tristate
rlabel metal2 s 42145 7600 42173 8000 6 ROW_SEL[27]
port 20 nsew signal tristate
rlabel metal2 s 43709 7600 43737 8000 6 ROW_SEL[28]
port 21 nsew signal tristate
rlabel metal2 s 45227 7600 45255 8000 6 ROW_SEL[29]
port 22 nsew signal tristate
rlabel metal2 s 3781 7600 3809 8000 6 ROW_SEL[2]
port 23 nsew signal tristate
rlabel metal2 s 46791 7600 46819 8000 6 ROW_SEL[30]
port 24 nsew signal tristate
rlabel metal2 s 48309 7600 48337 8000 6 ROW_SEL[31]
port 25 nsew signal tristate
rlabel metal2 s 49827 7600 49855 8000 6 ROW_SEL[32]
port 26 nsew signal tristate
rlabel metal2 s 51391 7600 51419 8000 6 ROW_SEL[33]
port 27 nsew signal tristate
rlabel metal2 s 52909 7600 52937 8000 6 ROW_SEL[34]
port 28 nsew signal tristate
rlabel metal2 s 54427 7600 54455 8000 6 ROW_SEL[35]
port 29 nsew signal tristate
rlabel metal2 s 55991 7600 56019 8000 6 ROW_SEL[36]
port 30 nsew signal tristate
rlabel metal2 s 57509 7600 57537 8000 6 ROW_SEL[37]
port 31 nsew signal tristate
rlabel metal2 s 59073 7600 59101 8000 6 ROW_SEL[38]
port 32 nsew signal tristate
rlabel metal2 s 60591 7600 60619 8000 6 ROW_SEL[39]
port 33 nsew signal tristate
rlabel metal2 s 5345 7600 5373 8000 6 ROW_SEL[3]
port 34 nsew signal tristate
rlabel metal2 s 62109 7600 62137 8000 6 ROW_SEL[40]
port 35 nsew signal tristate
rlabel metal2 s 63673 7600 63701 8000 6 ROW_SEL[41]
port 36 nsew signal tristate
rlabel metal2 s 65191 7600 65219 8000 6 ROW_SEL[42]
port 37 nsew signal tristate
rlabel metal2 s 66709 7600 66737 8000 6 ROW_SEL[43]
port 38 nsew signal tristate
rlabel metal2 s 68273 7600 68301 8000 6 ROW_SEL[44]
port 39 nsew signal tristate
rlabel metal2 s 69791 7600 69819 8000 6 ROW_SEL[45]
port 40 nsew signal tristate
rlabel metal2 s 71355 7600 71383 8000 6 ROW_SEL[46]
port 41 nsew signal tristate
rlabel metal2 s 72873 7600 72901 8000 6 ROW_SEL[47]
port 42 nsew signal tristate
rlabel metal2 s 74391 7600 74419 8000 6 ROW_SEL[48]
port 43 nsew signal tristate
rlabel metal2 s 75955 7600 75983 8000 6 ROW_SEL[49]
port 44 nsew signal tristate
rlabel metal2 s 6863 7600 6891 8000 6 ROW_SEL[4]
port 45 nsew signal tristate
rlabel metal2 s 77473 7600 77501 8000 6 ROW_SEL[50]
port 46 nsew signal tristate
rlabel metal2 s 78991 7600 79019 8000 6 ROW_SEL[51]
port 47 nsew signal tristate
rlabel metal2 s 80555 7600 80583 8000 6 ROW_SEL[52]
port 48 nsew signal tristate
rlabel metal2 s 82073 7600 82101 8000 6 ROW_SEL[53]
port 49 nsew signal tristate
rlabel metal2 s 83591 7600 83619 8000 6 ROW_SEL[54]
port 50 nsew signal tristate
rlabel metal2 s 85155 7600 85183 8000 6 ROW_SEL[55]
port 51 nsew signal tristate
rlabel metal2 s 86673 7600 86701 8000 6 ROW_SEL[56]
port 52 nsew signal tristate
rlabel metal2 s 88237 7600 88265 8000 6 ROW_SEL[57]
port 53 nsew signal tristate
rlabel metal2 s 89755 7600 89783 8000 6 ROW_SEL[58]
port 54 nsew signal tristate
rlabel metal2 s 91273 7600 91301 8000 6 ROW_SEL[59]
port 55 nsew signal tristate
rlabel metal2 s 8381 7600 8409 8000 6 ROW_SEL[5]
port 56 nsew signal tristate
rlabel metal2 s 92837 7600 92865 8000 6 ROW_SEL[60]
port 57 nsew signal tristate
rlabel metal2 s 94355 7600 94383 8000 6 ROW_SEL[61]
port 58 nsew signal tristate
rlabel metal2 s 95873 7600 95901 8000 6 ROW_SEL[62]
port 59 nsew signal tristate
rlabel metal2 s 97437 7600 97465 8000 6 ROW_SEL[63]
port 60 nsew signal tristate
rlabel metal2 s 98955 7600 98983 8000 6 ROW_SEL[64]
port 61 nsew signal tristate
rlabel metal2 s 100519 7600 100547 8000 6 ROW_SEL[65]
port 62 nsew signal tristate
rlabel metal2 s 102037 7600 102065 8000 6 ROW_SEL[66]
port 63 nsew signal tristate
rlabel metal2 s 103555 7600 103583 8000 6 ROW_SEL[67]
port 64 nsew signal tristate
rlabel metal2 s 105119 7600 105147 8000 6 ROW_SEL[68]
port 65 nsew signal tristate
rlabel metal2 s 106637 7600 106665 8000 6 ROW_SEL[69]
port 66 nsew signal tristate
rlabel metal2 s 9945 7600 9973 8000 6 ROW_SEL[6]
port 67 nsew signal tristate
rlabel metal2 s 108155 7600 108183 8000 6 ROW_SEL[70]
port 68 nsew signal tristate
rlabel metal2 s 109719 7600 109747 8000 6 ROW_SEL[71]
port 69 nsew signal tristate
rlabel metal2 s 111237 7600 111265 8000 6 ROW_SEL[72]
port 70 nsew signal tristate
rlabel metal2 s 112801 7600 112829 8000 6 ROW_SEL[73]
port 71 nsew signal tristate
rlabel metal2 s 114319 7600 114347 8000 6 ROW_SEL[74]
port 72 nsew signal tristate
rlabel metal2 s 115837 7600 115865 8000 6 ROW_SEL[75]
port 73 nsew signal tristate
rlabel metal2 s 117401 7600 117429 8000 6 ROW_SEL[76]
port 74 nsew signal tristate
rlabel metal2 s 118919 7600 118947 8000 6 ROW_SEL[77]
port 75 nsew signal tristate
rlabel metal2 s 120437 7600 120465 8000 6 ROW_SEL[78]
port 76 nsew signal tristate
rlabel metal2 s 122001 7600 122029 8000 6 ROW_SEL[79]
port 77 nsew signal tristate
rlabel metal2 s 11463 7600 11491 8000 6 ROW_SEL[7]
port 78 nsew signal tristate
rlabel metal2 s 123519 7600 123547 8000 6 ROW_SEL[80]
port 79 nsew signal tristate
rlabel metal2 s 125037 7600 125065 8000 6 ROW_SEL[81]
port 80 nsew signal tristate
rlabel metal2 s 126601 7600 126629 8000 6 ROW_SEL[82]
port 81 nsew signal tristate
rlabel metal2 s 128119 7600 128147 8000 6 ROW_SEL[83]
port 82 nsew signal tristate
rlabel metal2 s 129683 7600 129711 8000 6 ROW_SEL[84]
port 83 nsew signal tristate
rlabel metal2 s 131201 7600 131229 8000 6 ROW_SEL[85]
port 84 nsew signal tristate
rlabel metal2 s 132719 7600 132747 8000 6 ROW_SEL[86]
port 85 nsew signal tristate
rlabel metal2 s 134283 7600 134311 8000 6 ROW_SEL[87]
port 86 nsew signal tristate
rlabel metal2 s 135801 7600 135829 8000 6 ROW_SEL[88]
port 87 nsew signal tristate
rlabel metal2 s 137319 7600 137347 8000 6 ROW_SEL[89]
port 88 nsew signal tristate
rlabel metal2 s 12981 7600 13009 8000 6 ROW_SEL[8]
port 89 nsew signal tristate
rlabel metal2 s 138883 7600 138911 8000 6 ROW_SEL[90]
port 90 nsew signal tristate
rlabel metal2 s 140401 7600 140429 8000 6 ROW_SEL[91]
port 91 nsew signal tristate
rlabel metal2 s 141965 7600 141993 8000 6 ROW_SEL[92]
port 92 nsew signal tristate
rlabel metal2 s 143483 7600 143511 8000 6 ROW_SEL[93]
port 93 nsew signal tristate
rlabel metal2 s 145001 7600 145029 8000 6 ROW_SEL[94]
port 94 nsew signal tristate
rlabel metal2 s 146565 7600 146593 8000 6 ROW_SEL[95]
port 95 nsew signal tristate
rlabel metal2 s 148083 7600 148111 8000 6 ROW_SEL[96]
port 96 nsew signal tristate
rlabel metal2 s 149601 7600 149629 8000 6 ROW_SEL[97]
port 97 nsew signal tristate
rlabel metal2 s 151165 7600 151193 8000 6 ROW_SEL[98]
port 98 nsew signal tristate
rlabel metal2 s 152683 7600 152711 8000 6 ROW_SEL[99]
port 99 nsew signal tristate
rlabel metal2 s 14545 7600 14573 8000 6 ROW_SEL[9]
port 100 nsew signal tristate
rlabel metal4 s -208 328 -48 7560 4 VDD
port 101 nsew power bidirectional
rlabel metal5 s -208 328 153664 488 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -208 7400 153664 7560 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 153504 328 153664 7560 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 19521 -2 19681 7890 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 57620 -2 57780 7890 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 95719 -2 95879 7890 6 VDD
port 101 nsew power bidirectional
rlabel metal4 s 133818 -2 133978 7890 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -538 1736 153994 1896 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -538 3192 153994 3352 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -538 4648 153994 4808 6 VDD
port 101 nsew power bidirectional
rlabel metal5 s -538 6104 153994 6264 6 VDD
port 101 nsew power bidirectional
rlabel metal3 s 153100 956 153500 1016 6 clk
port 102 nsew signal input
rlabel metal3 s 153100 6940 153500 7000 6 data_in
port 103 nsew signal input
rlabel metal3 s 0 4016 400 4076 6 data_out
port 104 nsew signal tristate
rlabel metal3 s 153100 2928 153500 2988 6 ena
port 105 nsew signal input
rlabel metal3 s 153100 4968 153500 5028 6 rst
port 106 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 153500 8000
<< end >>
