magic
tech sky130A
timestamp 1758130718
<< metal5 >>
rect 18800 56200 21000 56400
rect 22700 56200 23000 56400
rect 51100 56200 51600 56400
rect 18400 55900 21500 56200
rect 22600 55900 23200 56200
rect 23900 55900 30700 56200
rect 18000 55700 21800 55900
rect 22400 55700 23200 55900
rect 23800 55700 30700 55900
rect 31700 55900 34100 56200
rect 37600 55900 40700 56200
rect 41000 55900 45600 56200
rect 31700 55700 34200 55900
rect 17800 55400 23200 55700
rect 23900 55400 30800 55700
rect 31700 55400 34300 55700
rect 37600 55400 40800 55900
rect 40960 55700 46100 55900
rect 51100 55700 51700 56200
rect 41000 55400 46600 55700
rect 17500 55100 23200 55400
rect 24500 55100 30800 55400
rect 32300 55100 34400 55400
rect 38200 55100 40300 55400
rect 41500 55100 46800 55400
rect 51000 55100 51800 55700
rect 17400 54900 19300 55100
rect 20800 54900 23200 55100
rect 24700 54900 30800 55100
rect 32500 54900 34600 55100
rect 17200 54600 19100 54900
rect 21100 54600 23200 54900
rect 17000 54400 18700 54600
rect 21400 54400 23200 54600
rect 24800 54400 26400 54900
rect 29400 54600 30800 54900
rect 32600 54600 34600 54900
rect 38500 54900 40000 55100
rect 41900 54900 46900 55100
rect 38500 54600 39800 54900
rect 29900 54400 30800 54600
rect 32800 54400 34700 54600
rect 16900 54100 18600 54400
rect 21600 54100 23200 54400
rect 16800 53800 18400 54100
rect 21700 53800 23200 54100
rect 16700 53600 18200 53800
rect 21800 53600 23200 53800
rect 16600 53300 18100 53600
rect 22000 53300 23200 53600
rect 16400 53100 18000 53300
rect 22100 53100 23200 53300
rect 16300 52800 17900 53100
rect 16200 52500 17900 52800
rect 22200 52500 23200 53100
rect 16200 52300 17800 52500
rect 22300 52300 23200 52500
rect 16100 52000 17600 52300
rect 16000 51800 17600 52000
rect 22400 51800 23200 52300
rect 16000 51500 17500 51800
rect 15800 51000 17400 51500
rect 22600 51200 23200 51800
rect 15700 50700 17400 51000
rect 15700 50200 17300 50700
rect 22700 50400 23300 51200
rect 15600 49900 17300 50200
rect 22800 50200 23300 50400
rect 22800 49900 23200 50200
rect 15600 49400 17200 49900
rect 15500 48400 17200 49400
rect 15500 47600 17000 48400
rect 6400 45160 6600 46300
rect 15400 46000 17000 47600
rect 6340 45000 6600 45160
rect 15500 45000 17000 46000
rect 25000 48100 26400 54400
rect 30000 54100 30800 54400
rect 30100 53300 30800 54100
rect 30200 52800 30800 53300
rect 30400 52000 30800 52800
rect 32900 54100 34800 54400
rect 38600 54100 39700 54600
rect 42000 54100 43600 54900
rect 44900 54600 47200 54900
rect 45400 54400 47400 54600
rect 50900 54400 52000 55100
rect 45600 54100 47400 54400
rect 32900 53800 34900 54100
rect 38800 53800 39700 54100
rect 32900 53600 35000 53800
rect 32900 53100 35200 53600
rect 32900 52800 35300 53100
rect 32900 52500 35400 52800
rect 32900 52300 35500 52500
rect 32900 52000 35600 52300
rect 32900 51640 33540 52000
rect 33700 51800 35600 52000
rect 29600 49900 30100 50700
rect 29500 49100 30100 49900
rect 32900 49400 33600 51640
rect 33800 51500 35800 51800
rect 34000 51200 35900 51500
rect 34100 51000 36000 51200
rect 34100 50700 36100 51000
rect 34200 50400 36100 50700
rect 34300 50200 36200 50400
rect 34400 49900 36400 50200
rect 34600 49700 36500 49900
rect 29400 48600 30100 49100
rect 29300 48400 30100 48600
rect 29200 48100 30100 48400
rect 25000 46800 30100 48100
rect 6200 44200 6500 45000
rect 15500 44200 17200 45000
rect 6100 43560 6400 44200
rect 7800 43900 8400 44200
rect 7600 43857 8400 43900
rect 7600 43700 8500 43857
rect 6040 43400 6400 43560
rect 7400 43400 7800 43700
rect 6100 42400 6260 43400
rect 7200 43100 7700 43400
rect 7100 42900 7400 43100
rect 7000 42760 7300 42900
rect 8300 42760 8500 43700
rect 15600 43700 17200 44200
rect 15600 43400 17300 43700
rect 6940 42600 7300 42760
rect 8240 42600 8500 42760
rect 15700 42900 17300 43400
rect 15700 42600 17400 42900
rect 6700 42400 7100 42600
rect 6100 42100 7000 42400
rect 6200 41800 6700 42100
rect 8200 41800 8400 42600
rect 15800 42400 17400 42600
rect 15800 42100 17500 42400
rect 8000 41600 8400 41800
rect 16000 41800 17500 42100
rect 16000 41600 17600 41800
rect 8000 41100 8300 41600
rect 9700 41300 10100 41600
rect 16100 41300 17800 41600
rect 9500 41100 10300 41300
rect 16200 41100 17800 41300
rect 22900 41100 23300 41300
rect 7900 40800 8300 41100
rect 9400 40800 10400 41100
rect 16200 40800 17900 41100
rect 22800 40800 23400 41100
rect 7900 39500 8200 40800
rect 9100 40500 9800 40800
rect 10000 40500 10400 40800
rect 16300 40500 18000 40800
rect 22700 40500 23400 40800
rect 9000 40300 9600 40500
rect 8900 40000 9400 40300
rect 10100 40000 10400 40500
rect 16400 40300 18100 40500
rect 22600 40300 23300 40500
rect 8600 39800 9200 40000
rect 8500 39500 9100 39800
rect 10000 39500 10400 40000
rect 16600 40000 18200 40300
rect 22300 40000 23200 40300
rect 16600 39800 18400 40000
rect 22200 39800 23000 40000
rect 16700 39500 18600 39800
rect 22000 39500 22900 39800
rect 7900 39200 8900 39500
rect 8000 39000 8600 39200
rect 10000 39000 10300 39500
rect 16800 39200 18700 39500
rect 21700 39200 22800 39500
rect 25000 39200 26400 46800
rect 28700 46500 30100 46800
rect 29200 46300 30100 46500
rect 29300 46000 30100 46300
rect 29400 45500 30100 46000
rect 29500 44700 30100 45500
rect 29600 44200 30100 44700
rect 29600 43900 30000 44200
rect 31100 42400 31400 42600
rect 31000 42100 31400 42400
rect 30800 41600 31400 42100
rect 30700 41300 31400 41600
rect 30700 41100 31300 41300
rect 33000 41100 33600 49400
rect 34700 49100 36600 49700
rect 34800 48900 36700 49100
rect 34900 48600 36800 48900
rect 35000 48400 37000 48600
rect 35200 48100 37000 48400
rect 35200 47800 37100 48100
rect 35300 47600 37200 47800
rect 35400 47300 37300 47600
rect 35500 47100 37400 47300
rect 35600 46500 37600 47100
rect 35800 46300 37700 46500
rect 35900 46000 37800 46300
rect 36000 45800 37900 46000
rect 36100 45200 38000 45800
rect 36200 45000 38200 45200
rect 36400 44700 38300 45000
rect 36500 44400 38300 44700
rect 36600 44200 38400 44400
rect 38800 44200 39600 53800
rect 42100 47800 43600 54100
rect 45700 53800 47500 54100
rect 50800 53800 52100 54400
rect 45800 53600 47600 53800
rect 46000 53300 47800 53600
rect 50600 53300 52200 53800
rect 46100 53100 47800 53300
rect 46200 52300 47900 53100
rect 50500 52500 52300 53300
rect 46300 49700 48000 52300
rect 50400 52000 52400 52500
rect 50300 51500 50940 52000
rect 51100 51500 52600 52000
rect 50300 51200 50900 51500
rect 50200 51000 50900 51200
rect 51200 51000 52700 51500
rect 50200 50700 50800 51000
rect 50000 50200 50800 50700
rect 51400 50700 52700 51000
rect 51400 50200 52800 50700
rect 49900 49700 50600 50200
rect 51500 49700 52900 50200
rect 46300 49400 47900 49700
rect 46200 48900 47900 49400
rect 49800 49400 50600 49700
rect 49800 48900 50500 49400
rect 51600 49100 53000 49700
rect 51600 48900 53200 49100
rect 46100 48400 47800 48900
rect 49700 48400 50400 48900
rect 51700 48400 53200 48900
rect 46000 48100 47600 48400
rect 49600 48100 50400 48400
rect 45800 47800 47500 48100
rect 42100 47100 43400 47800
rect 45700 47600 47400 47800
rect 49600 47600 50300 48100
rect 51800 47800 53300 48400
rect 45500 47300 47300 47600
rect 45100 47100 47200 47300
rect 49400 47100 50200 47600
rect 52000 47300 53400 47800
rect 52000 47100 53500 47300
rect 42100 46800 43900 47100
rect 44200 46800 46900 47100
rect 49300 46800 50200 47100
rect 52100 46800 53500 47100
rect 42100 46500 46700 46800
rect 49300 46500 50000 46800
rect 52100 46500 53600 46800
rect 42100 46300 46600 46500
rect 49200 46300 50000 46500
rect 42100 46000 46200 46300
rect 42100 45800 45700 46000
rect 49200 45800 49900 46300
rect 52200 46000 53600 46500
rect 42100 45500 43600 45800
rect 42100 45000 43400 45500
rect 49100 45200 49800 45800
rect 52300 45500 53800 46000
rect 52300 45200 53900 45500
rect 49000 45000 49800 45200
rect 52400 45000 53900 45200
rect 36600 43900 38500 44200
rect 36700 43700 38500 43900
rect 36800 43400 38600 43700
rect 38800 43400 39500 44200
rect 37000 43100 39500 43400
rect 37100 42900 39500 43100
rect 37200 42400 39500 42900
rect 37300 42100 39500 42400
rect 37400 41800 39500 42100
rect 37600 41300 39500 41800
rect 37700 41100 39500 41300
rect 30600 40800 31300 41100
rect 30500 40500 31300 40800
rect 30500 40300 31200 40500
rect 30400 40000 31200 40300
rect 30200 39800 31200 40000
rect 30000 39500 31200 39800
rect 32900 39500 33700 41100
rect 37800 40800 39500 41100
rect 37900 40500 39500 40800
rect 38000 40300 39500 40500
rect 38200 39800 39500 40300
rect 42100 39800 43600 45000
rect 49000 44700 54000 45000
rect 48800 44400 54000 44700
rect 48800 43900 54100 44400
rect 48700 43700 54100 43900
rect 48700 43400 49400 43700
rect 48600 42900 49400 43400
rect 52700 43100 54200 43700
rect 48500 42100 49300 42900
rect 52800 42600 54400 43100
rect 52900 42400 54400 42600
rect 48400 41600 49200 42100
rect 52900 41800 54500 42400
rect 48200 41300 49200 41600
rect 53000 41300 54600 41800
rect 48200 41100 49100 41300
rect 48100 40800 49100 41100
rect 53200 40800 54700 41300
rect 48100 40500 49000 40800
rect 48000 40300 49000 40500
rect 48000 40000 48800 40300
rect 53300 40000 54800 40800
rect 38300 39500 39500 39800
rect 29800 39200 31100 39500
rect 17000 39000 19000 39200
rect 21500 39000 22700 39200
rect 24800 39000 26500 39200
rect 29300 39000 31100 39200
rect 32800 39000 33800 39500
rect 38400 39200 39500 39500
rect 38500 39000 39500 39200
rect 42000 39200 43600 39800
rect 47900 39500 48800 40000
rect 42000 39000 43700 39200
rect 47800 39000 48800 39500
rect 8200 38700 8400 39000
rect 9800 38400 10200 39000
rect 17200 38700 19400 39000
rect 21000 38700 22400 39000
rect 24700 38700 31100 39000
rect 32600 38700 34000 39000
rect 11400 38400 12100 38700
rect 17300 38400 22300 38700
rect 24600 38400 31000 38700
rect 32400 38400 34200 38700
rect 38600 38400 39500 39000
rect 41900 38700 43700 39000
rect 47600 38700 48800 39000
rect 53400 39500 55000 40000
rect 53400 39200 55100 39500
rect 53400 38700 55200 39200
rect 41800 38400 43900 38700
rect 47400 38400 49000 38700
rect 53300 38400 55400 38700
rect 9700 37700 10200 38400
rect 11300 38200 12200 38400
rect 17500 38200 22100 38400
rect 23900 38200 31000 38400
rect 31800 38200 34800 38400
rect 38800 38200 39500 38400
rect 11000 37900 12200 38200
rect 17800 37900 21800 38200
rect 23800 37900 31000 38200
rect 10900 37700 12400 37900
rect 18000 37700 21600 37900
rect 23900 37700 31000 37900
rect 31700 37700 34800 38200
rect 38900 37900 39500 38200
rect 39000 37700 39500 37900
rect 41000 38200 44600 38400
rect 47000 38200 49600 38400
rect 52600 38200 55800 38400
rect 41000 37700 44800 38200
rect 46900 37700 49700 38200
rect 52600 37700 55900 38200
rect 9700 36900 10100 37700
rect 10800 37400 11500 37700
rect 10600 37100 11400 37400
rect 11900 37100 12400 37700
rect 18400 37400 21200 37700
rect 19000 37100 20800 37400
rect 39100 37100 39500 37700
rect 10400 36900 11200 37100
rect 11800 36900 12400 37100
rect 9700 36600 11000 36900
rect 9700 36400 10800 36600
rect 11800 36400 12200 36900
rect 9700 36100 10700 36400
rect 10000 35800 10400 36100
rect 11600 35800 12200 36400
rect 13400 35800 13900 36100
rect 11600 35600 12100 35800
rect 13200 35600 14000 35800
rect 11500 35100 12100 35600
rect 13000 35300 14200 35600
rect 12800 35100 14200 35300
rect 11500 34500 12000 35100
rect 12700 34800 14300 35100
rect 12500 34500 13400 34800
rect 11400 34460 12000 34500
rect 11400 34000 11940 34460
rect 12400 34300 13300 34500
rect 13700 34300 14300 34800
rect 12100 34000 13100 34300
rect 13600 34000 14300 34300
rect 11400 33800 13000 34000
rect 11500 33500 12800 33800
rect 13600 33500 14200 34000
rect 11500 33200 12600 33500
rect 13400 33200 14200 33500
rect 11600 33000 12400 33200
rect 13400 32700 14000 33200
rect 13300 32200 14000 32700
rect 57500 33000 57700 33200
rect 57500 32700 58000 33000
rect 57500 32400 58300 32700
rect 57600 32200 58600 32400
rect 13300 31400 13900 32200
rect 57600 31900 58800 32200
rect 57700 31700 59200 31900
rect 57700 31400 59400 31700
rect 13300 31100 59600 31400
rect 13300 30900 59900 31100
rect 13200 30600 59800 30900
rect 13000 30400 59500 30600
rect 12800 30100 13700 30400
rect 57700 30100 59200 30400
rect 12700 29800 13600 30100
rect 57600 29800 58900 30100
rect 12600 29600 13400 29800
rect 57600 29600 58600 29800
rect 12400 29300 13200 29600
rect 57500 29300 58300 29600
rect 12200 29100 13100 29300
rect 57500 29100 58100 29300
rect 12100 28800 13000 29100
rect 57500 28800 57700 29100
rect 11900 28500 12800 28800
rect 11800 28300 12600 28500
rect 11600 28000 12500 28300
rect 11500 27800 12400 28000
rect 11300 27500 12100 27800
rect 11200 27200 12000 27500
rect 11000 27000 11900 27200
rect 10900 26700 11800 27000
rect 10700 26400 11500 26700
rect 10600 26200 11400 26400
rect 10400 25900 11300 26200
rect 10200 25700 11200 25900
rect 10100 25400 10900 25700
rect 10000 25100 10800 25400
rect 9800 24900 10700 25100
rect 9600 24600 10400 24900
rect 9500 24400 10300 24600
rect 9400 24100 10200 24400
rect 9200 23800 10100 24100
rect 9100 23600 10000 23800
rect 8900 23300 9700 23600
rect 8800 23100 9600 23300
rect 8600 22800 9500 23100
rect 8500 22500 9200 22800
rect 8300 22300 9100 22500
rect 8200 22000 9000 22300
rect 8000 21800 8900 22000
rect 7800 21500 8600 21800
rect 7700 21200 8500 21500
rect 7600 21000 8400 21200
rect 7400 20700 8200 21000
rect 7200 20400 8000 20700
rect 7100 20200 7900 20400
rect 7000 19900 7800 20200
rect 6700 19700 7600 19900
rect 6600 19400 7400 19700
rect 6500 19100 7300 19400
rect 6400 18900 7200 19100
rect 6100 18600 7000 18900
rect 6000 18400 6800 18600
rect 5900 18100 6700 18400
rect 5600 17800 6500 18100
rect 5500 17600 6400 17800
rect 4100 17100 4300 17600
rect 5400 17300 6200 17600
rect 5300 17100 6100 17300
rect 4000 16500 4300 17100
rect 5000 16800 5900 17100
rect 4900 16500 5800 16800
rect 3800 16000 4400 16500
rect 4800 16300 5600 16500
rect 4700 16000 5500 16300
rect 3700 15800 5300 16000
rect 3600 15500 5200 15800
rect 3600 15200 5000 15500
rect 3500 15000 4800 15200
rect 3500 14700 4900 15000
rect 3400 14400 5000 14700
rect 3400 14200 5300 14400
rect 3200 13900 5400 14200
rect 3200 13700 5300 13900
rect 3100 13400 4900 13700
rect 3000 13100 4400 13400
rect 3000 12900 4000 13100
rect 2900 12600 3600 12900
rect 2900 12400 3100 12600
<< end >>
