magic
tech sky130A
timestamp 1757995770
<< nmoslvt >>
rect 270 -148900 1070 -148700
rect 1770 -148900 2570 -148700
rect 3270 -148900 4070 -148700
rect 4770 -148900 5570 -148700
rect 6270 -148900 7070 -148700
rect 7770 -148900 8570 -148700
rect 9270 -148900 10070 -148700
rect 10770 -148900 11570 -148700
rect 12270 -148900 13070 -148700
rect 13770 -148900 14570 -148700
rect 15270 -148900 16070 -148700
rect 16770 -148900 17570 -148700
rect 18270 -148900 19070 -148700
rect 19770 -148900 20570 -148700
rect 21270 -148900 22070 -148700
rect 22770 -148900 23570 -148700
rect 24270 -148900 25070 -148700
rect 25770 -148900 26570 -148700
rect 27270 -148900 28070 -148700
rect 28770 -148900 29570 -148700
rect 30270 -148900 31070 -148700
rect 31770 -148900 32570 -148700
rect 33270 -148900 34070 -148700
rect 34770 -148900 35570 -148700
rect 36270 -148900 37070 -148700
rect 37770 -148900 38570 -148700
rect 39270 -148900 40070 -148700
rect 40770 -148900 41570 -148700
rect 42270 -148900 43070 -148700
rect 43770 -148900 44570 -148700
rect 45270 -148900 46070 -148700
rect 46770 -148900 47570 -148700
rect 48270 -148900 49070 -148700
rect 49770 -148900 50570 -148700
rect 51270 -148900 52070 -148700
rect 52770 -148900 53570 -148700
rect 54270 -148900 55070 -148700
rect 55770 -148900 56570 -148700
rect 57270 -148900 58070 -148700
rect 58770 -148900 59570 -148700
rect 60270 -148900 61070 -148700
rect 61770 -148900 62570 -148700
rect 63270 -148900 64070 -148700
rect 64770 -148900 65570 -148700
rect 66270 -148900 67070 -148700
rect 67770 -148900 68570 -148700
rect 69270 -148900 70070 -148700
rect 70770 -148900 71570 -148700
rect 72270 -148900 73070 -148700
rect 73770 -148900 74570 -148700
rect 75270 -148900 76070 -148700
rect 76770 -148900 77570 -148700
rect 78270 -148900 79070 -148700
rect 79770 -148900 80570 -148700
rect 81270 -148900 82070 -148700
rect 82770 -148900 83570 -148700
rect 84270 -148900 85070 -148700
rect 85770 -148900 86570 -148700
rect 87270 -148900 88070 -148700
rect 88770 -148900 89570 -148700
rect 90270 -148900 91070 -148700
rect 91770 -148900 92570 -148700
rect 93270 -148900 94070 -148700
rect 94770 -148900 95570 -148700
rect 96270 -148900 97070 -148700
rect 97770 -148900 98570 -148700
rect 99270 -148900 100070 -148700
rect 100770 -148900 101570 -148700
rect 102270 -148900 103070 -148700
rect 103770 -148900 104570 -148700
rect 105270 -148900 106070 -148700
rect 106770 -148900 107570 -148700
rect 108270 -148900 109070 -148700
rect 109770 -148900 110570 -148700
rect 111270 -148900 112070 -148700
rect 112770 -148900 113570 -148700
rect 114270 -148900 115070 -148700
rect 115770 -148900 116570 -148700
rect 117270 -148900 118070 -148700
rect 118770 -148900 119570 -148700
rect 120270 -148900 121070 -148700
rect 121770 -148900 122570 -148700
rect 123270 -148900 124070 -148700
rect 124770 -148900 125570 -148700
rect 126270 -148900 127070 -148700
rect 127770 -148900 128570 -148700
rect 129270 -148900 130070 -148700
rect 130770 -148900 131570 -148700
rect 132270 -148900 133070 -148700
rect 133770 -148900 134570 -148700
rect 135270 -148900 136070 -148700
rect 136770 -148900 137570 -148700
rect 138270 -148900 139070 -148700
rect 139770 -148900 140570 -148700
rect 141270 -148900 142070 -148700
rect 142770 -148900 143570 -148700
rect 144270 -148900 145070 -148700
rect 145770 -148900 146570 -148700
rect 147270 -148900 148070 -148700
rect 148770 -148900 149570 -148700
<< ndiff >>
rect 270 -148660 1070 -148650
rect 270 -148690 280 -148660
rect 1060 -148690 1070 -148660
rect 270 -148700 1070 -148690
rect 1770 -148660 2570 -148650
rect 1770 -148690 1780 -148660
rect 2560 -148690 2570 -148660
rect 1770 -148700 2570 -148690
rect 3270 -148660 4070 -148650
rect 3270 -148690 3280 -148660
rect 4060 -148690 4070 -148660
rect 3270 -148700 4070 -148690
rect 4770 -148660 5570 -148650
rect 4770 -148690 4780 -148660
rect 5560 -148690 5570 -148660
rect 4770 -148700 5570 -148690
rect 6270 -148660 7070 -148650
rect 6270 -148690 6280 -148660
rect 7060 -148690 7070 -148660
rect 6270 -148700 7070 -148690
rect 7770 -148660 8570 -148650
rect 7770 -148690 7780 -148660
rect 8560 -148690 8570 -148660
rect 7770 -148700 8570 -148690
rect 9270 -148660 10070 -148650
rect 9270 -148690 9280 -148660
rect 10060 -148690 10070 -148660
rect 9270 -148700 10070 -148690
rect 10770 -148660 11570 -148650
rect 10770 -148690 10780 -148660
rect 11560 -148690 11570 -148660
rect 10770 -148700 11570 -148690
rect 12270 -148660 13070 -148650
rect 12270 -148690 12280 -148660
rect 13060 -148690 13070 -148660
rect 12270 -148700 13070 -148690
rect 13770 -148660 14570 -148650
rect 13770 -148690 13780 -148660
rect 14560 -148690 14570 -148660
rect 13770 -148700 14570 -148690
rect 15270 -148660 16070 -148650
rect 15270 -148690 15280 -148660
rect 16060 -148690 16070 -148660
rect 15270 -148700 16070 -148690
rect 16770 -148660 17570 -148650
rect 16770 -148690 16780 -148660
rect 17560 -148690 17570 -148660
rect 16770 -148700 17570 -148690
rect 18270 -148660 19070 -148650
rect 18270 -148690 18280 -148660
rect 19060 -148690 19070 -148660
rect 18270 -148700 19070 -148690
rect 19770 -148660 20570 -148650
rect 19770 -148690 19780 -148660
rect 20560 -148690 20570 -148660
rect 19770 -148700 20570 -148690
rect 21270 -148660 22070 -148650
rect 21270 -148690 21280 -148660
rect 22060 -148690 22070 -148660
rect 21270 -148700 22070 -148690
rect 22770 -148660 23570 -148650
rect 22770 -148690 22780 -148660
rect 23560 -148690 23570 -148660
rect 22770 -148700 23570 -148690
rect 24270 -148660 25070 -148650
rect 24270 -148690 24280 -148660
rect 25060 -148690 25070 -148660
rect 24270 -148700 25070 -148690
rect 25770 -148660 26570 -148650
rect 25770 -148690 25780 -148660
rect 26560 -148690 26570 -148660
rect 25770 -148700 26570 -148690
rect 27270 -148660 28070 -148650
rect 27270 -148690 27280 -148660
rect 28060 -148690 28070 -148660
rect 27270 -148700 28070 -148690
rect 28770 -148660 29570 -148650
rect 28770 -148690 28780 -148660
rect 29560 -148690 29570 -148660
rect 28770 -148700 29570 -148690
rect 30270 -148660 31070 -148650
rect 30270 -148690 30280 -148660
rect 31060 -148690 31070 -148660
rect 30270 -148700 31070 -148690
rect 31770 -148660 32570 -148650
rect 31770 -148690 31780 -148660
rect 32560 -148690 32570 -148660
rect 31770 -148700 32570 -148690
rect 33270 -148660 34070 -148650
rect 33270 -148690 33280 -148660
rect 34060 -148690 34070 -148660
rect 33270 -148700 34070 -148690
rect 34770 -148660 35570 -148650
rect 34770 -148690 34780 -148660
rect 35560 -148690 35570 -148660
rect 34770 -148700 35570 -148690
rect 36270 -148660 37070 -148650
rect 36270 -148690 36280 -148660
rect 37060 -148690 37070 -148660
rect 36270 -148700 37070 -148690
rect 37770 -148660 38570 -148650
rect 37770 -148690 37780 -148660
rect 38560 -148690 38570 -148660
rect 37770 -148700 38570 -148690
rect 39270 -148660 40070 -148650
rect 39270 -148690 39280 -148660
rect 40060 -148690 40070 -148660
rect 39270 -148700 40070 -148690
rect 40770 -148660 41570 -148650
rect 40770 -148690 40780 -148660
rect 41560 -148690 41570 -148660
rect 40770 -148700 41570 -148690
rect 42270 -148660 43070 -148650
rect 42270 -148690 42280 -148660
rect 43060 -148690 43070 -148660
rect 42270 -148700 43070 -148690
rect 43770 -148660 44570 -148650
rect 43770 -148690 43780 -148660
rect 44560 -148690 44570 -148660
rect 43770 -148700 44570 -148690
rect 45270 -148660 46070 -148650
rect 45270 -148690 45280 -148660
rect 46060 -148690 46070 -148660
rect 45270 -148700 46070 -148690
rect 46770 -148660 47570 -148650
rect 46770 -148690 46780 -148660
rect 47560 -148690 47570 -148660
rect 46770 -148700 47570 -148690
rect 48270 -148660 49070 -148650
rect 48270 -148690 48280 -148660
rect 49060 -148690 49070 -148660
rect 48270 -148700 49070 -148690
rect 49770 -148660 50570 -148650
rect 49770 -148690 49780 -148660
rect 50560 -148690 50570 -148660
rect 49770 -148700 50570 -148690
rect 51270 -148660 52070 -148650
rect 51270 -148690 51280 -148660
rect 52060 -148690 52070 -148660
rect 51270 -148700 52070 -148690
rect 52770 -148660 53570 -148650
rect 52770 -148690 52780 -148660
rect 53560 -148690 53570 -148660
rect 52770 -148700 53570 -148690
rect 54270 -148660 55070 -148650
rect 54270 -148690 54280 -148660
rect 55060 -148690 55070 -148660
rect 54270 -148700 55070 -148690
rect 55770 -148660 56570 -148650
rect 55770 -148690 55780 -148660
rect 56560 -148690 56570 -148660
rect 55770 -148700 56570 -148690
rect 57270 -148660 58070 -148650
rect 57270 -148690 57280 -148660
rect 58060 -148690 58070 -148660
rect 57270 -148700 58070 -148690
rect 58770 -148660 59570 -148650
rect 58770 -148690 58780 -148660
rect 59560 -148690 59570 -148660
rect 58770 -148700 59570 -148690
rect 60270 -148660 61070 -148650
rect 60270 -148690 60280 -148660
rect 61060 -148690 61070 -148660
rect 60270 -148700 61070 -148690
rect 61770 -148660 62570 -148650
rect 61770 -148690 61780 -148660
rect 62560 -148690 62570 -148660
rect 61770 -148700 62570 -148690
rect 63270 -148660 64070 -148650
rect 63270 -148690 63280 -148660
rect 64060 -148690 64070 -148660
rect 63270 -148700 64070 -148690
rect 64770 -148660 65570 -148650
rect 64770 -148690 64780 -148660
rect 65560 -148690 65570 -148660
rect 64770 -148700 65570 -148690
rect 66270 -148660 67070 -148650
rect 66270 -148690 66280 -148660
rect 67060 -148690 67070 -148660
rect 66270 -148700 67070 -148690
rect 67770 -148660 68570 -148650
rect 67770 -148690 67780 -148660
rect 68560 -148690 68570 -148660
rect 67770 -148700 68570 -148690
rect 69270 -148660 70070 -148650
rect 69270 -148690 69280 -148660
rect 70060 -148690 70070 -148660
rect 69270 -148700 70070 -148690
rect 70770 -148660 71570 -148650
rect 70770 -148690 70780 -148660
rect 71560 -148690 71570 -148660
rect 70770 -148700 71570 -148690
rect 72270 -148660 73070 -148650
rect 72270 -148690 72280 -148660
rect 73060 -148690 73070 -148660
rect 72270 -148700 73070 -148690
rect 73770 -148660 74570 -148650
rect 73770 -148690 73780 -148660
rect 74560 -148690 74570 -148660
rect 73770 -148700 74570 -148690
rect 75270 -148660 76070 -148650
rect 75270 -148690 75280 -148660
rect 76060 -148690 76070 -148660
rect 75270 -148700 76070 -148690
rect 76770 -148660 77570 -148650
rect 76770 -148690 76780 -148660
rect 77560 -148690 77570 -148660
rect 76770 -148700 77570 -148690
rect 78270 -148660 79070 -148650
rect 78270 -148690 78280 -148660
rect 79060 -148690 79070 -148660
rect 78270 -148700 79070 -148690
rect 79770 -148660 80570 -148650
rect 79770 -148690 79780 -148660
rect 80560 -148690 80570 -148660
rect 79770 -148700 80570 -148690
rect 81270 -148660 82070 -148650
rect 81270 -148690 81280 -148660
rect 82060 -148690 82070 -148660
rect 81270 -148700 82070 -148690
rect 82770 -148660 83570 -148650
rect 82770 -148690 82780 -148660
rect 83560 -148690 83570 -148660
rect 82770 -148700 83570 -148690
rect 84270 -148660 85070 -148650
rect 84270 -148690 84280 -148660
rect 85060 -148690 85070 -148660
rect 84270 -148700 85070 -148690
rect 85770 -148660 86570 -148650
rect 85770 -148690 85780 -148660
rect 86560 -148690 86570 -148660
rect 85770 -148700 86570 -148690
rect 87270 -148660 88070 -148650
rect 87270 -148690 87280 -148660
rect 88060 -148690 88070 -148660
rect 87270 -148700 88070 -148690
rect 88770 -148660 89570 -148650
rect 88770 -148690 88780 -148660
rect 89560 -148690 89570 -148660
rect 88770 -148700 89570 -148690
rect 90270 -148660 91070 -148650
rect 90270 -148690 90280 -148660
rect 91060 -148690 91070 -148660
rect 90270 -148700 91070 -148690
rect 91770 -148660 92570 -148650
rect 91770 -148690 91780 -148660
rect 92560 -148690 92570 -148660
rect 91770 -148700 92570 -148690
rect 93270 -148660 94070 -148650
rect 93270 -148690 93280 -148660
rect 94060 -148690 94070 -148660
rect 93270 -148700 94070 -148690
rect 94770 -148660 95570 -148650
rect 94770 -148690 94780 -148660
rect 95560 -148690 95570 -148660
rect 94770 -148700 95570 -148690
rect 96270 -148660 97070 -148650
rect 96270 -148690 96280 -148660
rect 97060 -148690 97070 -148660
rect 96270 -148700 97070 -148690
rect 97770 -148660 98570 -148650
rect 97770 -148690 97780 -148660
rect 98560 -148690 98570 -148660
rect 97770 -148700 98570 -148690
rect 99270 -148660 100070 -148650
rect 99270 -148690 99280 -148660
rect 100060 -148690 100070 -148660
rect 99270 -148700 100070 -148690
rect 100770 -148660 101570 -148650
rect 100770 -148690 100780 -148660
rect 101560 -148690 101570 -148660
rect 100770 -148700 101570 -148690
rect 102270 -148660 103070 -148650
rect 102270 -148690 102280 -148660
rect 103060 -148690 103070 -148660
rect 102270 -148700 103070 -148690
rect 103770 -148660 104570 -148650
rect 103770 -148690 103780 -148660
rect 104560 -148690 104570 -148660
rect 103770 -148700 104570 -148690
rect 105270 -148660 106070 -148650
rect 105270 -148690 105280 -148660
rect 106060 -148690 106070 -148660
rect 105270 -148700 106070 -148690
rect 106770 -148660 107570 -148650
rect 106770 -148690 106780 -148660
rect 107560 -148690 107570 -148660
rect 106770 -148700 107570 -148690
rect 108270 -148660 109070 -148650
rect 108270 -148690 108280 -148660
rect 109060 -148690 109070 -148660
rect 108270 -148700 109070 -148690
rect 109770 -148660 110570 -148650
rect 109770 -148690 109780 -148660
rect 110560 -148690 110570 -148660
rect 109770 -148700 110570 -148690
rect 111270 -148660 112070 -148650
rect 111270 -148690 111280 -148660
rect 112060 -148690 112070 -148660
rect 111270 -148700 112070 -148690
rect 112770 -148660 113570 -148650
rect 112770 -148690 112780 -148660
rect 113560 -148690 113570 -148660
rect 112770 -148700 113570 -148690
rect 114270 -148660 115070 -148650
rect 114270 -148690 114280 -148660
rect 115060 -148690 115070 -148660
rect 114270 -148700 115070 -148690
rect 115770 -148660 116570 -148650
rect 115770 -148690 115780 -148660
rect 116560 -148690 116570 -148660
rect 115770 -148700 116570 -148690
rect 117270 -148660 118070 -148650
rect 117270 -148690 117280 -148660
rect 118060 -148690 118070 -148660
rect 117270 -148700 118070 -148690
rect 118770 -148660 119570 -148650
rect 118770 -148690 118780 -148660
rect 119560 -148690 119570 -148660
rect 118770 -148700 119570 -148690
rect 120270 -148660 121070 -148650
rect 120270 -148690 120280 -148660
rect 121060 -148690 121070 -148660
rect 120270 -148700 121070 -148690
rect 121770 -148660 122570 -148650
rect 121770 -148690 121780 -148660
rect 122560 -148690 122570 -148660
rect 121770 -148700 122570 -148690
rect 123270 -148660 124070 -148650
rect 123270 -148690 123280 -148660
rect 124060 -148690 124070 -148660
rect 123270 -148700 124070 -148690
rect 124770 -148660 125570 -148650
rect 124770 -148690 124780 -148660
rect 125560 -148690 125570 -148660
rect 124770 -148700 125570 -148690
rect 126270 -148660 127070 -148650
rect 126270 -148690 126280 -148660
rect 127060 -148690 127070 -148660
rect 126270 -148700 127070 -148690
rect 127770 -148660 128570 -148650
rect 127770 -148690 127780 -148660
rect 128560 -148690 128570 -148660
rect 127770 -148700 128570 -148690
rect 129270 -148660 130070 -148650
rect 129270 -148690 129280 -148660
rect 130060 -148690 130070 -148660
rect 129270 -148700 130070 -148690
rect 130770 -148660 131570 -148650
rect 130770 -148690 130780 -148660
rect 131560 -148690 131570 -148660
rect 130770 -148700 131570 -148690
rect 132270 -148660 133070 -148650
rect 132270 -148690 132280 -148660
rect 133060 -148690 133070 -148660
rect 132270 -148700 133070 -148690
rect 133770 -148660 134570 -148650
rect 133770 -148690 133780 -148660
rect 134560 -148690 134570 -148660
rect 133770 -148700 134570 -148690
rect 135270 -148660 136070 -148650
rect 135270 -148690 135280 -148660
rect 136060 -148690 136070 -148660
rect 135270 -148700 136070 -148690
rect 136770 -148660 137570 -148650
rect 136770 -148690 136780 -148660
rect 137560 -148690 137570 -148660
rect 136770 -148700 137570 -148690
rect 138270 -148660 139070 -148650
rect 138270 -148690 138280 -148660
rect 139060 -148690 139070 -148660
rect 138270 -148700 139070 -148690
rect 139770 -148660 140570 -148650
rect 139770 -148690 139780 -148660
rect 140560 -148690 140570 -148660
rect 139770 -148700 140570 -148690
rect 141270 -148660 142070 -148650
rect 141270 -148690 141280 -148660
rect 142060 -148690 142070 -148660
rect 141270 -148700 142070 -148690
rect 142770 -148660 143570 -148650
rect 142770 -148690 142780 -148660
rect 143560 -148690 143570 -148660
rect 142770 -148700 143570 -148690
rect 144270 -148660 145070 -148650
rect 144270 -148690 144280 -148660
rect 145060 -148690 145070 -148660
rect 144270 -148700 145070 -148690
rect 145770 -148660 146570 -148650
rect 145770 -148690 145780 -148660
rect 146560 -148690 146570 -148660
rect 145770 -148700 146570 -148690
rect 147270 -148660 148070 -148650
rect 147270 -148690 147280 -148660
rect 148060 -148690 148070 -148660
rect 147270 -148700 148070 -148690
rect 148770 -148660 149570 -148650
rect 148770 -148690 148780 -148660
rect 149560 -148690 149570 -148660
rect 148770 -148700 149570 -148690
rect 270 -148915 1070 -148900
rect 270 -148935 280 -148915
rect 1060 -148935 1070 -148915
rect 270 -148940 1070 -148935
rect 1770 -148915 2570 -148900
rect 1770 -148935 1780 -148915
rect 2560 -148935 2570 -148915
rect 1770 -148940 2570 -148935
rect 3270 -148915 4070 -148900
rect 3270 -148935 3280 -148915
rect 4060 -148935 4070 -148915
rect 3270 -148940 4070 -148935
rect 4770 -148915 5570 -148900
rect 4770 -148935 4780 -148915
rect 5560 -148935 5570 -148915
rect 4770 -148940 5570 -148935
rect 6270 -148915 7070 -148900
rect 6270 -148935 6280 -148915
rect 7060 -148935 7070 -148915
rect 6270 -148940 7070 -148935
rect 7770 -148915 8570 -148900
rect 7770 -148935 7780 -148915
rect 8560 -148935 8570 -148915
rect 7770 -148940 8570 -148935
rect 9270 -148915 10070 -148900
rect 9270 -148935 9280 -148915
rect 10060 -148935 10070 -148915
rect 9270 -148940 10070 -148935
rect 10770 -148915 11570 -148900
rect 10770 -148935 10780 -148915
rect 11560 -148935 11570 -148915
rect 10770 -148940 11570 -148935
rect 12270 -148915 13070 -148900
rect 12270 -148935 12280 -148915
rect 13060 -148935 13070 -148915
rect 12270 -148940 13070 -148935
rect 13770 -148915 14570 -148900
rect 13770 -148935 13780 -148915
rect 14560 -148935 14570 -148915
rect 13770 -148940 14570 -148935
rect 15270 -148915 16070 -148900
rect 15270 -148935 15280 -148915
rect 16060 -148935 16070 -148915
rect 15270 -148940 16070 -148935
rect 16770 -148915 17570 -148900
rect 16770 -148935 16780 -148915
rect 17560 -148935 17570 -148915
rect 16770 -148940 17570 -148935
rect 18270 -148915 19070 -148900
rect 18270 -148935 18280 -148915
rect 19060 -148935 19070 -148915
rect 18270 -148940 19070 -148935
rect 19770 -148915 20570 -148900
rect 19770 -148935 19780 -148915
rect 20560 -148935 20570 -148915
rect 19770 -148940 20570 -148935
rect 21270 -148915 22070 -148900
rect 21270 -148935 21280 -148915
rect 22060 -148935 22070 -148915
rect 21270 -148940 22070 -148935
rect 22770 -148915 23570 -148900
rect 22770 -148935 22780 -148915
rect 23560 -148935 23570 -148915
rect 22770 -148940 23570 -148935
rect 24270 -148915 25070 -148900
rect 24270 -148935 24280 -148915
rect 25060 -148935 25070 -148915
rect 24270 -148940 25070 -148935
rect 25770 -148915 26570 -148900
rect 25770 -148935 25780 -148915
rect 26560 -148935 26570 -148915
rect 25770 -148940 26570 -148935
rect 27270 -148915 28070 -148900
rect 27270 -148935 27280 -148915
rect 28060 -148935 28070 -148915
rect 27270 -148940 28070 -148935
rect 28770 -148915 29570 -148900
rect 28770 -148935 28780 -148915
rect 29560 -148935 29570 -148915
rect 28770 -148940 29570 -148935
rect 30270 -148915 31070 -148900
rect 30270 -148935 30280 -148915
rect 31060 -148935 31070 -148915
rect 30270 -148940 31070 -148935
rect 31770 -148915 32570 -148900
rect 31770 -148935 31780 -148915
rect 32560 -148935 32570 -148915
rect 31770 -148940 32570 -148935
rect 33270 -148915 34070 -148900
rect 33270 -148935 33280 -148915
rect 34060 -148935 34070 -148915
rect 33270 -148940 34070 -148935
rect 34770 -148915 35570 -148900
rect 34770 -148935 34780 -148915
rect 35560 -148935 35570 -148915
rect 34770 -148940 35570 -148935
rect 36270 -148915 37070 -148900
rect 36270 -148935 36280 -148915
rect 37060 -148935 37070 -148915
rect 36270 -148940 37070 -148935
rect 37770 -148915 38570 -148900
rect 37770 -148935 37780 -148915
rect 38560 -148935 38570 -148915
rect 37770 -148940 38570 -148935
rect 39270 -148915 40070 -148900
rect 39270 -148935 39280 -148915
rect 40060 -148935 40070 -148915
rect 39270 -148940 40070 -148935
rect 40770 -148915 41570 -148900
rect 40770 -148935 40780 -148915
rect 41560 -148935 41570 -148915
rect 40770 -148940 41570 -148935
rect 42270 -148915 43070 -148900
rect 42270 -148935 42280 -148915
rect 43060 -148935 43070 -148915
rect 42270 -148940 43070 -148935
rect 43770 -148915 44570 -148900
rect 43770 -148935 43780 -148915
rect 44560 -148935 44570 -148915
rect 43770 -148940 44570 -148935
rect 45270 -148915 46070 -148900
rect 45270 -148935 45280 -148915
rect 46060 -148935 46070 -148915
rect 45270 -148940 46070 -148935
rect 46770 -148915 47570 -148900
rect 46770 -148935 46780 -148915
rect 47560 -148935 47570 -148915
rect 46770 -148940 47570 -148935
rect 48270 -148915 49070 -148900
rect 48270 -148935 48280 -148915
rect 49060 -148935 49070 -148915
rect 48270 -148940 49070 -148935
rect 49770 -148915 50570 -148900
rect 49770 -148935 49780 -148915
rect 50560 -148935 50570 -148915
rect 49770 -148940 50570 -148935
rect 51270 -148915 52070 -148900
rect 51270 -148935 51280 -148915
rect 52060 -148935 52070 -148915
rect 51270 -148940 52070 -148935
rect 52770 -148915 53570 -148900
rect 52770 -148935 52780 -148915
rect 53560 -148935 53570 -148915
rect 52770 -148940 53570 -148935
rect 54270 -148915 55070 -148900
rect 54270 -148935 54280 -148915
rect 55060 -148935 55070 -148915
rect 54270 -148940 55070 -148935
rect 55770 -148915 56570 -148900
rect 55770 -148935 55780 -148915
rect 56560 -148935 56570 -148915
rect 55770 -148940 56570 -148935
rect 57270 -148915 58070 -148900
rect 57270 -148935 57280 -148915
rect 58060 -148935 58070 -148915
rect 57270 -148940 58070 -148935
rect 58770 -148915 59570 -148900
rect 58770 -148935 58780 -148915
rect 59560 -148935 59570 -148915
rect 58770 -148940 59570 -148935
rect 60270 -148915 61070 -148900
rect 60270 -148935 60280 -148915
rect 61060 -148935 61070 -148915
rect 60270 -148940 61070 -148935
rect 61770 -148915 62570 -148900
rect 61770 -148935 61780 -148915
rect 62560 -148935 62570 -148915
rect 61770 -148940 62570 -148935
rect 63270 -148915 64070 -148900
rect 63270 -148935 63280 -148915
rect 64060 -148935 64070 -148915
rect 63270 -148940 64070 -148935
rect 64770 -148915 65570 -148900
rect 64770 -148935 64780 -148915
rect 65560 -148935 65570 -148915
rect 64770 -148940 65570 -148935
rect 66270 -148915 67070 -148900
rect 66270 -148935 66280 -148915
rect 67060 -148935 67070 -148915
rect 66270 -148940 67070 -148935
rect 67770 -148915 68570 -148900
rect 67770 -148935 67780 -148915
rect 68560 -148935 68570 -148915
rect 67770 -148940 68570 -148935
rect 69270 -148915 70070 -148900
rect 69270 -148935 69280 -148915
rect 70060 -148935 70070 -148915
rect 69270 -148940 70070 -148935
rect 70770 -148915 71570 -148900
rect 70770 -148935 70780 -148915
rect 71560 -148935 71570 -148915
rect 70770 -148940 71570 -148935
rect 72270 -148915 73070 -148900
rect 72270 -148935 72280 -148915
rect 73060 -148935 73070 -148915
rect 72270 -148940 73070 -148935
rect 73770 -148915 74570 -148900
rect 73770 -148935 73780 -148915
rect 74560 -148935 74570 -148915
rect 73770 -148940 74570 -148935
rect 75270 -148915 76070 -148900
rect 75270 -148935 75280 -148915
rect 76060 -148935 76070 -148915
rect 75270 -148940 76070 -148935
rect 76770 -148915 77570 -148900
rect 76770 -148935 76780 -148915
rect 77560 -148935 77570 -148915
rect 76770 -148940 77570 -148935
rect 78270 -148915 79070 -148900
rect 78270 -148935 78280 -148915
rect 79060 -148935 79070 -148915
rect 78270 -148940 79070 -148935
rect 79770 -148915 80570 -148900
rect 79770 -148935 79780 -148915
rect 80560 -148935 80570 -148915
rect 79770 -148940 80570 -148935
rect 81270 -148915 82070 -148900
rect 81270 -148935 81280 -148915
rect 82060 -148935 82070 -148915
rect 81270 -148940 82070 -148935
rect 82770 -148915 83570 -148900
rect 82770 -148935 82780 -148915
rect 83560 -148935 83570 -148915
rect 82770 -148940 83570 -148935
rect 84270 -148915 85070 -148900
rect 84270 -148935 84280 -148915
rect 85060 -148935 85070 -148915
rect 84270 -148940 85070 -148935
rect 85770 -148915 86570 -148900
rect 85770 -148935 85780 -148915
rect 86560 -148935 86570 -148915
rect 85770 -148940 86570 -148935
rect 87270 -148915 88070 -148900
rect 87270 -148935 87280 -148915
rect 88060 -148935 88070 -148915
rect 87270 -148940 88070 -148935
rect 88770 -148915 89570 -148900
rect 88770 -148935 88780 -148915
rect 89560 -148935 89570 -148915
rect 88770 -148940 89570 -148935
rect 90270 -148915 91070 -148900
rect 90270 -148935 90280 -148915
rect 91060 -148935 91070 -148915
rect 90270 -148940 91070 -148935
rect 91770 -148915 92570 -148900
rect 91770 -148935 91780 -148915
rect 92560 -148935 92570 -148915
rect 91770 -148940 92570 -148935
rect 93270 -148915 94070 -148900
rect 93270 -148935 93280 -148915
rect 94060 -148935 94070 -148915
rect 93270 -148940 94070 -148935
rect 94770 -148915 95570 -148900
rect 94770 -148935 94780 -148915
rect 95560 -148935 95570 -148915
rect 94770 -148940 95570 -148935
rect 96270 -148915 97070 -148900
rect 96270 -148935 96280 -148915
rect 97060 -148935 97070 -148915
rect 96270 -148940 97070 -148935
rect 97770 -148915 98570 -148900
rect 97770 -148935 97780 -148915
rect 98560 -148935 98570 -148915
rect 97770 -148940 98570 -148935
rect 99270 -148915 100070 -148900
rect 99270 -148935 99280 -148915
rect 100060 -148935 100070 -148915
rect 99270 -148940 100070 -148935
rect 100770 -148915 101570 -148900
rect 100770 -148935 100780 -148915
rect 101560 -148935 101570 -148915
rect 100770 -148940 101570 -148935
rect 102270 -148915 103070 -148900
rect 102270 -148935 102280 -148915
rect 103060 -148935 103070 -148915
rect 102270 -148940 103070 -148935
rect 103770 -148915 104570 -148900
rect 103770 -148935 103780 -148915
rect 104560 -148935 104570 -148915
rect 103770 -148940 104570 -148935
rect 105270 -148915 106070 -148900
rect 105270 -148935 105280 -148915
rect 106060 -148935 106070 -148915
rect 105270 -148940 106070 -148935
rect 106770 -148915 107570 -148900
rect 106770 -148935 106780 -148915
rect 107560 -148935 107570 -148915
rect 106770 -148940 107570 -148935
rect 108270 -148915 109070 -148900
rect 108270 -148935 108280 -148915
rect 109060 -148935 109070 -148915
rect 108270 -148940 109070 -148935
rect 109770 -148915 110570 -148900
rect 109770 -148935 109780 -148915
rect 110560 -148935 110570 -148915
rect 109770 -148940 110570 -148935
rect 111270 -148915 112070 -148900
rect 111270 -148935 111280 -148915
rect 112060 -148935 112070 -148915
rect 111270 -148940 112070 -148935
rect 112770 -148915 113570 -148900
rect 112770 -148935 112780 -148915
rect 113560 -148935 113570 -148915
rect 112770 -148940 113570 -148935
rect 114270 -148915 115070 -148900
rect 114270 -148935 114280 -148915
rect 115060 -148935 115070 -148915
rect 114270 -148940 115070 -148935
rect 115770 -148915 116570 -148900
rect 115770 -148935 115780 -148915
rect 116560 -148935 116570 -148915
rect 115770 -148940 116570 -148935
rect 117270 -148915 118070 -148900
rect 117270 -148935 117280 -148915
rect 118060 -148935 118070 -148915
rect 117270 -148940 118070 -148935
rect 118770 -148915 119570 -148900
rect 118770 -148935 118780 -148915
rect 119560 -148935 119570 -148915
rect 118770 -148940 119570 -148935
rect 120270 -148915 121070 -148900
rect 120270 -148935 120280 -148915
rect 121060 -148935 121070 -148915
rect 120270 -148940 121070 -148935
rect 121770 -148915 122570 -148900
rect 121770 -148935 121780 -148915
rect 122560 -148935 122570 -148915
rect 121770 -148940 122570 -148935
rect 123270 -148915 124070 -148900
rect 123270 -148935 123280 -148915
rect 124060 -148935 124070 -148915
rect 123270 -148940 124070 -148935
rect 124770 -148915 125570 -148900
rect 124770 -148935 124780 -148915
rect 125560 -148935 125570 -148915
rect 124770 -148940 125570 -148935
rect 126270 -148915 127070 -148900
rect 126270 -148935 126280 -148915
rect 127060 -148935 127070 -148915
rect 126270 -148940 127070 -148935
rect 127770 -148915 128570 -148900
rect 127770 -148935 127780 -148915
rect 128560 -148935 128570 -148915
rect 127770 -148940 128570 -148935
rect 129270 -148915 130070 -148900
rect 129270 -148935 129280 -148915
rect 130060 -148935 130070 -148915
rect 129270 -148940 130070 -148935
rect 130770 -148915 131570 -148900
rect 130770 -148935 130780 -148915
rect 131560 -148935 131570 -148915
rect 130770 -148940 131570 -148935
rect 132270 -148915 133070 -148900
rect 132270 -148935 132280 -148915
rect 133060 -148935 133070 -148915
rect 132270 -148940 133070 -148935
rect 133770 -148915 134570 -148900
rect 133770 -148935 133780 -148915
rect 134560 -148935 134570 -148915
rect 133770 -148940 134570 -148935
rect 135270 -148915 136070 -148900
rect 135270 -148935 135280 -148915
rect 136060 -148935 136070 -148915
rect 135270 -148940 136070 -148935
rect 136770 -148915 137570 -148900
rect 136770 -148935 136780 -148915
rect 137560 -148935 137570 -148915
rect 136770 -148940 137570 -148935
rect 138270 -148915 139070 -148900
rect 138270 -148935 138280 -148915
rect 139060 -148935 139070 -148915
rect 138270 -148940 139070 -148935
rect 139770 -148915 140570 -148900
rect 139770 -148935 139780 -148915
rect 140560 -148935 140570 -148915
rect 139770 -148940 140570 -148935
rect 141270 -148915 142070 -148900
rect 141270 -148935 141280 -148915
rect 142060 -148935 142070 -148915
rect 141270 -148940 142070 -148935
rect 142770 -148915 143570 -148900
rect 142770 -148935 142780 -148915
rect 143560 -148935 143570 -148915
rect 142770 -148940 143570 -148935
rect 144270 -148915 145070 -148900
rect 144270 -148935 144280 -148915
rect 145060 -148935 145070 -148915
rect 144270 -148940 145070 -148935
rect 145770 -148915 146570 -148900
rect 145770 -148935 145780 -148915
rect 146560 -148935 146570 -148915
rect 145770 -148940 146570 -148935
rect 147270 -148915 148070 -148900
rect 147270 -148935 147280 -148915
rect 148060 -148935 148070 -148915
rect 147270 -148940 148070 -148935
rect 148770 -148915 149570 -148900
rect 148770 -148935 148780 -148915
rect 149560 -148935 149570 -148915
rect 148770 -148940 149570 -148935
<< ndiffc >>
rect 280 -148690 1060 -148660
rect 1780 -148690 2560 -148660
rect 3280 -148690 4060 -148660
rect 4780 -148690 5560 -148660
rect 6280 -148690 7060 -148660
rect 7780 -148690 8560 -148660
rect 9280 -148690 10060 -148660
rect 10780 -148690 11560 -148660
rect 12280 -148690 13060 -148660
rect 13780 -148690 14560 -148660
rect 15280 -148690 16060 -148660
rect 16780 -148690 17560 -148660
rect 18280 -148690 19060 -148660
rect 19780 -148690 20560 -148660
rect 21280 -148690 22060 -148660
rect 22780 -148690 23560 -148660
rect 24280 -148690 25060 -148660
rect 25780 -148690 26560 -148660
rect 27280 -148690 28060 -148660
rect 28780 -148690 29560 -148660
rect 30280 -148690 31060 -148660
rect 31780 -148690 32560 -148660
rect 33280 -148690 34060 -148660
rect 34780 -148690 35560 -148660
rect 36280 -148690 37060 -148660
rect 37780 -148690 38560 -148660
rect 39280 -148690 40060 -148660
rect 40780 -148690 41560 -148660
rect 42280 -148690 43060 -148660
rect 43780 -148690 44560 -148660
rect 45280 -148690 46060 -148660
rect 46780 -148690 47560 -148660
rect 48280 -148690 49060 -148660
rect 49780 -148690 50560 -148660
rect 51280 -148690 52060 -148660
rect 52780 -148690 53560 -148660
rect 54280 -148690 55060 -148660
rect 55780 -148690 56560 -148660
rect 57280 -148690 58060 -148660
rect 58780 -148690 59560 -148660
rect 60280 -148690 61060 -148660
rect 61780 -148690 62560 -148660
rect 63280 -148690 64060 -148660
rect 64780 -148690 65560 -148660
rect 66280 -148690 67060 -148660
rect 67780 -148690 68560 -148660
rect 69280 -148690 70060 -148660
rect 70780 -148690 71560 -148660
rect 72280 -148690 73060 -148660
rect 73780 -148690 74560 -148660
rect 75280 -148690 76060 -148660
rect 76780 -148690 77560 -148660
rect 78280 -148690 79060 -148660
rect 79780 -148690 80560 -148660
rect 81280 -148690 82060 -148660
rect 82780 -148690 83560 -148660
rect 84280 -148690 85060 -148660
rect 85780 -148690 86560 -148660
rect 87280 -148690 88060 -148660
rect 88780 -148690 89560 -148660
rect 90280 -148690 91060 -148660
rect 91780 -148690 92560 -148660
rect 93280 -148690 94060 -148660
rect 94780 -148690 95560 -148660
rect 96280 -148690 97060 -148660
rect 97780 -148690 98560 -148660
rect 99280 -148690 100060 -148660
rect 100780 -148690 101560 -148660
rect 102280 -148690 103060 -148660
rect 103780 -148690 104560 -148660
rect 105280 -148690 106060 -148660
rect 106780 -148690 107560 -148660
rect 108280 -148690 109060 -148660
rect 109780 -148690 110560 -148660
rect 111280 -148690 112060 -148660
rect 112780 -148690 113560 -148660
rect 114280 -148690 115060 -148660
rect 115780 -148690 116560 -148660
rect 117280 -148690 118060 -148660
rect 118780 -148690 119560 -148660
rect 120280 -148690 121060 -148660
rect 121780 -148690 122560 -148660
rect 123280 -148690 124060 -148660
rect 124780 -148690 125560 -148660
rect 126280 -148690 127060 -148660
rect 127780 -148690 128560 -148660
rect 129280 -148690 130060 -148660
rect 130780 -148690 131560 -148660
rect 132280 -148690 133060 -148660
rect 133780 -148690 134560 -148660
rect 135280 -148690 136060 -148660
rect 136780 -148690 137560 -148660
rect 138280 -148690 139060 -148660
rect 139780 -148690 140560 -148660
rect 141280 -148690 142060 -148660
rect 142780 -148690 143560 -148660
rect 144280 -148690 145060 -148660
rect 145780 -148690 146560 -148660
rect 147280 -148690 148060 -148660
rect 148780 -148690 149560 -148660
rect 280 -148935 1060 -148915
rect 1780 -148935 2560 -148915
rect 3280 -148935 4060 -148915
rect 4780 -148935 5560 -148915
rect 6280 -148935 7060 -148915
rect 7780 -148935 8560 -148915
rect 9280 -148935 10060 -148915
rect 10780 -148935 11560 -148915
rect 12280 -148935 13060 -148915
rect 13780 -148935 14560 -148915
rect 15280 -148935 16060 -148915
rect 16780 -148935 17560 -148915
rect 18280 -148935 19060 -148915
rect 19780 -148935 20560 -148915
rect 21280 -148935 22060 -148915
rect 22780 -148935 23560 -148915
rect 24280 -148935 25060 -148915
rect 25780 -148935 26560 -148915
rect 27280 -148935 28060 -148915
rect 28780 -148935 29560 -148915
rect 30280 -148935 31060 -148915
rect 31780 -148935 32560 -148915
rect 33280 -148935 34060 -148915
rect 34780 -148935 35560 -148915
rect 36280 -148935 37060 -148915
rect 37780 -148935 38560 -148915
rect 39280 -148935 40060 -148915
rect 40780 -148935 41560 -148915
rect 42280 -148935 43060 -148915
rect 43780 -148935 44560 -148915
rect 45280 -148935 46060 -148915
rect 46780 -148935 47560 -148915
rect 48280 -148935 49060 -148915
rect 49780 -148935 50560 -148915
rect 51280 -148935 52060 -148915
rect 52780 -148935 53560 -148915
rect 54280 -148935 55060 -148915
rect 55780 -148935 56560 -148915
rect 57280 -148935 58060 -148915
rect 58780 -148935 59560 -148915
rect 60280 -148935 61060 -148915
rect 61780 -148935 62560 -148915
rect 63280 -148935 64060 -148915
rect 64780 -148935 65560 -148915
rect 66280 -148935 67060 -148915
rect 67780 -148935 68560 -148915
rect 69280 -148935 70060 -148915
rect 70780 -148935 71560 -148915
rect 72280 -148935 73060 -148915
rect 73780 -148935 74560 -148915
rect 75280 -148935 76060 -148915
rect 76780 -148935 77560 -148915
rect 78280 -148935 79060 -148915
rect 79780 -148935 80560 -148915
rect 81280 -148935 82060 -148915
rect 82780 -148935 83560 -148915
rect 84280 -148935 85060 -148915
rect 85780 -148935 86560 -148915
rect 87280 -148935 88060 -148915
rect 88780 -148935 89560 -148915
rect 90280 -148935 91060 -148915
rect 91780 -148935 92560 -148915
rect 93280 -148935 94060 -148915
rect 94780 -148935 95560 -148915
rect 96280 -148935 97060 -148915
rect 97780 -148935 98560 -148915
rect 99280 -148935 100060 -148915
rect 100780 -148935 101560 -148915
rect 102280 -148935 103060 -148915
rect 103780 -148935 104560 -148915
rect 105280 -148935 106060 -148915
rect 106780 -148935 107560 -148915
rect 108280 -148935 109060 -148915
rect 109780 -148935 110560 -148915
rect 111280 -148935 112060 -148915
rect 112780 -148935 113560 -148915
rect 114280 -148935 115060 -148915
rect 115780 -148935 116560 -148915
rect 117280 -148935 118060 -148915
rect 118780 -148935 119560 -148915
rect 120280 -148935 121060 -148915
rect 121780 -148935 122560 -148915
rect 123280 -148935 124060 -148915
rect 124780 -148935 125560 -148915
rect 126280 -148935 127060 -148915
rect 127780 -148935 128560 -148915
rect 129280 -148935 130060 -148915
rect 130780 -148935 131560 -148915
rect 132280 -148935 133060 -148915
rect 133780 -148935 134560 -148915
rect 135280 -148935 136060 -148915
rect 136780 -148935 137560 -148915
rect 138280 -148935 139060 -148915
rect 139780 -148935 140560 -148915
rect 141280 -148935 142060 -148915
rect 142780 -148935 143560 -148915
rect 144280 -148935 145060 -148915
rect 145780 -148935 146560 -148915
rect 147280 -148935 148060 -148915
rect 148780 -148935 149560 -148915
<< poly >>
rect 255 -148745 270 -148700
rect 110 -148750 270 -148745
rect 110 -148850 120 -148750
rect 210 -148850 270 -148750
rect 110 -148855 270 -148850
rect 255 -148900 270 -148855
rect 1070 -148900 1085 -148700
rect 1755 -148745 1770 -148700
rect 1610 -148750 1770 -148745
rect 1610 -148850 1620 -148750
rect 1710 -148850 1770 -148750
rect 1610 -148855 1770 -148850
rect 1755 -148900 1770 -148855
rect 2570 -148900 2585 -148700
rect 3255 -148745 3270 -148700
rect 3110 -148750 3270 -148745
rect 3110 -148850 3120 -148750
rect 3210 -148850 3270 -148750
rect 3110 -148855 3270 -148850
rect 3255 -148900 3270 -148855
rect 4070 -148900 4085 -148700
rect 4755 -148745 4770 -148700
rect 4610 -148750 4770 -148745
rect 4610 -148850 4620 -148750
rect 4710 -148850 4770 -148750
rect 4610 -148855 4770 -148850
rect 4755 -148900 4770 -148855
rect 5570 -148900 5585 -148700
rect 6255 -148745 6270 -148700
rect 6110 -148750 6270 -148745
rect 6110 -148850 6120 -148750
rect 6210 -148850 6270 -148750
rect 6110 -148855 6270 -148850
rect 6255 -148900 6270 -148855
rect 7070 -148900 7085 -148700
rect 7755 -148745 7770 -148700
rect 7610 -148750 7770 -148745
rect 7610 -148850 7620 -148750
rect 7710 -148850 7770 -148750
rect 7610 -148855 7770 -148850
rect 7755 -148900 7770 -148855
rect 8570 -148900 8585 -148700
rect 9255 -148745 9270 -148700
rect 9110 -148750 9270 -148745
rect 9110 -148850 9120 -148750
rect 9210 -148850 9270 -148750
rect 9110 -148855 9270 -148850
rect 9255 -148900 9270 -148855
rect 10070 -148900 10085 -148700
rect 10755 -148745 10770 -148700
rect 10610 -148750 10770 -148745
rect 10610 -148850 10620 -148750
rect 10710 -148850 10770 -148750
rect 10610 -148855 10770 -148850
rect 10755 -148900 10770 -148855
rect 11570 -148900 11585 -148700
rect 12255 -148745 12270 -148700
rect 12110 -148750 12270 -148745
rect 12110 -148850 12120 -148750
rect 12210 -148850 12270 -148750
rect 12110 -148855 12270 -148850
rect 12255 -148900 12270 -148855
rect 13070 -148900 13085 -148700
rect 13755 -148745 13770 -148700
rect 13610 -148750 13770 -148745
rect 13610 -148850 13620 -148750
rect 13710 -148850 13770 -148750
rect 13610 -148855 13770 -148850
rect 13755 -148900 13770 -148855
rect 14570 -148900 14585 -148700
rect 15255 -148745 15270 -148700
rect 15110 -148750 15270 -148745
rect 15110 -148850 15120 -148750
rect 15210 -148850 15270 -148750
rect 15110 -148855 15270 -148850
rect 15255 -148900 15270 -148855
rect 16070 -148900 16085 -148700
rect 16755 -148745 16770 -148700
rect 16610 -148750 16770 -148745
rect 16610 -148850 16620 -148750
rect 16710 -148850 16770 -148750
rect 16610 -148855 16770 -148850
rect 16755 -148900 16770 -148855
rect 17570 -148900 17585 -148700
rect 18255 -148745 18270 -148700
rect 18110 -148750 18270 -148745
rect 18110 -148850 18120 -148750
rect 18210 -148850 18270 -148750
rect 18110 -148855 18270 -148850
rect 18255 -148900 18270 -148855
rect 19070 -148900 19085 -148700
rect 19755 -148745 19770 -148700
rect 19610 -148750 19770 -148745
rect 19610 -148850 19620 -148750
rect 19710 -148850 19770 -148750
rect 19610 -148855 19770 -148850
rect 19755 -148900 19770 -148855
rect 20570 -148900 20585 -148700
rect 21255 -148745 21270 -148700
rect 21110 -148750 21270 -148745
rect 21110 -148850 21120 -148750
rect 21210 -148850 21270 -148750
rect 21110 -148855 21270 -148850
rect 21255 -148900 21270 -148855
rect 22070 -148900 22085 -148700
rect 22755 -148745 22770 -148700
rect 22610 -148750 22770 -148745
rect 22610 -148850 22620 -148750
rect 22710 -148850 22770 -148750
rect 22610 -148855 22770 -148850
rect 22755 -148900 22770 -148855
rect 23570 -148900 23585 -148700
rect 24255 -148745 24270 -148700
rect 24110 -148750 24270 -148745
rect 24110 -148850 24120 -148750
rect 24210 -148850 24270 -148750
rect 24110 -148855 24270 -148850
rect 24255 -148900 24270 -148855
rect 25070 -148900 25085 -148700
rect 25755 -148745 25770 -148700
rect 25610 -148750 25770 -148745
rect 25610 -148850 25620 -148750
rect 25710 -148850 25770 -148750
rect 25610 -148855 25770 -148850
rect 25755 -148900 25770 -148855
rect 26570 -148900 26585 -148700
rect 27255 -148745 27270 -148700
rect 27110 -148750 27270 -148745
rect 27110 -148850 27120 -148750
rect 27210 -148850 27270 -148750
rect 27110 -148855 27270 -148850
rect 27255 -148900 27270 -148855
rect 28070 -148900 28085 -148700
rect 28755 -148745 28770 -148700
rect 28610 -148750 28770 -148745
rect 28610 -148850 28620 -148750
rect 28710 -148850 28770 -148750
rect 28610 -148855 28770 -148850
rect 28755 -148900 28770 -148855
rect 29570 -148900 29585 -148700
rect 30255 -148745 30270 -148700
rect 30110 -148750 30270 -148745
rect 30110 -148850 30120 -148750
rect 30210 -148850 30270 -148750
rect 30110 -148855 30270 -148850
rect 30255 -148900 30270 -148855
rect 31070 -148900 31085 -148700
rect 31755 -148745 31770 -148700
rect 31610 -148750 31770 -148745
rect 31610 -148850 31620 -148750
rect 31710 -148850 31770 -148750
rect 31610 -148855 31770 -148850
rect 31755 -148900 31770 -148855
rect 32570 -148900 32585 -148700
rect 33255 -148745 33270 -148700
rect 33110 -148750 33270 -148745
rect 33110 -148850 33120 -148750
rect 33210 -148850 33270 -148750
rect 33110 -148855 33270 -148850
rect 33255 -148900 33270 -148855
rect 34070 -148900 34085 -148700
rect 34755 -148745 34770 -148700
rect 34610 -148750 34770 -148745
rect 34610 -148850 34620 -148750
rect 34710 -148850 34770 -148750
rect 34610 -148855 34770 -148850
rect 34755 -148900 34770 -148855
rect 35570 -148900 35585 -148700
rect 36255 -148745 36270 -148700
rect 36110 -148750 36270 -148745
rect 36110 -148850 36120 -148750
rect 36210 -148850 36270 -148750
rect 36110 -148855 36270 -148850
rect 36255 -148900 36270 -148855
rect 37070 -148900 37085 -148700
rect 37755 -148745 37770 -148700
rect 37610 -148750 37770 -148745
rect 37610 -148850 37620 -148750
rect 37710 -148850 37770 -148750
rect 37610 -148855 37770 -148850
rect 37755 -148900 37770 -148855
rect 38570 -148900 38585 -148700
rect 39255 -148745 39270 -148700
rect 39110 -148750 39270 -148745
rect 39110 -148850 39120 -148750
rect 39210 -148850 39270 -148750
rect 39110 -148855 39270 -148850
rect 39255 -148900 39270 -148855
rect 40070 -148900 40085 -148700
rect 40755 -148745 40770 -148700
rect 40610 -148750 40770 -148745
rect 40610 -148850 40620 -148750
rect 40710 -148850 40770 -148750
rect 40610 -148855 40770 -148850
rect 40755 -148900 40770 -148855
rect 41570 -148900 41585 -148700
rect 42255 -148745 42270 -148700
rect 42110 -148750 42270 -148745
rect 42110 -148850 42120 -148750
rect 42210 -148850 42270 -148750
rect 42110 -148855 42270 -148850
rect 42255 -148900 42270 -148855
rect 43070 -148900 43085 -148700
rect 43755 -148745 43770 -148700
rect 43610 -148750 43770 -148745
rect 43610 -148850 43620 -148750
rect 43710 -148850 43770 -148750
rect 43610 -148855 43770 -148850
rect 43755 -148900 43770 -148855
rect 44570 -148900 44585 -148700
rect 45255 -148745 45270 -148700
rect 45110 -148750 45270 -148745
rect 45110 -148850 45120 -148750
rect 45210 -148850 45270 -148750
rect 45110 -148855 45270 -148850
rect 45255 -148900 45270 -148855
rect 46070 -148900 46085 -148700
rect 46755 -148745 46770 -148700
rect 46610 -148750 46770 -148745
rect 46610 -148850 46620 -148750
rect 46710 -148850 46770 -148750
rect 46610 -148855 46770 -148850
rect 46755 -148900 46770 -148855
rect 47570 -148900 47585 -148700
rect 48255 -148745 48270 -148700
rect 48110 -148750 48270 -148745
rect 48110 -148850 48120 -148750
rect 48210 -148850 48270 -148750
rect 48110 -148855 48270 -148850
rect 48255 -148900 48270 -148855
rect 49070 -148900 49085 -148700
rect 49755 -148745 49770 -148700
rect 49610 -148750 49770 -148745
rect 49610 -148850 49620 -148750
rect 49710 -148850 49770 -148750
rect 49610 -148855 49770 -148850
rect 49755 -148900 49770 -148855
rect 50570 -148900 50585 -148700
rect 51255 -148745 51270 -148700
rect 51110 -148750 51270 -148745
rect 51110 -148850 51120 -148750
rect 51210 -148850 51270 -148750
rect 51110 -148855 51270 -148850
rect 51255 -148900 51270 -148855
rect 52070 -148900 52085 -148700
rect 52755 -148745 52770 -148700
rect 52610 -148750 52770 -148745
rect 52610 -148850 52620 -148750
rect 52710 -148850 52770 -148750
rect 52610 -148855 52770 -148850
rect 52755 -148900 52770 -148855
rect 53570 -148900 53585 -148700
rect 54255 -148745 54270 -148700
rect 54110 -148750 54270 -148745
rect 54110 -148850 54120 -148750
rect 54210 -148850 54270 -148750
rect 54110 -148855 54270 -148850
rect 54255 -148900 54270 -148855
rect 55070 -148900 55085 -148700
rect 55755 -148745 55770 -148700
rect 55610 -148750 55770 -148745
rect 55610 -148850 55620 -148750
rect 55710 -148850 55770 -148750
rect 55610 -148855 55770 -148850
rect 55755 -148900 55770 -148855
rect 56570 -148900 56585 -148700
rect 57255 -148745 57270 -148700
rect 57110 -148750 57270 -148745
rect 57110 -148850 57120 -148750
rect 57210 -148850 57270 -148750
rect 57110 -148855 57270 -148850
rect 57255 -148900 57270 -148855
rect 58070 -148900 58085 -148700
rect 58755 -148745 58770 -148700
rect 58610 -148750 58770 -148745
rect 58610 -148850 58620 -148750
rect 58710 -148850 58770 -148750
rect 58610 -148855 58770 -148850
rect 58755 -148900 58770 -148855
rect 59570 -148900 59585 -148700
rect 60255 -148745 60270 -148700
rect 60110 -148750 60270 -148745
rect 60110 -148850 60120 -148750
rect 60210 -148850 60270 -148750
rect 60110 -148855 60270 -148850
rect 60255 -148900 60270 -148855
rect 61070 -148900 61085 -148700
rect 61755 -148745 61770 -148700
rect 61610 -148750 61770 -148745
rect 61610 -148850 61620 -148750
rect 61710 -148850 61770 -148750
rect 61610 -148855 61770 -148850
rect 61755 -148900 61770 -148855
rect 62570 -148900 62585 -148700
rect 63255 -148745 63270 -148700
rect 63110 -148750 63270 -148745
rect 63110 -148850 63120 -148750
rect 63210 -148850 63270 -148750
rect 63110 -148855 63270 -148850
rect 63255 -148900 63270 -148855
rect 64070 -148900 64085 -148700
rect 64755 -148745 64770 -148700
rect 64610 -148750 64770 -148745
rect 64610 -148850 64620 -148750
rect 64710 -148850 64770 -148750
rect 64610 -148855 64770 -148850
rect 64755 -148900 64770 -148855
rect 65570 -148900 65585 -148700
rect 66255 -148745 66270 -148700
rect 66110 -148750 66270 -148745
rect 66110 -148850 66120 -148750
rect 66210 -148850 66270 -148750
rect 66110 -148855 66270 -148850
rect 66255 -148900 66270 -148855
rect 67070 -148900 67085 -148700
rect 67755 -148745 67770 -148700
rect 67610 -148750 67770 -148745
rect 67610 -148850 67620 -148750
rect 67710 -148850 67770 -148750
rect 67610 -148855 67770 -148850
rect 67755 -148900 67770 -148855
rect 68570 -148900 68585 -148700
rect 69255 -148745 69270 -148700
rect 69110 -148750 69270 -148745
rect 69110 -148850 69120 -148750
rect 69210 -148850 69270 -148750
rect 69110 -148855 69270 -148850
rect 69255 -148900 69270 -148855
rect 70070 -148900 70085 -148700
rect 70755 -148745 70770 -148700
rect 70610 -148750 70770 -148745
rect 70610 -148850 70620 -148750
rect 70710 -148850 70770 -148750
rect 70610 -148855 70770 -148850
rect 70755 -148900 70770 -148855
rect 71570 -148900 71585 -148700
rect 72255 -148745 72270 -148700
rect 72110 -148750 72270 -148745
rect 72110 -148850 72120 -148750
rect 72210 -148850 72270 -148750
rect 72110 -148855 72270 -148850
rect 72255 -148900 72270 -148855
rect 73070 -148900 73085 -148700
rect 73755 -148745 73770 -148700
rect 73610 -148750 73770 -148745
rect 73610 -148850 73620 -148750
rect 73710 -148850 73770 -148750
rect 73610 -148855 73770 -148850
rect 73755 -148900 73770 -148855
rect 74570 -148900 74585 -148700
rect 75255 -148745 75270 -148700
rect 75110 -148750 75270 -148745
rect 75110 -148850 75120 -148750
rect 75210 -148850 75270 -148750
rect 75110 -148855 75270 -148850
rect 75255 -148900 75270 -148855
rect 76070 -148900 76085 -148700
rect 76755 -148745 76770 -148700
rect 76610 -148750 76770 -148745
rect 76610 -148850 76620 -148750
rect 76710 -148850 76770 -148750
rect 76610 -148855 76770 -148850
rect 76755 -148900 76770 -148855
rect 77570 -148900 77585 -148700
rect 78255 -148745 78270 -148700
rect 78110 -148750 78270 -148745
rect 78110 -148850 78120 -148750
rect 78210 -148850 78270 -148750
rect 78110 -148855 78270 -148850
rect 78255 -148900 78270 -148855
rect 79070 -148900 79085 -148700
rect 79755 -148745 79770 -148700
rect 79610 -148750 79770 -148745
rect 79610 -148850 79620 -148750
rect 79710 -148850 79770 -148750
rect 79610 -148855 79770 -148850
rect 79755 -148900 79770 -148855
rect 80570 -148900 80585 -148700
rect 81255 -148745 81270 -148700
rect 81110 -148750 81270 -148745
rect 81110 -148850 81120 -148750
rect 81210 -148850 81270 -148750
rect 81110 -148855 81270 -148850
rect 81255 -148900 81270 -148855
rect 82070 -148900 82085 -148700
rect 82755 -148745 82770 -148700
rect 82610 -148750 82770 -148745
rect 82610 -148850 82620 -148750
rect 82710 -148850 82770 -148750
rect 82610 -148855 82770 -148850
rect 82755 -148900 82770 -148855
rect 83570 -148900 83585 -148700
rect 84255 -148745 84270 -148700
rect 84110 -148750 84270 -148745
rect 84110 -148850 84120 -148750
rect 84210 -148850 84270 -148750
rect 84110 -148855 84270 -148850
rect 84255 -148900 84270 -148855
rect 85070 -148900 85085 -148700
rect 85755 -148745 85770 -148700
rect 85610 -148750 85770 -148745
rect 85610 -148850 85620 -148750
rect 85710 -148850 85770 -148750
rect 85610 -148855 85770 -148850
rect 85755 -148900 85770 -148855
rect 86570 -148900 86585 -148700
rect 87255 -148745 87270 -148700
rect 87110 -148750 87270 -148745
rect 87110 -148850 87120 -148750
rect 87210 -148850 87270 -148750
rect 87110 -148855 87270 -148850
rect 87255 -148900 87270 -148855
rect 88070 -148900 88085 -148700
rect 88755 -148745 88770 -148700
rect 88610 -148750 88770 -148745
rect 88610 -148850 88620 -148750
rect 88710 -148850 88770 -148750
rect 88610 -148855 88770 -148850
rect 88755 -148900 88770 -148855
rect 89570 -148900 89585 -148700
rect 90255 -148745 90270 -148700
rect 90110 -148750 90270 -148745
rect 90110 -148850 90120 -148750
rect 90210 -148850 90270 -148750
rect 90110 -148855 90270 -148850
rect 90255 -148900 90270 -148855
rect 91070 -148900 91085 -148700
rect 91755 -148745 91770 -148700
rect 91610 -148750 91770 -148745
rect 91610 -148850 91620 -148750
rect 91710 -148850 91770 -148750
rect 91610 -148855 91770 -148850
rect 91755 -148900 91770 -148855
rect 92570 -148900 92585 -148700
rect 93255 -148745 93270 -148700
rect 93110 -148750 93270 -148745
rect 93110 -148850 93120 -148750
rect 93210 -148850 93270 -148750
rect 93110 -148855 93270 -148850
rect 93255 -148900 93270 -148855
rect 94070 -148900 94085 -148700
rect 94755 -148745 94770 -148700
rect 94610 -148750 94770 -148745
rect 94610 -148850 94620 -148750
rect 94710 -148850 94770 -148750
rect 94610 -148855 94770 -148850
rect 94755 -148900 94770 -148855
rect 95570 -148900 95585 -148700
rect 96255 -148745 96270 -148700
rect 96110 -148750 96270 -148745
rect 96110 -148850 96120 -148750
rect 96210 -148850 96270 -148750
rect 96110 -148855 96270 -148850
rect 96255 -148900 96270 -148855
rect 97070 -148900 97085 -148700
rect 97755 -148745 97770 -148700
rect 97610 -148750 97770 -148745
rect 97610 -148850 97620 -148750
rect 97710 -148850 97770 -148750
rect 97610 -148855 97770 -148850
rect 97755 -148900 97770 -148855
rect 98570 -148900 98585 -148700
rect 99255 -148745 99270 -148700
rect 99110 -148750 99270 -148745
rect 99110 -148850 99120 -148750
rect 99210 -148850 99270 -148750
rect 99110 -148855 99270 -148850
rect 99255 -148900 99270 -148855
rect 100070 -148900 100085 -148700
rect 100755 -148745 100770 -148700
rect 100610 -148750 100770 -148745
rect 100610 -148850 100620 -148750
rect 100710 -148850 100770 -148750
rect 100610 -148855 100770 -148850
rect 100755 -148900 100770 -148855
rect 101570 -148900 101585 -148700
rect 102255 -148745 102270 -148700
rect 102110 -148750 102270 -148745
rect 102110 -148850 102120 -148750
rect 102210 -148850 102270 -148750
rect 102110 -148855 102270 -148850
rect 102255 -148900 102270 -148855
rect 103070 -148900 103085 -148700
rect 103755 -148745 103770 -148700
rect 103610 -148750 103770 -148745
rect 103610 -148850 103620 -148750
rect 103710 -148850 103770 -148750
rect 103610 -148855 103770 -148850
rect 103755 -148900 103770 -148855
rect 104570 -148900 104585 -148700
rect 105255 -148745 105270 -148700
rect 105110 -148750 105270 -148745
rect 105110 -148850 105120 -148750
rect 105210 -148850 105270 -148750
rect 105110 -148855 105270 -148850
rect 105255 -148900 105270 -148855
rect 106070 -148900 106085 -148700
rect 106755 -148745 106770 -148700
rect 106610 -148750 106770 -148745
rect 106610 -148850 106620 -148750
rect 106710 -148850 106770 -148750
rect 106610 -148855 106770 -148850
rect 106755 -148900 106770 -148855
rect 107570 -148900 107585 -148700
rect 108255 -148745 108270 -148700
rect 108110 -148750 108270 -148745
rect 108110 -148850 108120 -148750
rect 108210 -148850 108270 -148750
rect 108110 -148855 108270 -148850
rect 108255 -148900 108270 -148855
rect 109070 -148900 109085 -148700
rect 109755 -148745 109770 -148700
rect 109610 -148750 109770 -148745
rect 109610 -148850 109620 -148750
rect 109710 -148850 109770 -148750
rect 109610 -148855 109770 -148850
rect 109755 -148900 109770 -148855
rect 110570 -148900 110585 -148700
rect 111255 -148745 111270 -148700
rect 111110 -148750 111270 -148745
rect 111110 -148850 111120 -148750
rect 111210 -148850 111270 -148750
rect 111110 -148855 111270 -148850
rect 111255 -148900 111270 -148855
rect 112070 -148900 112085 -148700
rect 112755 -148745 112770 -148700
rect 112610 -148750 112770 -148745
rect 112610 -148850 112620 -148750
rect 112710 -148850 112770 -148750
rect 112610 -148855 112770 -148850
rect 112755 -148900 112770 -148855
rect 113570 -148900 113585 -148700
rect 114255 -148745 114270 -148700
rect 114110 -148750 114270 -148745
rect 114110 -148850 114120 -148750
rect 114210 -148850 114270 -148750
rect 114110 -148855 114270 -148850
rect 114255 -148900 114270 -148855
rect 115070 -148900 115085 -148700
rect 115755 -148745 115770 -148700
rect 115610 -148750 115770 -148745
rect 115610 -148850 115620 -148750
rect 115710 -148850 115770 -148750
rect 115610 -148855 115770 -148850
rect 115755 -148900 115770 -148855
rect 116570 -148900 116585 -148700
rect 117255 -148745 117270 -148700
rect 117110 -148750 117270 -148745
rect 117110 -148850 117120 -148750
rect 117210 -148850 117270 -148750
rect 117110 -148855 117270 -148850
rect 117255 -148900 117270 -148855
rect 118070 -148900 118085 -148700
rect 118755 -148745 118770 -148700
rect 118610 -148750 118770 -148745
rect 118610 -148850 118620 -148750
rect 118710 -148850 118770 -148750
rect 118610 -148855 118770 -148850
rect 118755 -148900 118770 -148855
rect 119570 -148900 119585 -148700
rect 120255 -148745 120270 -148700
rect 120110 -148750 120270 -148745
rect 120110 -148850 120120 -148750
rect 120210 -148850 120270 -148750
rect 120110 -148855 120270 -148850
rect 120255 -148900 120270 -148855
rect 121070 -148900 121085 -148700
rect 121755 -148745 121770 -148700
rect 121610 -148750 121770 -148745
rect 121610 -148850 121620 -148750
rect 121710 -148850 121770 -148750
rect 121610 -148855 121770 -148850
rect 121755 -148900 121770 -148855
rect 122570 -148900 122585 -148700
rect 123255 -148745 123270 -148700
rect 123110 -148750 123270 -148745
rect 123110 -148850 123120 -148750
rect 123210 -148850 123270 -148750
rect 123110 -148855 123270 -148850
rect 123255 -148900 123270 -148855
rect 124070 -148900 124085 -148700
rect 124755 -148745 124770 -148700
rect 124610 -148750 124770 -148745
rect 124610 -148850 124620 -148750
rect 124710 -148850 124770 -148750
rect 124610 -148855 124770 -148850
rect 124755 -148900 124770 -148855
rect 125570 -148900 125585 -148700
rect 126255 -148745 126270 -148700
rect 126110 -148750 126270 -148745
rect 126110 -148850 126120 -148750
rect 126210 -148850 126270 -148750
rect 126110 -148855 126270 -148850
rect 126255 -148900 126270 -148855
rect 127070 -148900 127085 -148700
rect 127755 -148745 127770 -148700
rect 127610 -148750 127770 -148745
rect 127610 -148850 127620 -148750
rect 127710 -148850 127770 -148750
rect 127610 -148855 127770 -148850
rect 127755 -148900 127770 -148855
rect 128570 -148900 128585 -148700
rect 129255 -148745 129270 -148700
rect 129110 -148750 129270 -148745
rect 129110 -148850 129120 -148750
rect 129210 -148850 129270 -148750
rect 129110 -148855 129270 -148850
rect 129255 -148900 129270 -148855
rect 130070 -148900 130085 -148700
rect 130755 -148745 130770 -148700
rect 130610 -148750 130770 -148745
rect 130610 -148850 130620 -148750
rect 130710 -148850 130770 -148750
rect 130610 -148855 130770 -148850
rect 130755 -148900 130770 -148855
rect 131570 -148900 131585 -148700
rect 132255 -148745 132270 -148700
rect 132110 -148750 132270 -148745
rect 132110 -148850 132120 -148750
rect 132210 -148850 132270 -148750
rect 132110 -148855 132270 -148850
rect 132255 -148900 132270 -148855
rect 133070 -148900 133085 -148700
rect 133755 -148745 133770 -148700
rect 133610 -148750 133770 -148745
rect 133610 -148850 133620 -148750
rect 133710 -148850 133770 -148750
rect 133610 -148855 133770 -148850
rect 133755 -148900 133770 -148855
rect 134570 -148900 134585 -148700
rect 135255 -148745 135270 -148700
rect 135110 -148750 135270 -148745
rect 135110 -148850 135120 -148750
rect 135210 -148850 135270 -148750
rect 135110 -148855 135270 -148850
rect 135255 -148900 135270 -148855
rect 136070 -148900 136085 -148700
rect 136755 -148745 136770 -148700
rect 136610 -148750 136770 -148745
rect 136610 -148850 136620 -148750
rect 136710 -148850 136770 -148750
rect 136610 -148855 136770 -148850
rect 136755 -148900 136770 -148855
rect 137570 -148900 137585 -148700
rect 138255 -148745 138270 -148700
rect 138110 -148750 138270 -148745
rect 138110 -148850 138120 -148750
rect 138210 -148850 138270 -148750
rect 138110 -148855 138270 -148850
rect 138255 -148900 138270 -148855
rect 139070 -148900 139085 -148700
rect 139755 -148745 139770 -148700
rect 139610 -148750 139770 -148745
rect 139610 -148850 139620 -148750
rect 139710 -148850 139770 -148750
rect 139610 -148855 139770 -148850
rect 139755 -148900 139770 -148855
rect 140570 -148900 140585 -148700
rect 141255 -148745 141270 -148700
rect 141110 -148750 141270 -148745
rect 141110 -148850 141120 -148750
rect 141210 -148850 141270 -148750
rect 141110 -148855 141270 -148850
rect 141255 -148900 141270 -148855
rect 142070 -148900 142085 -148700
rect 142755 -148745 142770 -148700
rect 142610 -148750 142770 -148745
rect 142610 -148850 142620 -148750
rect 142710 -148850 142770 -148750
rect 142610 -148855 142770 -148850
rect 142755 -148900 142770 -148855
rect 143570 -148900 143585 -148700
rect 144255 -148745 144270 -148700
rect 144110 -148750 144270 -148745
rect 144110 -148850 144120 -148750
rect 144210 -148850 144270 -148750
rect 144110 -148855 144270 -148850
rect 144255 -148900 144270 -148855
rect 145070 -148900 145085 -148700
rect 145755 -148745 145770 -148700
rect 145610 -148750 145770 -148745
rect 145610 -148850 145620 -148750
rect 145710 -148850 145770 -148750
rect 145610 -148855 145770 -148850
rect 145755 -148900 145770 -148855
rect 146570 -148900 146585 -148700
rect 147255 -148745 147270 -148700
rect 147110 -148750 147270 -148745
rect 147110 -148850 147120 -148750
rect 147210 -148850 147270 -148750
rect 147110 -148855 147270 -148850
rect 147255 -148900 147270 -148855
rect 148070 -148900 148085 -148700
rect 148755 -148745 148770 -148700
rect 148610 -148750 148770 -148745
rect 148610 -148850 148620 -148750
rect 148710 -148850 148770 -148750
rect 148610 -148855 148770 -148850
rect 148755 -148900 148770 -148855
rect 149570 -148900 149585 -148700
<< polycont >>
rect 120 -148850 210 -148750
rect 1620 -148850 1710 -148750
rect 3120 -148850 3210 -148750
rect 4620 -148850 4710 -148750
rect 6120 -148850 6210 -148750
rect 7620 -148850 7710 -148750
rect 9120 -148850 9210 -148750
rect 10620 -148850 10710 -148750
rect 12120 -148850 12210 -148750
rect 13620 -148850 13710 -148750
rect 15120 -148850 15210 -148750
rect 16620 -148850 16710 -148750
rect 18120 -148850 18210 -148750
rect 19620 -148850 19710 -148750
rect 21120 -148850 21210 -148750
rect 22620 -148850 22710 -148750
rect 24120 -148850 24210 -148750
rect 25620 -148850 25710 -148750
rect 27120 -148850 27210 -148750
rect 28620 -148850 28710 -148750
rect 30120 -148850 30210 -148750
rect 31620 -148850 31710 -148750
rect 33120 -148850 33210 -148750
rect 34620 -148850 34710 -148750
rect 36120 -148850 36210 -148750
rect 37620 -148850 37710 -148750
rect 39120 -148850 39210 -148750
rect 40620 -148850 40710 -148750
rect 42120 -148850 42210 -148750
rect 43620 -148850 43710 -148750
rect 45120 -148850 45210 -148750
rect 46620 -148850 46710 -148750
rect 48120 -148850 48210 -148750
rect 49620 -148850 49710 -148750
rect 51120 -148850 51210 -148750
rect 52620 -148850 52710 -148750
rect 54120 -148850 54210 -148750
rect 55620 -148850 55710 -148750
rect 57120 -148850 57210 -148750
rect 58620 -148850 58710 -148750
rect 60120 -148850 60210 -148750
rect 61620 -148850 61710 -148750
rect 63120 -148850 63210 -148750
rect 64620 -148850 64710 -148750
rect 66120 -148850 66210 -148750
rect 67620 -148850 67710 -148750
rect 69120 -148850 69210 -148750
rect 70620 -148850 70710 -148750
rect 72120 -148850 72210 -148750
rect 73620 -148850 73710 -148750
rect 75120 -148850 75210 -148750
rect 76620 -148850 76710 -148750
rect 78120 -148850 78210 -148750
rect 79620 -148850 79710 -148750
rect 81120 -148850 81210 -148750
rect 82620 -148850 82710 -148750
rect 84120 -148850 84210 -148750
rect 85620 -148850 85710 -148750
rect 87120 -148850 87210 -148750
rect 88620 -148850 88710 -148750
rect 90120 -148850 90210 -148750
rect 91620 -148850 91710 -148750
rect 93120 -148850 93210 -148750
rect 94620 -148850 94710 -148750
rect 96120 -148850 96210 -148750
rect 97620 -148850 97710 -148750
rect 99120 -148850 99210 -148750
rect 100620 -148850 100710 -148750
rect 102120 -148850 102210 -148750
rect 103620 -148850 103710 -148750
rect 105120 -148850 105210 -148750
rect 106620 -148850 106710 -148750
rect 108120 -148850 108210 -148750
rect 109620 -148850 109710 -148750
rect 111120 -148850 111210 -148750
rect 112620 -148850 112710 -148750
rect 114120 -148850 114210 -148750
rect 115620 -148850 115710 -148750
rect 117120 -148850 117210 -148750
rect 118620 -148850 118710 -148750
rect 120120 -148850 120210 -148750
rect 121620 -148850 121710 -148750
rect 123120 -148850 123210 -148750
rect 124620 -148850 124710 -148750
rect 126120 -148850 126210 -148750
rect 127620 -148850 127710 -148750
rect 129120 -148850 129210 -148750
rect 130620 -148850 130710 -148750
rect 132120 -148850 132210 -148750
rect 133620 -148850 133710 -148750
rect 135120 -148850 135210 -148750
rect 136620 -148850 136710 -148750
rect 138120 -148850 138210 -148750
rect 139620 -148850 139710 -148750
rect 141120 -148850 141210 -148750
rect 142620 -148850 142710 -148750
rect 144120 -148850 144210 -148750
rect 145620 -148850 145710 -148750
rect 147120 -148850 147210 -148750
rect 148620 -148850 148710 -148750
<< locali >>
rect 270 -148645 280 -148615
rect 1060 -148645 1070 -148615
rect 270 -148660 1070 -148645
rect 270 -148690 280 -148660
rect 1060 -148690 1070 -148660
rect 1770 -148645 1780 -148615
rect 2560 -148645 2570 -148615
rect 1770 -148660 2570 -148645
rect 1770 -148690 1780 -148660
rect 2560 -148690 2570 -148660
rect 3270 -148645 3280 -148615
rect 4060 -148645 4070 -148615
rect 3270 -148660 4070 -148645
rect 3270 -148690 3280 -148660
rect 4060 -148690 4070 -148660
rect 4770 -148645 4780 -148615
rect 5560 -148645 5570 -148615
rect 4770 -148660 5570 -148645
rect 4770 -148690 4780 -148660
rect 5560 -148690 5570 -148660
rect 6270 -148645 6280 -148615
rect 7060 -148645 7070 -148615
rect 6270 -148660 7070 -148645
rect 6270 -148690 6280 -148660
rect 7060 -148690 7070 -148660
rect 7770 -148645 7780 -148615
rect 8560 -148645 8570 -148615
rect 7770 -148660 8570 -148645
rect 7770 -148690 7780 -148660
rect 8560 -148690 8570 -148660
rect 9270 -148645 9280 -148615
rect 10060 -148645 10070 -148615
rect 9270 -148660 10070 -148645
rect 9270 -148690 9280 -148660
rect 10060 -148690 10070 -148660
rect 10770 -148645 10780 -148615
rect 11560 -148645 11570 -148615
rect 10770 -148660 11570 -148645
rect 10770 -148690 10780 -148660
rect 11560 -148690 11570 -148660
rect 12270 -148645 12280 -148615
rect 13060 -148645 13070 -148615
rect 12270 -148660 13070 -148645
rect 12270 -148690 12280 -148660
rect 13060 -148690 13070 -148660
rect 13770 -148645 13780 -148615
rect 14560 -148645 14570 -148615
rect 13770 -148660 14570 -148645
rect 13770 -148690 13780 -148660
rect 14560 -148690 14570 -148660
rect 15270 -148645 15280 -148615
rect 16060 -148645 16070 -148615
rect 15270 -148660 16070 -148645
rect 15270 -148690 15280 -148660
rect 16060 -148690 16070 -148660
rect 16770 -148645 16780 -148615
rect 17560 -148645 17570 -148615
rect 16770 -148660 17570 -148645
rect 16770 -148690 16780 -148660
rect 17560 -148690 17570 -148660
rect 18270 -148645 18280 -148615
rect 19060 -148645 19070 -148615
rect 18270 -148660 19070 -148645
rect 18270 -148690 18280 -148660
rect 19060 -148690 19070 -148660
rect 19770 -148645 19780 -148615
rect 20560 -148645 20570 -148615
rect 19770 -148660 20570 -148645
rect 19770 -148690 19780 -148660
rect 20560 -148690 20570 -148660
rect 21270 -148645 21280 -148615
rect 22060 -148645 22070 -148615
rect 21270 -148660 22070 -148645
rect 21270 -148690 21280 -148660
rect 22060 -148690 22070 -148660
rect 22770 -148645 22780 -148615
rect 23560 -148645 23570 -148615
rect 22770 -148660 23570 -148645
rect 22770 -148690 22780 -148660
rect 23560 -148690 23570 -148660
rect 24270 -148645 24280 -148615
rect 25060 -148645 25070 -148615
rect 24270 -148660 25070 -148645
rect 24270 -148690 24280 -148660
rect 25060 -148690 25070 -148660
rect 25770 -148645 25780 -148615
rect 26560 -148645 26570 -148615
rect 25770 -148660 26570 -148645
rect 25770 -148690 25780 -148660
rect 26560 -148690 26570 -148660
rect 27270 -148645 27280 -148615
rect 28060 -148645 28070 -148615
rect 27270 -148660 28070 -148645
rect 27270 -148690 27280 -148660
rect 28060 -148690 28070 -148660
rect 28770 -148645 28780 -148615
rect 29560 -148645 29570 -148615
rect 28770 -148660 29570 -148645
rect 28770 -148690 28780 -148660
rect 29560 -148690 29570 -148660
rect 30270 -148645 30280 -148615
rect 31060 -148645 31070 -148615
rect 30270 -148660 31070 -148645
rect 30270 -148690 30280 -148660
rect 31060 -148690 31070 -148660
rect 31770 -148645 31780 -148615
rect 32560 -148645 32570 -148615
rect 31770 -148660 32570 -148645
rect 31770 -148690 31780 -148660
rect 32560 -148690 32570 -148660
rect 33270 -148645 33280 -148615
rect 34060 -148645 34070 -148615
rect 33270 -148660 34070 -148645
rect 33270 -148690 33280 -148660
rect 34060 -148690 34070 -148660
rect 34770 -148645 34780 -148615
rect 35560 -148645 35570 -148615
rect 34770 -148660 35570 -148645
rect 34770 -148690 34780 -148660
rect 35560 -148690 35570 -148660
rect 36270 -148645 36280 -148615
rect 37060 -148645 37070 -148615
rect 36270 -148660 37070 -148645
rect 36270 -148690 36280 -148660
rect 37060 -148690 37070 -148660
rect 37770 -148645 37780 -148615
rect 38560 -148645 38570 -148615
rect 37770 -148660 38570 -148645
rect 37770 -148690 37780 -148660
rect 38560 -148690 38570 -148660
rect 39270 -148645 39280 -148615
rect 40060 -148645 40070 -148615
rect 39270 -148660 40070 -148645
rect 39270 -148690 39280 -148660
rect 40060 -148690 40070 -148660
rect 40770 -148645 40780 -148615
rect 41560 -148645 41570 -148615
rect 40770 -148660 41570 -148645
rect 40770 -148690 40780 -148660
rect 41560 -148690 41570 -148660
rect 42270 -148645 42280 -148615
rect 43060 -148645 43070 -148615
rect 42270 -148660 43070 -148645
rect 42270 -148690 42280 -148660
rect 43060 -148690 43070 -148660
rect 43770 -148645 43780 -148615
rect 44560 -148645 44570 -148615
rect 43770 -148660 44570 -148645
rect 43770 -148690 43780 -148660
rect 44560 -148690 44570 -148660
rect 45270 -148645 45280 -148615
rect 46060 -148645 46070 -148615
rect 45270 -148660 46070 -148645
rect 45270 -148690 45280 -148660
rect 46060 -148690 46070 -148660
rect 46770 -148645 46780 -148615
rect 47560 -148645 47570 -148615
rect 46770 -148660 47570 -148645
rect 46770 -148690 46780 -148660
rect 47560 -148690 47570 -148660
rect 48270 -148645 48280 -148615
rect 49060 -148645 49070 -148615
rect 48270 -148660 49070 -148645
rect 48270 -148690 48280 -148660
rect 49060 -148690 49070 -148660
rect 49770 -148645 49780 -148615
rect 50560 -148645 50570 -148615
rect 49770 -148660 50570 -148645
rect 49770 -148690 49780 -148660
rect 50560 -148690 50570 -148660
rect 51270 -148645 51280 -148615
rect 52060 -148645 52070 -148615
rect 51270 -148660 52070 -148645
rect 51270 -148690 51280 -148660
rect 52060 -148690 52070 -148660
rect 52770 -148645 52780 -148615
rect 53560 -148645 53570 -148615
rect 52770 -148660 53570 -148645
rect 52770 -148690 52780 -148660
rect 53560 -148690 53570 -148660
rect 54270 -148645 54280 -148615
rect 55060 -148645 55070 -148615
rect 54270 -148660 55070 -148645
rect 54270 -148690 54280 -148660
rect 55060 -148690 55070 -148660
rect 55770 -148645 55780 -148615
rect 56560 -148645 56570 -148615
rect 55770 -148660 56570 -148645
rect 55770 -148690 55780 -148660
rect 56560 -148690 56570 -148660
rect 57270 -148645 57280 -148615
rect 58060 -148645 58070 -148615
rect 57270 -148660 58070 -148645
rect 57270 -148690 57280 -148660
rect 58060 -148690 58070 -148660
rect 58770 -148645 58780 -148615
rect 59560 -148645 59570 -148615
rect 58770 -148660 59570 -148645
rect 58770 -148690 58780 -148660
rect 59560 -148690 59570 -148660
rect 60270 -148645 60280 -148615
rect 61060 -148645 61070 -148615
rect 60270 -148660 61070 -148645
rect 60270 -148690 60280 -148660
rect 61060 -148690 61070 -148660
rect 61770 -148645 61780 -148615
rect 62560 -148645 62570 -148615
rect 61770 -148660 62570 -148645
rect 61770 -148690 61780 -148660
rect 62560 -148690 62570 -148660
rect 63270 -148645 63280 -148615
rect 64060 -148645 64070 -148615
rect 63270 -148660 64070 -148645
rect 63270 -148690 63280 -148660
rect 64060 -148690 64070 -148660
rect 64770 -148645 64780 -148615
rect 65560 -148645 65570 -148615
rect 64770 -148660 65570 -148645
rect 64770 -148690 64780 -148660
rect 65560 -148690 65570 -148660
rect 66270 -148645 66280 -148615
rect 67060 -148645 67070 -148615
rect 66270 -148660 67070 -148645
rect 66270 -148690 66280 -148660
rect 67060 -148690 67070 -148660
rect 67770 -148645 67780 -148615
rect 68560 -148645 68570 -148615
rect 67770 -148660 68570 -148645
rect 67770 -148690 67780 -148660
rect 68560 -148690 68570 -148660
rect 69270 -148645 69280 -148615
rect 70060 -148645 70070 -148615
rect 69270 -148660 70070 -148645
rect 69270 -148690 69280 -148660
rect 70060 -148690 70070 -148660
rect 70770 -148645 70780 -148615
rect 71560 -148645 71570 -148615
rect 70770 -148660 71570 -148645
rect 70770 -148690 70780 -148660
rect 71560 -148690 71570 -148660
rect 72270 -148645 72280 -148615
rect 73060 -148645 73070 -148615
rect 72270 -148660 73070 -148645
rect 72270 -148690 72280 -148660
rect 73060 -148690 73070 -148660
rect 73770 -148645 73780 -148615
rect 74560 -148645 74570 -148615
rect 73770 -148660 74570 -148645
rect 73770 -148690 73780 -148660
rect 74560 -148690 74570 -148660
rect 75270 -148645 75280 -148615
rect 76060 -148645 76070 -148615
rect 75270 -148660 76070 -148645
rect 75270 -148690 75280 -148660
rect 76060 -148690 76070 -148660
rect 76770 -148645 76780 -148615
rect 77560 -148645 77570 -148615
rect 76770 -148660 77570 -148645
rect 76770 -148690 76780 -148660
rect 77560 -148690 77570 -148660
rect 78270 -148645 78280 -148615
rect 79060 -148645 79070 -148615
rect 78270 -148660 79070 -148645
rect 78270 -148690 78280 -148660
rect 79060 -148690 79070 -148660
rect 79770 -148645 79780 -148615
rect 80560 -148645 80570 -148615
rect 79770 -148660 80570 -148645
rect 79770 -148690 79780 -148660
rect 80560 -148690 80570 -148660
rect 81270 -148645 81280 -148615
rect 82060 -148645 82070 -148615
rect 81270 -148660 82070 -148645
rect 81270 -148690 81280 -148660
rect 82060 -148690 82070 -148660
rect 82770 -148645 82780 -148615
rect 83560 -148645 83570 -148615
rect 82770 -148660 83570 -148645
rect 82770 -148690 82780 -148660
rect 83560 -148690 83570 -148660
rect 84270 -148645 84280 -148615
rect 85060 -148645 85070 -148615
rect 84270 -148660 85070 -148645
rect 84270 -148690 84280 -148660
rect 85060 -148690 85070 -148660
rect 85770 -148645 85780 -148615
rect 86560 -148645 86570 -148615
rect 85770 -148660 86570 -148645
rect 85770 -148690 85780 -148660
rect 86560 -148690 86570 -148660
rect 87270 -148645 87280 -148615
rect 88060 -148645 88070 -148615
rect 87270 -148660 88070 -148645
rect 87270 -148690 87280 -148660
rect 88060 -148690 88070 -148660
rect 88770 -148645 88780 -148615
rect 89560 -148645 89570 -148615
rect 88770 -148660 89570 -148645
rect 88770 -148690 88780 -148660
rect 89560 -148690 89570 -148660
rect 90270 -148645 90280 -148615
rect 91060 -148645 91070 -148615
rect 90270 -148660 91070 -148645
rect 90270 -148690 90280 -148660
rect 91060 -148690 91070 -148660
rect 91770 -148645 91780 -148615
rect 92560 -148645 92570 -148615
rect 91770 -148660 92570 -148645
rect 91770 -148690 91780 -148660
rect 92560 -148690 92570 -148660
rect 93270 -148645 93280 -148615
rect 94060 -148645 94070 -148615
rect 93270 -148660 94070 -148645
rect 93270 -148690 93280 -148660
rect 94060 -148690 94070 -148660
rect 94770 -148645 94780 -148615
rect 95560 -148645 95570 -148615
rect 94770 -148660 95570 -148645
rect 94770 -148690 94780 -148660
rect 95560 -148690 95570 -148660
rect 96270 -148645 96280 -148615
rect 97060 -148645 97070 -148615
rect 96270 -148660 97070 -148645
rect 96270 -148690 96280 -148660
rect 97060 -148690 97070 -148660
rect 97770 -148645 97780 -148615
rect 98560 -148645 98570 -148615
rect 97770 -148660 98570 -148645
rect 97770 -148690 97780 -148660
rect 98560 -148690 98570 -148660
rect 99270 -148645 99280 -148615
rect 100060 -148645 100070 -148615
rect 99270 -148660 100070 -148645
rect 99270 -148690 99280 -148660
rect 100060 -148690 100070 -148660
rect 100770 -148645 100780 -148615
rect 101560 -148645 101570 -148615
rect 100770 -148660 101570 -148645
rect 100770 -148690 100780 -148660
rect 101560 -148690 101570 -148660
rect 102270 -148645 102280 -148615
rect 103060 -148645 103070 -148615
rect 102270 -148660 103070 -148645
rect 102270 -148690 102280 -148660
rect 103060 -148690 103070 -148660
rect 103770 -148645 103780 -148615
rect 104560 -148645 104570 -148615
rect 103770 -148660 104570 -148645
rect 103770 -148690 103780 -148660
rect 104560 -148690 104570 -148660
rect 105270 -148645 105280 -148615
rect 106060 -148645 106070 -148615
rect 105270 -148660 106070 -148645
rect 105270 -148690 105280 -148660
rect 106060 -148690 106070 -148660
rect 106770 -148645 106780 -148615
rect 107560 -148645 107570 -148615
rect 106770 -148660 107570 -148645
rect 106770 -148690 106780 -148660
rect 107560 -148690 107570 -148660
rect 108270 -148645 108280 -148615
rect 109060 -148645 109070 -148615
rect 108270 -148660 109070 -148645
rect 108270 -148690 108280 -148660
rect 109060 -148690 109070 -148660
rect 109770 -148645 109780 -148615
rect 110560 -148645 110570 -148615
rect 109770 -148660 110570 -148645
rect 109770 -148690 109780 -148660
rect 110560 -148690 110570 -148660
rect 111270 -148645 111280 -148615
rect 112060 -148645 112070 -148615
rect 111270 -148660 112070 -148645
rect 111270 -148690 111280 -148660
rect 112060 -148690 112070 -148660
rect 112770 -148645 112780 -148615
rect 113560 -148645 113570 -148615
rect 112770 -148660 113570 -148645
rect 112770 -148690 112780 -148660
rect 113560 -148690 113570 -148660
rect 114270 -148645 114280 -148615
rect 115060 -148645 115070 -148615
rect 114270 -148660 115070 -148645
rect 114270 -148690 114280 -148660
rect 115060 -148690 115070 -148660
rect 115770 -148645 115780 -148615
rect 116560 -148645 116570 -148615
rect 115770 -148660 116570 -148645
rect 115770 -148690 115780 -148660
rect 116560 -148690 116570 -148660
rect 117270 -148645 117280 -148615
rect 118060 -148645 118070 -148615
rect 117270 -148660 118070 -148645
rect 117270 -148690 117280 -148660
rect 118060 -148690 118070 -148660
rect 118770 -148645 118780 -148615
rect 119560 -148645 119570 -148615
rect 118770 -148660 119570 -148645
rect 118770 -148690 118780 -148660
rect 119560 -148690 119570 -148660
rect 120270 -148645 120280 -148615
rect 121060 -148645 121070 -148615
rect 120270 -148660 121070 -148645
rect 120270 -148690 120280 -148660
rect 121060 -148690 121070 -148660
rect 121770 -148645 121780 -148615
rect 122560 -148645 122570 -148615
rect 121770 -148660 122570 -148645
rect 121770 -148690 121780 -148660
rect 122560 -148690 122570 -148660
rect 123270 -148645 123280 -148615
rect 124060 -148645 124070 -148615
rect 123270 -148660 124070 -148645
rect 123270 -148690 123280 -148660
rect 124060 -148690 124070 -148660
rect 124770 -148645 124780 -148615
rect 125560 -148645 125570 -148615
rect 124770 -148660 125570 -148645
rect 124770 -148690 124780 -148660
rect 125560 -148690 125570 -148660
rect 126270 -148645 126280 -148615
rect 127060 -148645 127070 -148615
rect 126270 -148660 127070 -148645
rect 126270 -148690 126280 -148660
rect 127060 -148690 127070 -148660
rect 127770 -148645 127780 -148615
rect 128560 -148645 128570 -148615
rect 127770 -148660 128570 -148645
rect 127770 -148690 127780 -148660
rect 128560 -148690 128570 -148660
rect 129270 -148645 129280 -148615
rect 130060 -148645 130070 -148615
rect 129270 -148660 130070 -148645
rect 129270 -148690 129280 -148660
rect 130060 -148690 130070 -148660
rect 130770 -148645 130780 -148615
rect 131560 -148645 131570 -148615
rect 130770 -148660 131570 -148645
rect 130770 -148690 130780 -148660
rect 131560 -148690 131570 -148660
rect 132270 -148645 132280 -148615
rect 133060 -148645 133070 -148615
rect 132270 -148660 133070 -148645
rect 132270 -148690 132280 -148660
rect 133060 -148690 133070 -148660
rect 133770 -148645 133780 -148615
rect 134560 -148645 134570 -148615
rect 133770 -148660 134570 -148645
rect 133770 -148690 133780 -148660
rect 134560 -148690 134570 -148660
rect 135270 -148645 135280 -148615
rect 136060 -148645 136070 -148615
rect 135270 -148660 136070 -148645
rect 135270 -148690 135280 -148660
rect 136060 -148690 136070 -148660
rect 136770 -148645 136780 -148615
rect 137560 -148645 137570 -148615
rect 136770 -148660 137570 -148645
rect 136770 -148690 136780 -148660
rect 137560 -148690 137570 -148660
rect 138270 -148645 138280 -148615
rect 139060 -148645 139070 -148615
rect 138270 -148660 139070 -148645
rect 138270 -148690 138280 -148660
rect 139060 -148690 139070 -148660
rect 139770 -148645 139780 -148615
rect 140560 -148645 140570 -148615
rect 139770 -148660 140570 -148645
rect 139770 -148690 139780 -148660
rect 140560 -148690 140570 -148660
rect 141270 -148645 141280 -148615
rect 142060 -148645 142070 -148615
rect 141270 -148660 142070 -148645
rect 141270 -148690 141280 -148660
rect 142060 -148690 142070 -148660
rect 142770 -148645 142780 -148615
rect 143560 -148645 143570 -148615
rect 142770 -148660 143570 -148645
rect 142770 -148690 142780 -148660
rect 143560 -148690 143570 -148660
rect 144270 -148645 144280 -148615
rect 145060 -148645 145070 -148615
rect 144270 -148660 145070 -148645
rect 144270 -148690 144280 -148660
rect 145060 -148690 145070 -148660
rect 145770 -148645 145780 -148615
rect 146560 -148645 146570 -148615
rect 145770 -148660 146570 -148645
rect 145770 -148690 145780 -148660
rect 146560 -148690 146570 -148660
rect 147270 -148645 147280 -148615
rect 148060 -148645 148070 -148615
rect 147270 -148660 148070 -148645
rect 147270 -148690 147280 -148660
rect 148060 -148690 148070 -148660
rect 148770 -148645 148780 -148615
rect 149560 -148645 149570 -148615
rect 148770 -148660 149570 -148645
rect 148770 -148690 148780 -148660
rect 149560 -148690 149570 -148660
rect 110 -148750 220 -148745
rect 110 -148850 120 -148750
rect 210 -148850 220 -148750
rect 110 -148855 220 -148850
rect 1610 -148750 1720 -148745
rect 1610 -148850 1620 -148750
rect 1710 -148850 1720 -148750
rect 1610 -148855 1720 -148850
rect 3110 -148750 3220 -148745
rect 3110 -148850 3120 -148750
rect 3210 -148850 3220 -148750
rect 3110 -148855 3220 -148850
rect 4610 -148750 4720 -148745
rect 4610 -148850 4620 -148750
rect 4710 -148850 4720 -148750
rect 4610 -148855 4720 -148850
rect 6110 -148750 6220 -148745
rect 6110 -148850 6120 -148750
rect 6210 -148850 6220 -148750
rect 6110 -148855 6220 -148850
rect 7610 -148750 7720 -148745
rect 7610 -148850 7620 -148750
rect 7710 -148850 7720 -148750
rect 7610 -148855 7720 -148850
rect 9110 -148750 9220 -148745
rect 9110 -148850 9120 -148750
rect 9210 -148850 9220 -148750
rect 9110 -148855 9220 -148850
rect 10610 -148750 10720 -148745
rect 10610 -148850 10620 -148750
rect 10710 -148850 10720 -148750
rect 10610 -148855 10720 -148850
rect 12110 -148750 12220 -148745
rect 12110 -148850 12120 -148750
rect 12210 -148850 12220 -148750
rect 12110 -148855 12220 -148850
rect 13610 -148750 13720 -148745
rect 13610 -148850 13620 -148750
rect 13710 -148850 13720 -148750
rect 13610 -148855 13720 -148850
rect 15110 -148750 15220 -148745
rect 15110 -148850 15120 -148750
rect 15210 -148850 15220 -148750
rect 15110 -148855 15220 -148850
rect 16610 -148750 16720 -148745
rect 16610 -148850 16620 -148750
rect 16710 -148850 16720 -148750
rect 16610 -148855 16720 -148850
rect 18110 -148750 18220 -148745
rect 18110 -148850 18120 -148750
rect 18210 -148850 18220 -148750
rect 18110 -148855 18220 -148850
rect 19610 -148750 19720 -148745
rect 19610 -148850 19620 -148750
rect 19710 -148850 19720 -148750
rect 19610 -148855 19720 -148850
rect 21110 -148750 21220 -148745
rect 21110 -148850 21120 -148750
rect 21210 -148850 21220 -148750
rect 21110 -148855 21220 -148850
rect 22610 -148750 22720 -148745
rect 22610 -148850 22620 -148750
rect 22710 -148850 22720 -148750
rect 22610 -148855 22720 -148850
rect 24110 -148750 24220 -148745
rect 24110 -148850 24120 -148750
rect 24210 -148850 24220 -148750
rect 24110 -148855 24220 -148850
rect 25610 -148750 25720 -148745
rect 25610 -148850 25620 -148750
rect 25710 -148850 25720 -148750
rect 25610 -148855 25720 -148850
rect 27110 -148750 27220 -148745
rect 27110 -148850 27120 -148750
rect 27210 -148850 27220 -148750
rect 27110 -148855 27220 -148850
rect 28610 -148750 28720 -148745
rect 28610 -148850 28620 -148750
rect 28710 -148850 28720 -148750
rect 28610 -148855 28720 -148850
rect 30110 -148750 30220 -148745
rect 30110 -148850 30120 -148750
rect 30210 -148850 30220 -148750
rect 30110 -148855 30220 -148850
rect 31610 -148750 31720 -148745
rect 31610 -148850 31620 -148750
rect 31710 -148850 31720 -148750
rect 31610 -148855 31720 -148850
rect 33110 -148750 33220 -148745
rect 33110 -148850 33120 -148750
rect 33210 -148850 33220 -148750
rect 33110 -148855 33220 -148850
rect 34610 -148750 34720 -148745
rect 34610 -148850 34620 -148750
rect 34710 -148850 34720 -148750
rect 34610 -148855 34720 -148850
rect 36110 -148750 36220 -148745
rect 36110 -148850 36120 -148750
rect 36210 -148850 36220 -148750
rect 36110 -148855 36220 -148850
rect 37610 -148750 37720 -148745
rect 37610 -148850 37620 -148750
rect 37710 -148850 37720 -148750
rect 37610 -148855 37720 -148850
rect 39110 -148750 39220 -148745
rect 39110 -148850 39120 -148750
rect 39210 -148850 39220 -148750
rect 39110 -148855 39220 -148850
rect 40610 -148750 40720 -148745
rect 40610 -148850 40620 -148750
rect 40710 -148850 40720 -148750
rect 40610 -148855 40720 -148850
rect 42110 -148750 42220 -148745
rect 42110 -148850 42120 -148750
rect 42210 -148850 42220 -148750
rect 42110 -148855 42220 -148850
rect 43610 -148750 43720 -148745
rect 43610 -148850 43620 -148750
rect 43710 -148850 43720 -148750
rect 43610 -148855 43720 -148850
rect 45110 -148750 45220 -148745
rect 45110 -148850 45120 -148750
rect 45210 -148850 45220 -148750
rect 45110 -148855 45220 -148850
rect 46610 -148750 46720 -148745
rect 46610 -148850 46620 -148750
rect 46710 -148850 46720 -148750
rect 46610 -148855 46720 -148850
rect 48110 -148750 48220 -148745
rect 48110 -148850 48120 -148750
rect 48210 -148850 48220 -148750
rect 48110 -148855 48220 -148850
rect 49610 -148750 49720 -148745
rect 49610 -148850 49620 -148750
rect 49710 -148850 49720 -148750
rect 49610 -148855 49720 -148850
rect 51110 -148750 51220 -148745
rect 51110 -148850 51120 -148750
rect 51210 -148850 51220 -148750
rect 51110 -148855 51220 -148850
rect 52610 -148750 52720 -148745
rect 52610 -148850 52620 -148750
rect 52710 -148850 52720 -148750
rect 52610 -148855 52720 -148850
rect 54110 -148750 54220 -148745
rect 54110 -148850 54120 -148750
rect 54210 -148850 54220 -148750
rect 54110 -148855 54220 -148850
rect 55610 -148750 55720 -148745
rect 55610 -148850 55620 -148750
rect 55710 -148850 55720 -148750
rect 55610 -148855 55720 -148850
rect 57110 -148750 57220 -148745
rect 57110 -148850 57120 -148750
rect 57210 -148850 57220 -148750
rect 57110 -148855 57220 -148850
rect 58610 -148750 58720 -148745
rect 58610 -148850 58620 -148750
rect 58710 -148850 58720 -148750
rect 58610 -148855 58720 -148850
rect 60110 -148750 60220 -148745
rect 60110 -148850 60120 -148750
rect 60210 -148850 60220 -148750
rect 60110 -148855 60220 -148850
rect 61610 -148750 61720 -148745
rect 61610 -148850 61620 -148750
rect 61710 -148850 61720 -148750
rect 61610 -148855 61720 -148850
rect 63110 -148750 63220 -148745
rect 63110 -148850 63120 -148750
rect 63210 -148850 63220 -148750
rect 63110 -148855 63220 -148850
rect 64610 -148750 64720 -148745
rect 64610 -148850 64620 -148750
rect 64710 -148850 64720 -148750
rect 64610 -148855 64720 -148850
rect 66110 -148750 66220 -148745
rect 66110 -148850 66120 -148750
rect 66210 -148850 66220 -148750
rect 66110 -148855 66220 -148850
rect 67610 -148750 67720 -148745
rect 67610 -148850 67620 -148750
rect 67710 -148850 67720 -148750
rect 67610 -148855 67720 -148850
rect 69110 -148750 69220 -148745
rect 69110 -148850 69120 -148750
rect 69210 -148850 69220 -148750
rect 69110 -148855 69220 -148850
rect 70610 -148750 70720 -148745
rect 70610 -148850 70620 -148750
rect 70710 -148850 70720 -148750
rect 70610 -148855 70720 -148850
rect 72110 -148750 72220 -148745
rect 72110 -148850 72120 -148750
rect 72210 -148850 72220 -148750
rect 72110 -148855 72220 -148850
rect 73610 -148750 73720 -148745
rect 73610 -148850 73620 -148750
rect 73710 -148850 73720 -148750
rect 73610 -148855 73720 -148850
rect 75110 -148750 75220 -148745
rect 75110 -148850 75120 -148750
rect 75210 -148850 75220 -148750
rect 75110 -148855 75220 -148850
rect 76610 -148750 76720 -148745
rect 76610 -148850 76620 -148750
rect 76710 -148850 76720 -148750
rect 76610 -148855 76720 -148850
rect 78110 -148750 78220 -148745
rect 78110 -148850 78120 -148750
rect 78210 -148850 78220 -148750
rect 78110 -148855 78220 -148850
rect 79610 -148750 79720 -148745
rect 79610 -148850 79620 -148750
rect 79710 -148850 79720 -148750
rect 79610 -148855 79720 -148850
rect 81110 -148750 81220 -148745
rect 81110 -148850 81120 -148750
rect 81210 -148850 81220 -148750
rect 81110 -148855 81220 -148850
rect 82610 -148750 82720 -148745
rect 82610 -148850 82620 -148750
rect 82710 -148850 82720 -148750
rect 82610 -148855 82720 -148850
rect 84110 -148750 84220 -148745
rect 84110 -148850 84120 -148750
rect 84210 -148850 84220 -148750
rect 84110 -148855 84220 -148850
rect 85610 -148750 85720 -148745
rect 85610 -148850 85620 -148750
rect 85710 -148850 85720 -148750
rect 85610 -148855 85720 -148850
rect 87110 -148750 87220 -148745
rect 87110 -148850 87120 -148750
rect 87210 -148850 87220 -148750
rect 87110 -148855 87220 -148850
rect 88610 -148750 88720 -148745
rect 88610 -148850 88620 -148750
rect 88710 -148850 88720 -148750
rect 88610 -148855 88720 -148850
rect 90110 -148750 90220 -148745
rect 90110 -148850 90120 -148750
rect 90210 -148850 90220 -148750
rect 90110 -148855 90220 -148850
rect 91610 -148750 91720 -148745
rect 91610 -148850 91620 -148750
rect 91710 -148850 91720 -148750
rect 91610 -148855 91720 -148850
rect 93110 -148750 93220 -148745
rect 93110 -148850 93120 -148750
rect 93210 -148850 93220 -148750
rect 93110 -148855 93220 -148850
rect 94610 -148750 94720 -148745
rect 94610 -148850 94620 -148750
rect 94710 -148850 94720 -148750
rect 94610 -148855 94720 -148850
rect 96110 -148750 96220 -148745
rect 96110 -148850 96120 -148750
rect 96210 -148850 96220 -148750
rect 96110 -148855 96220 -148850
rect 97610 -148750 97720 -148745
rect 97610 -148850 97620 -148750
rect 97710 -148850 97720 -148750
rect 97610 -148855 97720 -148850
rect 99110 -148750 99220 -148745
rect 99110 -148850 99120 -148750
rect 99210 -148850 99220 -148750
rect 99110 -148855 99220 -148850
rect 100610 -148750 100720 -148745
rect 100610 -148850 100620 -148750
rect 100710 -148850 100720 -148750
rect 100610 -148855 100720 -148850
rect 102110 -148750 102220 -148745
rect 102110 -148850 102120 -148750
rect 102210 -148850 102220 -148750
rect 102110 -148855 102220 -148850
rect 103610 -148750 103720 -148745
rect 103610 -148850 103620 -148750
rect 103710 -148850 103720 -148750
rect 103610 -148855 103720 -148850
rect 105110 -148750 105220 -148745
rect 105110 -148850 105120 -148750
rect 105210 -148850 105220 -148750
rect 105110 -148855 105220 -148850
rect 106610 -148750 106720 -148745
rect 106610 -148850 106620 -148750
rect 106710 -148850 106720 -148750
rect 106610 -148855 106720 -148850
rect 108110 -148750 108220 -148745
rect 108110 -148850 108120 -148750
rect 108210 -148850 108220 -148750
rect 108110 -148855 108220 -148850
rect 109610 -148750 109720 -148745
rect 109610 -148850 109620 -148750
rect 109710 -148850 109720 -148750
rect 109610 -148855 109720 -148850
rect 111110 -148750 111220 -148745
rect 111110 -148850 111120 -148750
rect 111210 -148850 111220 -148750
rect 111110 -148855 111220 -148850
rect 112610 -148750 112720 -148745
rect 112610 -148850 112620 -148750
rect 112710 -148850 112720 -148750
rect 112610 -148855 112720 -148850
rect 114110 -148750 114220 -148745
rect 114110 -148850 114120 -148750
rect 114210 -148850 114220 -148750
rect 114110 -148855 114220 -148850
rect 115610 -148750 115720 -148745
rect 115610 -148850 115620 -148750
rect 115710 -148850 115720 -148750
rect 115610 -148855 115720 -148850
rect 117110 -148750 117220 -148745
rect 117110 -148850 117120 -148750
rect 117210 -148850 117220 -148750
rect 117110 -148855 117220 -148850
rect 118610 -148750 118720 -148745
rect 118610 -148850 118620 -148750
rect 118710 -148850 118720 -148750
rect 118610 -148855 118720 -148850
rect 120110 -148750 120220 -148745
rect 120110 -148850 120120 -148750
rect 120210 -148850 120220 -148750
rect 120110 -148855 120220 -148850
rect 121610 -148750 121720 -148745
rect 121610 -148850 121620 -148750
rect 121710 -148850 121720 -148750
rect 121610 -148855 121720 -148850
rect 123110 -148750 123220 -148745
rect 123110 -148850 123120 -148750
rect 123210 -148850 123220 -148750
rect 123110 -148855 123220 -148850
rect 124610 -148750 124720 -148745
rect 124610 -148850 124620 -148750
rect 124710 -148850 124720 -148750
rect 124610 -148855 124720 -148850
rect 126110 -148750 126220 -148745
rect 126110 -148850 126120 -148750
rect 126210 -148850 126220 -148750
rect 126110 -148855 126220 -148850
rect 127610 -148750 127720 -148745
rect 127610 -148850 127620 -148750
rect 127710 -148850 127720 -148750
rect 127610 -148855 127720 -148850
rect 129110 -148750 129220 -148745
rect 129110 -148850 129120 -148750
rect 129210 -148850 129220 -148750
rect 129110 -148855 129220 -148850
rect 130610 -148750 130720 -148745
rect 130610 -148850 130620 -148750
rect 130710 -148850 130720 -148750
rect 130610 -148855 130720 -148850
rect 132110 -148750 132220 -148745
rect 132110 -148850 132120 -148750
rect 132210 -148850 132220 -148750
rect 132110 -148855 132220 -148850
rect 133610 -148750 133720 -148745
rect 133610 -148850 133620 -148750
rect 133710 -148850 133720 -148750
rect 133610 -148855 133720 -148850
rect 135110 -148750 135220 -148745
rect 135110 -148850 135120 -148750
rect 135210 -148850 135220 -148750
rect 135110 -148855 135220 -148850
rect 136610 -148750 136720 -148745
rect 136610 -148850 136620 -148750
rect 136710 -148850 136720 -148750
rect 136610 -148855 136720 -148850
rect 138110 -148750 138220 -148745
rect 138110 -148850 138120 -148750
rect 138210 -148850 138220 -148750
rect 138110 -148855 138220 -148850
rect 139610 -148750 139720 -148745
rect 139610 -148850 139620 -148750
rect 139710 -148850 139720 -148750
rect 139610 -148855 139720 -148850
rect 141110 -148750 141220 -148745
rect 141110 -148850 141120 -148750
rect 141210 -148850 141220 -148750
rect 141110 -148855 141220 -148850
rect 142610 -148750 142720 -148745
rect 142610 -148850 142620 -148750
rect 142710 -148850 142720 -148750
rect 142610 -148855 142720 -148850
rect 144110 -148750 144220 -148745
rect 144110 -148850 144120 -148750
rect 144210 -148850 144220 -148750
rect 144110 -148855 144220 -148850
rect 145610 -148750 145720 -148745
rect 145610 -148850 145620 -148750
rect 145710 -148850 145720 -148750
rect 145610 -148855 145720 -148850
rect 147110 -148750 147220 -148745
rect 147110 -148850 147120 -148750
rect 147210 -148850 147220 -148750
rect 147110 -148855 147220 -148850
rect 148610 -148750 148720 -148745
rect 148610 -148850 148620 -148750
rect 148710 -148850 148720 -148750
rect 148610 -148855 148720 -148850
rect 270 -148915 1070 -148900
rect 270 -148935 280 -148915
rect 1060 -148935 1070 -148915
rect 270 -148960 1070 -148935
rect 270 -148990 280 -148960
rect 1060 -148990 1070 -148960
rect 270 -149000 1070 -148990
rect 1770 -148915 2570 -148900
rect 1770 -148935 1780 -148915
rect 2560 -148935 2570 -148915
rect 1770 -148960 2570 -148935
rect 1770 -148990 1780 -148960
rect 2560 -148990 2570 -148960
rect 1770 -149000 2570 -148990
rect 3270 -148915 4070 -148900
rect 3270 -148935 3280 -148915
rect 4060 -148935 4070 -148915
rect 3270 -148960 4070 -148935
rect 3270 -148990 3280 -148960
rect 4060 -148990 4070 -148960
rect 3270 -149000 4070 -148990
rect 4770 -148915 5570 -148900
rect 4770 -148935 4780 -148915
rect 5560 -148935 5570 -148915
rect 4770 -148960 5570 -148935
rect 4770 -148990 4780 -148960
rect 5560 -148990 5570 -148960
rect 4770 -149000 5570 -148990
rect 6270 -148915 7070 -148900
rect 6270 -148935 6280 -148915
rect 7060 -148935 7070 -148915
rect 6270 -148960 7070 -148935
rect 6270 -148990 6280 -148960
rect 7060 -148990 7070 -148960
rect 6270 -149000 7070 -148990
rect 7770 -148915 8570 -148900
rect 7770 -148935 7780 -148915
rect 8560 -148935 8570 -148915
rect 7770 -148960 8570 -148935
rect 7770 -148990 7780 -148960
rect 8560 -148990 8570 -148960
rect 7770 -149000 8570 -148990
rect 9270 -148915 10070 -148900
rect 9270 -148935 9280 -148915
rect 10060 -148935 10070 -148915
rect 9270 -148960 10070 -148935
rect 9270 -148990 9280 -148960
rect 10060 -148990 10070 -148960
rect 9270 -149000 10070 -148990
rect 10770 -148915 11570 -148900
rect 10770 -148935 10780 -148915
rect 11560 -148935 11570 -148915
rect 10770 -148960 11570 -148935
rect 10770 -148990 10780 -148960
rect 11560 -148990 11570 -148960
rect 10770 -149000 11570 -148990
rect 12270 -148915 13070 -148900
rect 12270 -148935 12280 -148915
rect 13060 -148935 13070 -148915
rect 12270 -148960 13070 -148935
rect 12270 -148990 12280 -148960
rect 13060 -148990 13070 -148960
rect 12270 -149000 13070 -148990
rect 13770 -148915 14570 -148900
rect 13770 -148935 13780 -148915
rect 14560 -148935 14570 -148915
rect 13770 -148960 14570 -148935
rect 13770 -148990 13780 -148960
rect 14560 -148990 14570 -148960
rect 13770 -149000 14570 -148990
rect 15270 -148915 16070 -148900
rect 15270 -148935 15280 -148915
rect 16060 -148935 16070 -148915
rect 15270 -148960 16070 -148935
rect 15270 -148990 15280 -148960
rect 16060 -148990 16070 -148960
rect 15270 -149000 16070 -148990
rect 16770 -148915 17570 -148900
rect 16770 -148935 16780 -148915
rect 17560 -148935 17570 -148915
rect 16770 -148960 17570 -148935
rect 16770 -148990 16780 -148960
rect 17560 -148990 17570 -148960
rect 16770 -149000 17570 -148990
rect 18270 -148915 19070 -148900
rect 18270 -148935 18280 -148915
rect 19060 -148935 19070 -148915
rect 18270 -148960 19070 -148935
rect 18270 -148990 18280 -148960
rect 19060 -148990 19070 -148960
rect 18270 -149000 19070 -148990
rect 19770 -148915 20570 -148900
rect 19770 -148935 19780 -148915
rect 20560 -148935 20570 -148915
rect 19770 -148960 20570 -148935
rect 19770 -148990 19780 -148960
rect 20560 -148990 20570 -148960
rect 19770 -149000 20570 -148990
rect 21270 -148915 22070 -148900
rect 21270 -148935 21280 -148915
rect 22060 -148935 22070 -148915
rect 21270 -148960 22070 -148935
rect 21270 -148990 21280 -148960
rect 22060 -148990 22070 -148960
rect 21270 -149000 22070 -148990
rect 22770 -148915 23570 -148900
rect 22770 -148935 22780 -148915
rect 23560 -148935 23570 -148915
rect 22770 -148960 23570 -148935
rect 22770 -148990 22780 -148960
rect 23560 -148990 23570 -148960
rect 22770 -149000 23570 -148990
rect 24270 -148915 25070 -148900
rect 24270 -148935 24280 -148915
rect 25060 -148935 25070 -148915
rect 24270 -148960 25070 -148935
rect 24270 -148990 24280 -148960
rect 25060 -148990 25070 -148960
rect 24270 -149000 25070 -148990
rect 25770 -148915 26570 -148900
rect 25770 -148935 25780 -148915
rect 26560 -148935 26570 -148915
rect 25770 -148960 26570 -148935
rect 25770 -148990 25780 -148960
rect 26560 -148990 26570 -148960
rect 25770 -149000 26570 -148990
rect 27270 -148915 28070 -148900
rect 27270 -148935 27280 -148915
rect 28060 -148935 28070 -148915
rect 27270 -148960 28070 -148935
rect 27270 -148990 27280 -148960
rect 28060 -148990 28070 -148960
rect 27270 -149000 28070 -148990
rect 28770 -148915 29570 -148900
rect 28770 -148935 28780 -148915
rect 29560 -148935 29570 -148915
rect 28770 -148960 29570 -148935
rect 28770 -148990 28780 -148960
rect 29560 -148990 29570 -148960
rect 28770 -149000 29570 -148990
rect 30270 -148915 31070 -148900
rect 30270 -148935 30280 -148915
rect 31060 -148935 31070 -148915
rect 30270 -148960 31070 -148935
rect 30270 -148990 30280 -148960
rect 31060 -148990 31070 -148960
rect 30270 -149000 31070 -148990
rect 31770 -148915 32570 -148900
rect 31770 -148935 31780 -148915
rect 32560 -148935 32570 -148915
rect 31770 -148960 32570 -148935
rect 31770 -148990 31780 -148960
rect 32560 -148990 32570 -148960
rect 31770 -149000 32570 -148990
rect 33270 -148915 34070 -148900
rect 33270 -148935 33280 -148915
rect 34060 -148935 34070 -148915
rect 33270 -148960 34070 -148935
rect 33270 -148990 33280 -148960
rect 34060 -148990 34070 -148960
rect 33270 -149000 34070 -148990
rect 34770 -148915 35570 -148900
rect 34770 -148935 34780 -148915
rect 35560 -148935 35570 -148915
rect 34770 -148960 35570 -148935
rect 34770 -148990 34780 -148960
rect 35560 -148990 35570 -148960
rect 34770 -149000 35570 -148990
rect 36270 -148915 37070 -148900
rect 36270 -148935 36280 -148915
rect 37060 -148935 37070 -148915
rect 36270 -148960 37070 -148935
rect 36270 -148990 36280 -148960
rect 37060 -148990 37070 -148960
rect 36270 -149000 37070 -148990
rect 37770 -148915 38570 -148900
rect 37770 -148935 37780 -148915
rect 38560 -148935 38570 -148915
rect 37770 -148960 38570 -148935
rect 37770 -148990 37780 -148960
rect 38560 -148990 38570 -148960
rect 37770 -149000 38570 -148990
rect 39270 -148915 40070 -148900
rect 39270 -148935 39280 -148915
rect 40060 -148935 40070 -148915
rect 39270 -148960 40070 -148935
rect 39270 -148990 39280 -148960
rect 40060 -148990 40070 -148960
rect 39270 -149000 40070 -148990
rect 40770 -148915 41570 -148900
rect 40770 -148935 40780 -148915
rect 41560 -148935 41570 -148915
rect 40770 -148960 41570 -148935
rect 40770 -148990 40780 -148960
rect 41560 -148990 41570 -148960
rect 40770 -149000 41570 -148990
rect 42270 -148915 43070 -148900
rect 42270 -148935 42280 -148915
rect 43060 -148935 43070 -148915
rect 42270 -148960 43070 -148935
rect 42270 -148990 42280 -148960
rect 43060 -148990 43070 -148960
rect 42270 -149000 43070 -148990
rect 43770 -148915 44570 -148900
rect 43770 -148935 43780 -148915
rect 44560 -148935 44570 -148915
rect 43770 -148960 44570 -148935
rect 43770 -148990 43780 -148960
rect 44560 -148990 44570 -148960
rect 43770 -149000 44570 -148990
rect 45270 -148915 46070 -148900
rect 45270 -148935 45280 -148915
rect 46060 -148935 46070 -148915
rect 45270 -148960 46070 -148935
rect 45270 -148990 45280 -148960
rect 46060 -148990 46070 -148960
rect 45270 -149000 46070 -148990
rect 46770 -148915 47570 -148900
rect 46770 -148935 46780 -148915
rect 47560 -148935 47570 -148915
rect 46770 -148960 47570 -148935
rect 46770 -148990 46780 -148960
rect 47560 -148990 47570 -148960
rect 46770 -149000 47570 -148990
rect 48270 -148915 49070 -148900
rect 48270 -148935 48280 -148915
rect 49060 -148935 49070 -148915
rect 48270 -148960 49070 -148935
rect 48270 -148990 48280 -148960
rect 49060 -148990 49070 -148960
rect 48270 -149000 49070 -148990
rect 49770 -148915 50570 -148900
rect 49770 -148935 49780 -148915
rect 50560 -148935 50570 -148915
rect 49770 -148960 50570 -148935
rect 49770 -148990 49780 -148960
rect 50560 -148990 50570 -148960
rect 49770 -149000 50570 -148990
rect 51270 -148915 52070 -148900
rect 51270 -148935 51280 -148915
rect 52060 -148935 52070 -148915
rect 51270 -148960 52070 -148935
rect 51270 -148990 51280 -148960
rect 52060 -148990 52070 -148960
rect 51270 -149000 52070 -148990
rect 52770 -148915 53570 -148900
rect 52770 -148935 52780 -148915
rect 53560 -148935 53570 -148915
rect 52770 -148960 53570 -148935
rect 52770 -148990 52780 -148960
rect 53560 -148990 53570 -148960
rect 52770 -149000 53570 -148990
rect 54270 -148915 55070 -148900
rect 54270 -148935 54280 -148915
rect 55060 -148935 55070 -148915
rect 54270 -148960 55070 -148935
rect 54270 -148990 54280 -148960
rect 55060 -148990 55070 -148960
rect 54270 -149000 55070 -148990
rect 55770 -148915 56570 -148900
rect 55770 -148935 55780 -148915
rect 56560 -148935 56570 -148915
rect 55770 -148960 56570 -148935
rect 55770 -148990 55780 -148960
rect 56560 -148990 56570 -148960
rect 55770 -149000 56570 -148990
rect 57270 -148915 58070 -148900
rect 57270 -148935 57280 -148915
rect 58060 -148935 58070 -148915
rect 57270 -148960 58070 -148935
rect 57270 -148990 57280 -148960
rect 58060 -148990 58070 -148960
rect 57270 -149000 58070 -148990
rect 58770 -148915 59570 -148900
rect 58770 -148935 58780 -148915
rect 59560 -148935 59570 -148915
rect 58770 -148960 59570 -148935
rect 58770 -148990 58780 -148960
rect 59560 -148990 59570 -148960
rect 58770 -149000 59570 -148990
rect 60270 -148915 61070 -148900
rect 60270 -148935 60280 -148915
rect 61060 -148935 61070 -148915
rect 60270 -148960 61070 -148935
rect 60270 -148990 60280 -148960
rect 61060 -148990 61070 -148960
rect 60270 -149000 61070 -148990
rect 61770 -148915 62570 -148900
rect 61770 -148935 61780 -148915
rect 62560 -148935 62570 -148915
rect 61770 -148960 62570 -148935
rect 61770 -148990 61780 -148960
rect 62560 -148990 62570 -148960
rect 61770 -149000 62570 -148990
rect 63270 -148915 64070 -148900
rect 63270 -148935 63280 -148915
rect 64060 -148935 64070 -148915
rect 63270 -148960 64070 -148935
rect 63270 -148990 63280 -148960
rect 64060 -148990 64070 -148960
rect 63270 -149000 64070 -148990
rect 64770 -148915 65570 -148900
rect 64770 -148935 64780 -148915
rect 65560 -148935 65570 -148915
rect 64770 -148960 65570 -148935
rect 64770 -148990 64780 -148960
rect 65560 -148990 65570 -148960
rect 64770 -149000 65570 -148990
rect 66270 -148915 67070 -148900
rect 66270 -148935 66280 -148915
rect 67060 -148935 67070 -148915
rect 66270 -148960 67070 -148935
rect 66270 -148990 66280 -148960
rect 67060 -148990 67070 -148960
rect 66270 -149000 67070 -148990
rect 67770 -148915 68570 -148900
rect 67770 -148935 67780 -148915
rect 68560 -148935 68570 -148915
rect 67770 -148960 68570 -148935
rect 67770 -148990 67780 -148960
rect 68560 -148990 68570 -148960
rect 67770 -149000 68570 -148990
rect 69270 -148915 70070 -148900
rect 69270 -148935 69280 -148915
rect 70060 -148935 70070 -148915
rect 69270 -148960 70070 -148935
rect 69270 -148990 69280 -148960
rect 70060 -148990 70070 -148960
rect 69270 -149000 70070 -148990
rect 70770 -148915 71570 -148900
rect 70770 -148935 70780 -148915
rect 71560 -148935 71570 -148915
rect 70770 -148960 71570 -148935
rect 70770 -148990 70780 -148960
rect 71560 -148990 71570 -148960
rect 70770 -149000 71570 -148990
rect 72270 -148915 73070 -148900
rect 72270 -148935 72280 -148915
rect 73060 -148935 73070 -148915
rect 72270 -148960 73070 -148935
rect 72270 -148990 72280 -148960
rect 73060 -148990 73070 -148960
rect 72270 -149000 73070 -148990
rect 73770 -148915 74570 -148900
rect 73770 -148935 73780 -148915
rect 74560 -148935 74570 -148915
rect 73770 -148960 74570 -148935
rect 73770 -148990 73780 -148960
rect 74560 -148990 74570 -148960
rect 73770 -149000 74570 -148990
rect 75270 -148915 76070 -148900
rect 75270 -148935 75280 -148915
rect 76060 -148935 76070 -148915
rect 75270 -148960 76070 -148935
rect 75270 -148990 75280 -148960
rect 76060 -148990 76070 -148960
rect 75270 -149000 76070 -148990
rect 76770 -148915 77570 -148900
rect 76770 -148935 76780 -148915
rect 77560 -148935 77570 -148915
rect 76770 -148960 77570 -148935
rect 76770 -148990 76780 -148960
rect 77560 -148990 77570 -148960
rect 76770 -149000 77570 -148990
rect 78270 -148915 79070 -148900
rect 78270 -148935 78280 -148915
rect 79060 -148935 79070 -148915
rect 78270 -148960 79070 -148935
rect 78270 -148990 78280 -148960
rect 79060 -148990 79070 -148960
rect 78270 -149000 79070 -148990
rect 79770 -148915 80570 -148900
rect 79770 -148935 79780 -148915
rect 80560 -148935 80570 -148915
rect 79770 -148960 80570 -148935
rect 79770 -148990 79780 -148960
rect 80560 -148990 80570 -148960
rect 79770 -149000 80570 -148990
rect 81270 -148915 82070 -148900
rect 81270 -148935 81280 -148915
rect 82060 -148935 82070 -148915
rect 81270 -148960 82070 -148935
rect 81270 -148990 81280 -148960
rect 82060 -148990 82070 -148960
rect 81270 -149000 82070 -148990
rect 82770 -148915 83570 -148900
rect 82770 -148935 82780 -148915
rect 83560 -148935 83570 -148915
rect 82770 -148960 83570 -148935
rect 82770 -148990 82780 -148960
rect 83560 -148990 83570 -148960
rect 82770 -149000 83570 -148990
rect 84270 -148915 85070 -148900
rect 84270 -148935 84280 -148915
rect 85060 -148935 85070 -148915
rect 84270 -148960 85070 -148935
rect 84270 -148990 84280 -148960
rect 85060 -148990 85070 -148960
rect 84270 -149000 85070 -148990
rect 85770 -148915 86570 -148900
rect 85770 -148935 85780 -148915
rect 86560 -148935 86570 -148915
rect 85770 -148960 86570 -148935
rect 85770 -148990 85780 -148960
rect 86560 -148990 86570 -148960
rect 85770 -149000 86570 -148990
rect 87270 -148915 88070 -148900
rect 87270 -148935 87280 -148915
rect 88060 -148935 88070 -148915
rect 87270 -148960 88070 -148935
rect 87270 -148990 87280 -148960
rect 88060 -148990 88070 -148960
rect 87270 -149000 88070 -148990
rect 88770 -148915 89570 -148900
rect 88770 -148935 88780 -148915
rect 89560 -148935 89570 -148915
rect 88770 -148960 89570 -148935
rect 88770 -148990 88780 -148960
rect 89560 -148990 89570 -148960
rect 88770 -149000 89570 -148990
rect 90270 -148915 91070 -148900
rect 90270 -148935 90280 -148915
rect 91060 -148935 91070 -148915
rect 90270 -148960 91070 -148935
rect 90270 -148990 90280 -148960
rect 91060 -148990 91070 -148960
rect 90270 -149000 91070 -148990
rect 91770 -148915 92570 -148900
rect 91770 -148935 91780 -148915
rect 92560 -148935 92570 -148915
rect 91770 -148960 92570 -148935
rect 91770 -148990 91780 -148960
rect 92560 -148990 92570 -148960
rect 91770 -149000 92570 -148990
rect 93270 -148915 94070 -148900
rect 93270 -148935 93280 -148915
rect 94060 -148935 94070 -148915
rect 93270 -148960 94070 -148935
rect 93270 -148990 93280 -148960
rect 94060 -148990 94070 -148960
rect 93270 -149000 94070 -148990
rect 94770 -148915 95570 -148900
rect 94770 -148935 94780 -148915
rect 95560 -148935 95570 -148915
rect 94770 -148960 95570 -148935
rect 94770 -148990 94780 -148960
rect 95560 -148990 95570 -148960
rect 94770 -149000 95570 -148990
rect 96270 -148915 97070 -148900
rect 96270 -148935 96280 -148915
rect 97060 -148935 97070 -148915
rect 96270 -148960 97070 -148935
rect 96270 -148990 96280 -148960
rect 97060 -148990 97070 -148960
rect 96270 -149000 97070 -148990
rect 97770 -148915 98570 -148900
rect 97770 -148935 97780 -148915
rect 98560 -148935 98570 -148915
rect 97770 -148960 98570 -148935
rect 97770 -148990 97780 -148960
rect 98560 -148990 98570 -148960
rect 97770 -149000 98570 -148990
rect 99270 -148915 100070 -148900
rect 99270 -148935 99280 -148915
rect 100060 -148935 100070 -148915
rect 99270 -148960 100070 -148935
rect 99270 -148990 99280 -148960
rect 100060 -148990 100070 -148960
rect 99270 -149000 100070 -148990
rect 100770 -148915 101570 -148900
rect 100770 -148935 100780 -148915
rect 101560 -148935 101570 -148915
rect 100770 -148960 101570 -148935
rect 100770 -148990 100780 -148960
rect 101560 -148990 101570 -148960
rect 100770 -149000 101570 -148990
rect 102270 -148915 103070 -148900
rect 102270 -148935 102280 -148915
rect 103060 -148935 103070 -148915
rect 102270 -148960 103070 -148935
rect 102270 -148990 102280 -148960
rect 103060 -148990 103070 -148960
rect 102270 -149000 103070 -148990
rect 103770 -148915 104570 -148900
rect 103770 -148935 103780 -148915
rect 104560 -148935 104570 -148915
rect 103770 -148960 104570 -148935
rect 103770 -148990 103780 -148960
rect 104560 -148990 104570 -148960
rect 103770 -149000 104570 -148990
rect 105270 -148915 106070 -148900
rect 105270 -148935 105280 -148915
rect 106060 -148935 106070 -148915
rect 105270 -148960 106070 -148935
rect 105270 -148990 105280 -148960
rect 106060 -148990 106070 -148960
rect 105270 -149000 106070 -148990
rect 106770 -148915 107570 -148900
rect 106770 -148935 106780 -148915
rect 107560 -148935 107570 -148915
rect 106770 -148960 107570 -148935
rect 106770 -148990 106780 -148960
rect 107560 -148990 107570 -148960
rect 106770 -149000 107570 -148990
rect 108270 -148915 109070 -148900
rect 108270 -148935 108280 -148915
rect 109060 -148935 109070 -148915
rect 108270 -148960 109070 -148935
rect 108270 -148990 108280 -148960
rect 109060 -148990 109070 -148960
rect 108270 -149000 109070 -148990
rect 109770 -148915 110570 -148900
rect 109770 -148935 109780 -148915
rect 110560 -148935 110570 -148915
rect 109770 -148960 110570 -148935
rect 109770 -148990 109780 -148960
rect 110560 -148990 110570 -148960
rect 109770 -149000 110570 -148990
rect 111270 -148915 112070 -148900
rect 111270 -148935 111280 -148915
rect 112060 -148935 112070 -148915
rect 111270 -148960 112070 -148935
rect 111270 -148990 111280 -148960
rect 112060 -148990 112070 -148960
rect 111270 -149000 112070 -148990
rect 112770 -148915 113570 -148900
rect 112770 -148935 112780 -148915
rect 113560 -148935 113570 -148915
rect 112770 -148960 113570 -148935
rect 112770 -148990 112780 -148960
rect 113560 -148990 113570 -148960
rect 112770 -149000 113570 -148990
rect 114270 -148915 115070 -148900
rect 114270 -148935 114280 -148915
rect 115060 -148935 115070 -148915
rect 114270 -148960 115070 -148935
rect 114270 -148990 114280 -148960
rect 115060 -148990 115070 -148960
rect 114270 -149000 115070 -148990
rect 115770 -148915 116570 -148900
rect 115770 -148935 115780 -148915
rect 116560 -148935 116570 -148915
rect 115770 -148960 116570 -148935
rect 115770 -148990 115780 -148960
rect 116560 -148990 116570 -148960
rect 115770 -149000 116570 -148990
rect 117270 -148915 118070 -148900
rect 117270 -148935 117280 -148915
rect 118060 -148935 118070 -148915
rect 117270 -148960 118070 -148935
rect 117270 -148990 117280 -148960
rect 118060 -148990 118070 -148960
rect 117270 -149000 118070 -148990
rect 118770 -148915 119570 -148900
rect 118770 -148935 118780 -148915
rect 119560 -148935 119570 -148915
rect 118770 -148960 119570 -148935
rect 118770 -148990 118780 -148960
rect 119560 -148990 119570 -148960
rect 118770 -149000 119570 -148990
rect 120270 -148915 121070 -148900
rect 120270 -148935 120280 -148915
rect 121060 -148935 121070 -148915
rect 120270 -148960 121070 -148935
rect 120270 -148990 120280 -148960
rect 121060 -148990 121070 -148960
rect 120270 -149000 121070 -148990
rect 121770 -148915 122570 -148900
rect 121770 -148935 121780 -148915
rect 122560 -148935 122570 -148915
rect 121770 -148960 122570 -148935
rect 121770 -148990 121780 -148960
rect 122560 -148990 122570 -148960
rect 121770 -149000 122570 -148990
rect 123270 -148915 124070 -148900
rect 123270 -148935 123280 -148915
rect 124060 -148935 124070 -148915
rect 123270 -148960 124070 -148935
rect 123270 -148990 123280 -148960
rect 124060 -148990 124070 -148960
rect 123270 -149000 124070 -148990
rect 124770 -148915 125570 -148900
rect 124770 -148935 124780 -148915
rect 125560 -148935 125570 -148915
rect 124770 -148960 125570 -148935
rect 124770 -148990 124780 -148960
rect 125560 -148990 125570 -148960
rect 124770 -149000 125570 -148990
rect 126270 -148915 127070 -148900
rect 126270 -148935 126280 -148915
rect 127060 -148935 127070 -148915
rect 126270 -148960 127070 -148935
rect 126270 -148990 126280 -148960
rect 127060 -148990 127070 -148960
rect 126270 -149000 127070 -148990
rect 127770 -148915 128570 -148900
rect 127770 -148935 127780 -148915
rect 128560 -148935 128570 -148915
rect 127770 -148960 128570 -148935
rect 127770 -148990 127780 -148960
rect 128560 -148990 128570 -148960
rect 127770 -149000 128570 -148990
rect 129270 -148915 130070 -148900
rect 129270 -148935 129280 -148915
rect 130060 -148935 130070 -148915
rect 129270 -148960 130070 -148935
rect 129270 -148990 129280 -148960
rect 130060 -148990 130070 -148960
rect 129270 -149000 130070 -148990
rect 130770 -148915 131570 -148900
rect 130770 -148935 130780 -148915
rect 131560 -148935 131570 -148915
rect 130770 -148960 131570 -148935
rect 130770 -148990 130780 -148960
rect 131560 -148990 131570 -148960
rect 130770 -149000 131570 -148990
rect 132270 -148915 133070 -148900
rect 132270 -148935 132280 -148915
rect 133060 -148935 133070 -148915
rect 132270 -148960 133070 -148935
rect 132270 -148990 132280 -148960
rect 133060 -148990 133070 -148960
rect 132270 -149000 133070 -148990
rect 133770 -148915 134570 -148900
rect 133770 -148935 133780 -148915
rect 134560 -148935 134570 -148915
rect 133770 -148960 134570 -148935
rect 133770 -148990 133780 -148960
rect 134560 -148990 134570 -148960
rect 133770 -149000 134570 -148990
rect 135270 -148915 136070 -148900
rect 135270 -148935 135280 -148915
rect 136060 -148935 136070 -148915
rect 135270 -148960 136070 -148935
rect 135270 -148990 135280 -148960
rect 136060 -148990 136070 -148960
rect 135270 -149000 136070 -148990
rect 136770 -148915 137570 -148900
rect 136770 -148935 136780 -148915
rect 137560 -148935 137570 -148915
rect 136770 -148960 137570 -148935
rect 136770 -148990 136780 -148960
rect 137560 -148990 137570 -148960
rect 136770 -149000 137570 -148990
rect 138270 -148915 139070 -148900
rect 138270 -148935 138280 -148915
rect 139060 -148935 139070 -148915
rect 138270 -148960 139070 -148935
rect 138270 -148990 138280 -148960
rect 139060 -148990 139070 -148960
rect 138270 -149000 139070 -148990
rect 139770 -148915 140570 -148900
rect 139770 -148935 139780 -148915
rect 140560 -148935 140570 -148915
rect 139770 -148960 140570 -148935
rect 139770 -148990 139780 -148960
rect 140560 -148990 140570 -148960
rect 139770 -149000 140570 -148990
rect 141270 -148915 142070 -148900
rect 141270 -148935 141280 -148915
rect 142060 -148935 142070 -148915
rect 141270 -148960 142070 -148935
rect 141270 -148990 141280 -148960
rect 142060 -148990 142070 -148960
rect 141270 -149000 142070 -148990
rect 142770 -148915 143570 -148900
rect 142770 -148935 142780 -148915
rect 143560 -148935 143570 -148915
rect 142770 -148960 143570 -148935
rect 142770 -148990 142780 -148960
rect 143560 -148990 143570 -148960
rect 142770 -149000 143570 -148990
rect 144270 -148915 145070 -148900
rect 144270 -148935 144280 -148915
rect 145060 -148935 145070 -148915
rect 144270 -148960 145070 -148935
rect 144270 -148990 144280 -148960
rect 145060 -148990 145070 -148960
rect 144270 -149000 145070 -148990
rect 145770 -148915 146570 -148900
rect 145770 -148935 145780 -148915
rect 146560 -148935 146570 -148915
rect 145770 -148960 146570 -148935
rect 145770 -148990 145780 -148960
rect 146560 -148990 146570 -148960
rect 145770 -149000 146570 -148990
rect 147270 -148915 148070 -148900
rect 147270 -148935 147280 -148915
rect 148060 -148935 148070 -148915
rect 147270 -148960 148070 -148935
rect 147270 -148990 147280 -148960
rect 148060 -148990 148070 -148960
rect 147270 -149000 148070 -148990
rect 148770 -148915 149570 -148900
rect 148770 -148935 148780 -148915
rect 149560 -148935 149570 -148915
rect 148770 -148960 149570 -148935
rect 148770 -148990 148780 -148960
rect 149560 -148990 149570 -148960
rect 148770 -149000 149570 -148990
<< viali >>
rect 280 -148645 1060 -148615
rect 1780 -148645 2560 -148615
rect 3280 -148645 4060 -148615
rect 4780 -148645 5560 -148615
rect 6280 -148645 7060 -148615
rect 7780 -148645 8560 -148615
rect 9280 -148645 10060 -148615
rect 10780 -148645 11560 -148615
rect 12280 -148645 13060 -148615
rect 13780 -148645 14560 -148615
rect 15280 -148645 16060 -148615
rect 16780 -148645 17560 -148615
rect 18280 -148645 19060 -148615
rect 19780 -148645 20560 -148615
rect 21280 -148645 22060 -148615
rect 22780 -148645 23560 -148615
rect 24280 -148645 25060 -148615
rect 25780 -148645 26560 -148615
rect 27280 -148645 28060 -148615
rect 28780 -148645 29560 -148615
rect 30280 -148645 31060 -148615
rect 31780 -148645 32560 -148615
rect 33280 -148645 34060 -148615
rect 34780 -148645 35560 -148615
rect 36280 -148645 37060 -148615
rect 37780 -148645 38560 -148615
rect 39280 -148645 40060 -148615
rect 40780 -148645 41560 -148615
rect 42280 -148645 43060 -148615
rect 43780 -148645 44560 -148615
rect 45280 -148645 46060 -148615
rect 46780 -148645 47560 -148615
rect 48280 -148645 49060 -148615
rect 49780 -148645 50560 -148615
rect 51280 -148645 52060 -148615
rect 52780 -148645 53560 -148615
rect 54280 -148645 55060 -148615
rect 55780 -148645 56560 -148615
rect 57280 -148645 58060 -148615
rect 58780 -148645 59560 -148615
rect 60280 -148645 61060 -148615
rect 61780 -148645 62560 -148615
rect 63280 -148645 64060 -148615
rect 64780 -148645 65560 -148615
rect 66280 -148645 67060 -148615
rect 67780 -148645 68560 -148615
rect 69280 -148645 70060 -148615
rect 70780 -148645 71560 -148615
rect 72280 -148645 73060 -148615
rect 73780 -148645 74560 -148615
rect 75280 -148645 76060 -148615
rect 76780 -148645 77560 -148615
rect 78280 -148645 79060 -148615
rect 79780 -148645 80560 -148615
rect 81280 -148645 82060 -148615
rect 82780 -148645 83560 -148615
rect 84280 -148645 85060 -148615
rect 85780 -148645 86560 -148615
rect 87280 -148645 88060 -148615
rect 88780 -148645 89560 -148615
rect 90280 -148645 91060 -148615
rect 91780 -148645 92560 -148615
rect 93280 -148645 94060 -148615
rect 94780 -148645 95560 -148615
rect 96280 -148645 97060 -148615
rect 97780 -148645 98560 -148615
rect 99280 -148645 100060 -148615
rect 100780 -148645 101560 -148615
rect 102280 -148645 103060 -148615
rect 103780 -148645 104560 -148615
rect 105280 -148645 106060 -148615
rect 106780 -148645 107560 -148615
rect 108280 -148645 109060 -148615
rect 109780 -148645 110560 -148615
rect 111280 -148645 112060 -148615
rect 112780 -148645 113560 -148615
rect 114280 -148645 115060 -148615
rect 115780 -148645 116560 -148615
rect 117280 -148645 118060 -148615
rect 118780 -148645 119560 -148615
rect 120280 -148645 121060 -148615
rect 121780 -148645 122560 -148615
rect 123280 -148645 124060 -148615
rect 124780 -148645 125560 -148615
rect 126280 -148645 127060 -148615
rect 127780 -148645 128560 -148615
rect 129280 -148645 130060 -148615
rect 130780 -148645 131560 -148615
rect 132280 -148645 133060 -148615
rect 133780 -148645 134560 -148615
rect 135280 -148645 136060 -148615
rect 136780 -148645 137560 -148615
rect 138280 -148645 139060 -148615
rect 139780 -148645 140560 -148615
rect 141280 -148645 142060 -148615
rect 142780 -148645 143560 -148615
rect 144280 -148645 145060 -148615
rect 145780 -148645 146560 -148615
rect 147280 -148645 148060 -148615
rect 148780 -148645 149560 -148615
rect 120 -148850 210 -148750
rect 1620 -148850 1710 -148750
rect 3120 -148850 3210 -148750
rect 4620 -148850 4710 -148750
rect 6120 -148850 6210 -148750
rect 7620 -148850 7710 -148750
rect 9120 -148850 9210 -148750
rect 10620 -148850 10710 -148750
rect 12120 -148850 12210 -148750
rect 13620 -148850 13710 -148750
rect 15120 -148850 15210 -148750
rect 16620 -148850 16710 -148750
rect 18120 -148850 18210 -148750
rect 19620 -148850 19710 -148750
rect 21120 -148850 21210 -148750
rect 22620 -148850 22710 -148750
rect 24120 -148850 24210 -148750
rect 25620 -148850 25710 -148750
rect 27120 -148850 27210 -148750
rect 28620 -148850 28710 -148750
rect 30120 -148850 30210 -148750
rect 31620 -148850 31710 -148750
rect 33120 -148850 33210 -148750
rect 34620 -148850 34710 -148750
rect 36120 -148850 36210 -148750
rect 37620 -148850 37710 -148750
rect 39120 -148850 39210 -148750
rect 40620 -148850 40710 -148750
rect 42120 -148850 42210 -148750
rect 43620 -148850 43710 -148750
rect 45120 -148850 45210 -148750
rect 46620 -148850 46710 -148750
rect 48120 -148850 48210 -148750
rect 49620 -148850 49710 -148750
rect 51120 -148850 51210 -148750
rect 52620 -148850 52710 -148750
rect 54120 -148850 54210 -148750
rect 55620 -148850 55710 -148750
rect 57120 -148850 57210 -148750
rect 58620 -148850 58710 -148750
rect 60120 -148850 60210 -148750
rect 61620 -148850 61710 -148750
rect 63120 -148850 63210 -148750
rect 64620 -148850 64710 -148750
rect 66120 -148850 66210 -148750
rect 67620 -148850 67710 -148750
rect 69120 -148850 69210 -148750
rect 70620 -148850 70710 -148750
rect 72120 -148850 72210 -148750
rect 73620 -148850 73710 -148750
rect 75120 -148850 75210 -148750
rect 76620 -148850 76710 -148750
rect 78120 -148850 78210 -148750
rect 79620 -148850 79710 -148750
rect 81120 -148850 81210 -148750
rect 82620 -148850 82710 -148750
rect 84120 -148850 84210 -148750
rect 85620 -148850 85710 -148750
rect 87120 -148850 87210 -148750
rect 88620 -148850 88710 -148750
rect 90120 -148850 90210 -148750
rect 91620 -148850 91710 -148750
rect 93120 -148850 93210 -148750
rect 94620 -148850 94710 -148750
rect 96120 -148850 96210 -148750
rect 97620 -148850 97710 -148750
rect 99120 -148850 99210 -148750
rect 100620 -148850 100710 -148750
rect 102120 -148850 102210 -148750
rect 103620 -148850 103710 -148750
rect 105120 -148850 105210 -148750
rect 106620 -148850 106710 -148750
rect 108120 -148850 108210 -148750
rect 109620 -148850 109710 -148750
rect 111120 -148850 111210 -148750
rect 112620 -148850 112710 -148750
rect 114120 -148850 114210 -148750
rect 115620 -148850 115710 -148750
rect 117120 -148850 117210 -148750
rect 118620 -148850 118710 -148750
rect 120120 -148850 120210 -148750
rect 121620 -148850 121710 -148750
rect 123120 -148850 123210 -148750
rect 124620 -148850 124710 -148750
rect 126120 -148850 126210 -148750
rect 127620 -148850 127710 -148750
rect 129120 -148850 129210 -148750
rect 130620 -148850 130710 -148750
rect 132120 -148850 132210 -148750
rect 133620 -148850 133710 -148750
rect 135120 -148850 135210 -148750
rect 136620 -148850 136710 -148750
rect 138120 -148850 138210 -148750
rect 139620 -148850 139710 -148750
rect 141120 -148850 141210 -148750
rect 142620 -148850 142710 -148750
rect 144120 -148850 144210 -148750
rect 145620 -148850 145710 -148750
rect 147120 -148850 147210 -148750
rect 148620 -148850 148710 -148750
rect 280 -148990 1060 -148960
rect 1780 -148990 2560 -148960
rect 3280 -148990 4060 -148960
rect 4780 -148990 5560 -148960
rect 6280 -148990 7060 -148960
rect 7780 -148990 8560 -148960
rect 9280 -148990 10060 -148960
rect 10780 -148990 11560 -148960
rect 12280 -148990 13060 -148960
rect 13780 -148990 14560 -148960
rect 15280 -148990 16060 -148960
rect 16780 -148990 17560 -148960
rect 18280 -148990 19060 -148960
rect 19780 -148990 20560 -148960
rect 21280 -148990 22060 -148960
rect 22780 -148990 23560 -148960
rect 24280 -148990 25060 -148960
rect 25780 -148990 26560 -148960
rect 27280 -148990 28060 -148960
rect 28780 -148990 29560 -148960
rect 30280 -148990 31060 -148960
rect 31780 -148990 32560 -148960
rect 33280 -148990 34060 -148960
rect 34780 -148990 35560 -148960
rect 36280 -148990 37060 -148960
rect 37780 -148990 38560 -148960
rect 39280 -148990 40060 -148960
rect 40780 -148990 41560 -148960
rect 42280 -148990 43060 -148960
rect 43780 -148990 44560 -148960
rect 45280 -148990 46060 -148960
rect 46780 -148990 47560 -148960
rect 48280 -148990 49060 -148960
rect 49780 -148990 50560 -148960
rect 51280 -148990 52060 -148960
rect 52780 -148990 53560 -148960
rect 54280 -148990 55060 -148960
rect 55780 -148990 56560 -148960
rect 57280 -148990 58060 -148960
rect 58780 -148990 59560 -148960
rect 60280 -148990 61060 -148960
rect 61780 -148990 62560 -148960
rect 63280 -148990 64060 -148960
rect 64780 -148990 65560 -148960
rect 66280 -148990 67060 -148960
rect 67780 -148990 68560 -148960
rect 69280 -148990 70060 -148960
rect 70780 -148990 71560 -148960
rect 72280 -148990 73060 -148960
rect 73780 -148990 74560 -148960
rect 75280 -148990 76060 -148960
rect 76780 -148990 77560 -148960
rect 78280 -148990 79060 -148960
rect 79780 -148990 80560 -148960
rect 81280 -148990 82060 -148960
rect 82780 -148990 83560 -148960
rect 84280 -148990 85060 -148960
rect 85780 -148990 86560 -148960
rect 87280 -148990 88060 -148960
rect 88780 -148990 89560 -148960
rect 90280 -148990 91060 -148960
rect 91780 -148990 92560 -148960
rect 93280 -148990 94060 -148960
rect 94780 -148990 95560 -148960
rect 96280 -148990 97060 -148960
rect 97780 -148990 98560 -148960
rect 99280 -148990 100060 -148960
rect 100780 -148990 101560 -148960
rect 102280 -148990 103060 -148960
rect 103780 -148990 104560 -148960
rect 105280 -148990 106060 -148960
rect 106780 -148990 107560 -148960
rect 108280 -148990 109060 -148960
rect 109780 -148990 110560 -148960
rect 111280 -148990 112060 -148960
rect 112780 -148990 113560 -148960
rect 114280 -148990 115060 -148960
rect 115780 -148990 116560 -148960
rect 117280 -148990 118060 -148960
rect 118780 -148990 119560 -148960
rect 120280 -148990 121060 -148960
rect 121780 -148990 122560 -148960
rect 123280 -148990 124060 -148960
rect 124780 -148990 125560 -148960
rect 126280 -148990 127060 -148960
rect 127780 -148990 128560 -148960
rect 129280 -148990 130060 -148960
rect 130780 -148990 131560 -148960
rect 132280 -148990 133060 -148960
rect 133780 -148990 134560 -148960
rect 135280 -148990 136060 -148960
rect 136780 -148990 137560 -148960
rect 138280 -148990 139060 -148960
rect 139780 -148990 140560 -148960
rect 141280 -148990 142060 -148960
rect 142780 -148990 143560 -148960
rect 144280 -148990 145060 -148960
rect 145780 -148990 146560 -148960
rect 147280 -148990 148060 -148960
rect 148780 -148990 149560 -148960
<< metal1 >>
rect -970 1725 149500 1730
rect -970 1680 -960 1725
rect -450 1680 25 1725
rect 70 1680 1525 1725
rect 1570 1680 3025 1725
rect 3070 1680 4525 1725
rect 4570 1680 6025 1725
rect 6070 1680 7525 1725
rect 7570 1680 9025 1725
rect 9070 1680 10525 1725
rect 10570 1680 12025 1725
rect 12070 1680 13525 1725
rect 13570 1680 15025 1725
rect 15070 1680 16525 1725
rect 16570 1680 18025 1725
rect 18070 1680 19525 1725
rect 19570 1680 21025 1725
rect 21070 1680 22525 1725
rect 22570 1680 24025 1725
rect 24070 1680 25525 1725
rect 25570 1680 27025 1725
rect 27070 1680 28525 1725
rect 28570 1680 30025 1725
rect 30070 1680 31525 1725
rect 31570 1680 33025 1725
rect 33070 1680 34525 1725
rect 34570 1680 36025 1725
rect 36070 1680 37525 1725
rect 37570 1680 39025 1725
rect 39070 1680 40525 1725
rect 40570 1680 42025 1725
rect 42070 1680 43525 1725
rect 43570 1680 45025 1725
rect 45070 1680 46525 1725
rect 46570 1680 48025 1725
rect 48070 1680 49525 1725
rect 49570 1680 51025 1725
rect 51070 1680 52525 1725
rect 52570 1680 54025 1725
rect 54070 1680 55525 1725
rect 55570 1680 57025 1725
rect 57070 1680 58525 1725
rect 58570 1680 60025 1725
rect 60070 1680 61525 1725
rect 61570 1680 63025 1725
rect 63070 1680 64525 1725
rect 64570 1680 66025 1725
rect 66070 1680 67525 1725
rect 67570 1680 69025 1725
rect 69070 1680 70525 1725
rect 70570 1680 72025 1725
rect 72070 1680 73525 1725
rect 73570 1680 75025 1725
rect 75070 1680 76525 1725
rect 76570 1680 78025 1725
rect 78070 1680 79525 1725
rect 79570 1680 81025 1725
rect 81070 1680 82525 1725
rect 82570 1680 84025 1725
rect 84070 1680 85525 1725
rect 85570 1680 87025 1725
rect 87070 1680 88525 1725
rect 88570 1680 90025 1725
rect 90070 1680 91525 1725
rect 91570 1680 93025 1725
rect 93070 1680 94525 1725
rect 94570 1680 96025 1725
rect 96070 1680 97525 1725
rect 97570 1680 99025 1725
rect 99070 1680 100525 1725
rect 100570 1680 102025 1725
rect 102070 1680 103525 1725
rect 103570 1680 105025 1725
rect 105070 1680 106525 1725
rect 106570 1680 108025 1725
rect 108070 1680 109525 1725
rect 109570 1680 111025 1725
rect 111070 1680 112525 1725
rect 112570 1680 114025 1725
rect 114070 1680 115525 1725
rect 115570 1680 117025 1725
rect 117070 1680 118525 1725
rect 118570 1680 120025 1725
rect 120070 1680 121525 1725
rect 121570 1680 123025 1725
rect 123070 1680 124525 1725
rect 124570 1680 126025 1725
rect 126070 1680 127525 1725
rect 127570 1680 129025 1725
rect 129070 1680 130525 1725
rect 130570 1680 132025 1725
rect 132070 1680 133525 1725
rect 133570 1680 135025 1725
rect 135070 1680 136525 1725
rect 136570 1680 138025 1725
rect 138070 1680 139525 1725
rect 139570 1680 141025 1725
rect 141070 1680 142525 1725
rect 142570 1680 144025 1725
rect 144070 1680 145525 1725
rect 145570 1680 147025 1725
rect 147070 1680 148525 1725
rect 148570 1680 149500 1725
rect -970 1675 149500 1680
rect -1000 1485 -900 1500
rect -1000 1410 0 1485
rect -1000 -15 -900 1410
rect -800 780 0 785
rect -800 745 -790 780
rect -590 745 -270 780
rect -130 745 0 780
rect -800 740 0 745
rect 150200 90 150300 1515
rect 150000 15 150300 90
rect -1000 -90 0 -15
rect -1000 -1515 -900 -90
rect -800 -720 0 -715
rect -800 -755 -790 -720
rect -590 -755 -270 -720
rect -130 -755 0 -720
rect -800 -760 0 -755
rect 150200 -1410 150300 15
rect 150000 -1485 150300 -1410
rect -1000 -1590 0 -1515
rect -1000 -3015 -900 -1590
rect -800 -2220 0 -2215
rect -800 -2255 -790 -2220
rect -590 -2255 -270 -2220
rect -130 -2255 0 -2220
rect -800 -2260 0 -2255
rect 150200 -2910 150300 -1485
rect 150000 -2985 150300 -2910
rect -1000 -3090 0 -3015
rect -1000 -4515 -900 -3090
rect -800 -3720 0 -3715
rect -800 -3755 -790 -3720
rect -590 -3755 -270 -3720
rect -130 -3755 0 -3720
rect -800 -3760 0 -3755
rect 150200 -4410 150300 -2985
rect 150000 -4485 150300 -4410
rect -1000 -4590 0 -4515
rect -1000 -6015 -900 -4590
rect -800 -5220 0 -5215
rect -800 -5255 -790 -5220
rect -590 -5255 -270 -5220
rect -130 -5255 0 -5220
rect -800 -5260 0 -5255
rect 150200 -5910 150300 -4485
rect 150000 -5985 150300 -5910
rect -1000 -6090 0 -6015
rect -1000 -7515 -900 -6090
rect -800 -6720 0 -6715
rect -800 -6755 -790 -6720
rect -590 -6755 -270 -6720
rect -130 -6755 0 -6720
rect -800 -6760 0 -6755
rect 150200 -7410 150300 -5985
rect 150000 -7485 150300 -7410
rect -1000 -7590 0 -7515
rect -1000 -9015 -900 -7590
rect -800 -8220 0 -8215
rect -800 -8255 -790 -8220
rect -590 -8255 -270 -8220
rect -130 -8255 0 -8220
rect -800 -8260 0 -8255
rect 150200 -8910 150300 -7485
rect 150000 -8985 150300 -8910
rect -1000 -9090 0 -9015
rect -1000 -10515 -900 -9090
rect -800 -9720 0 -9715
rect -800 -9755 -790 -9720
rect -590 -9755 -270 -9720
rect -130 -9755 0 -9720
rect -800 -9760 0 -9755
rect 150200 -10410 150300 -8985
rect 150000 -10485 150300 -10410
rect -1000 -10590 0 -10515
rect -1000 -12015 -900 -10590
rect -800 -11220 0 -11215
rect -800 -11255 -790 -11220
rect -590 -11255 -270 -11220
rect -130 -11255 0 -11220
rect -800 -11260 0 -11255
rect 150200 -11910 150300 -10485
rect 150000 -11985 150300 -11910
rect -1000 -12090 0 -12015
rect -1000 -13515 -900 -12090
rect -800 -12720 0 -12715
rect -800 -12755 -790 -12720
rect -590 -12755 -270 -12720
rect -130 -12755 0 -12720
rect -800 -12760 0 -12755
rect 150200 -13410 150300 -11985
rect 150000 -13485 150300 -13410
rect -1000 -13590 0 -13515
rect -1000 -15015 -900 -13590
rect -800 -14220 0 -14215
rect -800 -14255 -790 -14220
rect -590 -14255 -270 -14220
rect -130 -14255 0 -14220
rect -800 -14260 0 -14255
rect 150200 -14910 150300 -13485
rect 150000 -14985 150300 -14910
rect -1000 -15090 0 -15015
rect -1000 -16515 -900 -15090
rect -800 -15720 0 -15715
rect -800 -15755 -790 -15720
rect -590 -15755 -270 -15720
rect -130 -15755 0 -15720
rect -800 -15760 0 -15755
rect 150200 -16410 150300 -14985
rect 150000 -16485 150300 -16410
rect -1000 -16590 0 -16515
rect -1000 -18015 -900 -16590
rect -800 -17220 0 -17215
rect -800 -17255 -790 -17220
rect -590 -17255 -270 -17220
rect -130 -17255 0 -17220
rect -800 -17260 0 -17255
rect 150200 -17910 150300 -16485
rect 150000 -17985 150300 -17910
rect -1000 -18090 0 -18015
rect -1000 -19515 -900 -18090
rect -800 -18720 0 -18715
rect -800 -18755 -790 -18720
rect -590 -18755 -270 -18720
rect -130 -18755 0 -18720
rect -800 -18760 0 -18755
rect 150200 -19410 150300 -17985
rect 150000 -19485 150300 -19410
rect -1000 -19590 0 -19515
rect -1000 -21015 -900 -19590
rect -800 -20220 0 -20215
rect -800 -20255 -790 -20220
rect -590 -20255 -270 -20220
rect -130 -20255 0 -20220
rect -800 -20260 0 -20255
rect 150200 -20910 150300 -19485
rect 150000 -20985 150300 -20910
rect -1000 -21090 0 -21015
rect -1000 -22515 -900 -21090
rect -800 -21720 0 -21715
rect -800 -21755 -790 -21720
rect -590 -21755 -270 -21720
rect -130 -21755 0 -21720
rect -800 -21760 0 -21755
rect 150200 -22410 150300 -20985
rect 150000 -22485 150300 -22410
rect -1000 -22590 0 -22515
rect -1000 -24015 -900 -22590
rect -800 -23220 0 -23215
rect -800 -23255 -790 -23220
rect -590 -23255 -270 -23220
rect -130 -23255 0 -23220
rect -800 -23260 0 -23255
rect 150200 -23910 150300 -22485
rect 150000 -23985 150300 -23910
rect -1000 -24090 0 -24015
rect -1000 -25515 -900 -24090
rect -800 -24720 0 -24715
rect -800 -24755 -790 -24720
rect -590 -24755 -270 -24720
rect -130 -24755 0 -24720
rect -800 -24760 0 -24755
rect 150200 -25410 150300 -23985
rect 150000 -25485 150300 -25410
rect -1000 -25590 0 -25515
rect -1000 -27015 -900 -25590
rect -800 -26220 0 -26215
rect -800 -26255 -790 -26220
rect -590 -26255 -270 -26220
rect -130 -26255 0 -26220
rect -800 -26260 0 -26255
rect 150200 -26910 150300 -25485
rect 150000 -26985 150300 -26910
rect -1000 -27090 0 -27015
rect -1000 -28515 -900 -27090
rect -800 -27720 0 -27715
rect -800 -27755 -790 -27720
rect -590 -27755 -270 -27720
rect -130 -27755 0 -27720
rect -800 -27760 0 -27755
rect 150200 -28410 150300 -26985
rect 150000 -28485 150300 -28410
rect -1000 -28590 0 -28515
rect -1000 -30015 -900 -28590
rect -800 -29220 0 -29215
rect -800 -29255 -790 -29220
rect -590 -29255 -270 -29220
rect -130 -29255 0 -29220
rect -800 -29260 0 -29255
rect 150200 -29910 150300 -28485
rect 150000 -29985 150300 -29910
rect -1000 -30090 0 -30015
rect -1000 -31515 -900 -30090
rect -800 -30720 0 -30715
rect -800 -30755 -790 -30720
rect -590 -30755 -270 -30720
rect -130 -30755 0 -30720
rect -800 -30760 0 -30755
rect 150200 -31410 150300 -29985
rect 150000 -31485 150300 -31410
rect -1000 -31590 0 -31515
rect -1000 -33015 -900 -31590
rect -800 -32220 0 -32215
rect -800 -32255 -790 -32220
rect -590 -32255 -270 -32220
rect -130 -32255 0 -32220
rect -800 -32260 0 -32255
rect 150200 -32910 150300 -31485
rect 150000 -32985 150300 -32910
rect -1000 -33090 0 -33015
rect -1000 -34515 -900 -33090
rect -800 -33720 0 -33715
rect -800 -33755 -790 -33720
rect -590 -33755 -270 -33720
rect -130 -33755 0 -33720
rect -800 -33760 0 -33755
rect 150200 -34410 150300 -32985
rect 150000 -34485 150300 -34410
rect -1000 -34590 0 -34515
rect -1000 -36015 -900 -34590
rect -800 -35220 0 -35215
rect -800 -35255 -790 -35220
rect -590 -35255 -270 -35220
rect -130 -35255 0 -35220
rect -800 -35260 0 -35255
rect 150200 -35910 150300 -34485
rect 150000 -35985 150300 -35910
rect -1000 -36090 0 -36015
rect -1000 -37515 -900 -36090
rect -800 -36720 0 -36715
rect -800 -36755 -790 -36720
rect -590 -36755 -270 -36720
rect -130 -36755 0 -36720
rect -800 -36760 0 -36755
rect 150200 -37410 150300 -35985
rect 150000 -37485 150300 -37410
rect -1000 -37590 0 -37515
rect -1000 -39015 -900 -37590
rect -800 -38220 0 -38215
rect -800 -38255 -790 -38220
rect -590 -38255 -270 -38220
rect -130 -38255 0 -38220
rect -800 -38260 0 -38255
rect 150200 -38910 150300 -37485
rect 150000 -38985 150300 -38910
rect -1000 -39090 0 -39015
rect -1000 -40515 -900 -39090
rect -800 -39720 0 -39715
rect -800 -39755 -790 -39720
rect -590 -39755 -270 -39720
rect -130 -39755 0 -39720
rect -800 -39760 0 -39755
rect 150200 -40410 150300 -38985
rect 150000 -40485 150300 -40410
rect -1000 -40590 0 -40515
rect -1000 -42015 -900 -40590
rect -800 -41220 0 -41215
rect -800 -41255 -790 -41220
rect -590 -41255 -270 -41220
rect -130 -41255 0 -41220
rect -800 -41260 0 -41255
rect 150200 -41910 150300 -40485
rect 150000 -41985 150300 -41910
rect -1000 -42090 0 -42015
rect -1000 -43515 -900 -42090
rect -800 -42720 0 -42715
rect -800 -42755 -790 -42720
rect -590 -42755 -270 -42720
rect -130 -42755 0 -42720
rect -800 -42760 0 -42755
rect 150200 -43410 150300 -41985
rect 150000 -43485 150300 -43410
rect -1000 -43590 0 -43515
rect -1000 -45015 -900 -43590
rect -800 -44220 0 -44215
rect -800 -44255 -790 -44220
rect -590 -44255 -270 -44220
rect -130 -44255 0 -44220
rect -800 -44260 0 -44255
rect 150200 -44910 150300 -43485
rect 150000 -44985 150300 -44910
rect -1000 -45090 0 -45015
rect -1000 -46515 -900 -45090
rect -800 -45720 0 -45715
rect -800 -45755 -790 -45720
rect -590 -45755 -270 -45720
rect -130 -45755 0 -45720
rect -800 -45760 0 -45755
rect 150200 -46410 150300 -44985
rect 150000 -46485 150300 -46410
rect -1000 -46590 0 -46515
rect -1000 -48015 -900 -46590
rect -800 -47220 0 -47215
rect -800 -47255 -790 -47220
rect -590 -47255 -270 -47220
rect -130 -47255 0 -47220
rect -800 -47260 0 -47255
rect 150200 -47910 150300 -46485
rect 150000 -47985 150300 -47910
rect -1000 -48090 0 -48015
rect -1000 -49515 -900 -48090
rect -800 -48720 0 -48715
rect -800 -48755 -790 -48720
rect -590 -48755 -270 -48720
rect -130 -48755 0 -48720
rect -800 -48760 0 -48755
rect 150200 -49410 150300 -47985
rect 150000 -49485 150300 -49410
rect -1000 -49590 0 -49515
rect -1000 -51015 -900 -49590
rect -800 -50220 0 -50215
rect -800 -50255 -790 -50220
rect -590 -50255 -270 -50220
rect -130 -50255 0 -50220
rect -800 -50260 0 -50255
rect 150200 -50910 150300 -49485
rect 150000 -50985 150300 -50910
rect -1000 -51090 0 -51015
rect -1000 -52515 -900 -51090
rect -800 -51720 0 -51715
rect -800 -51755 -790 -51720
rect -590 -51755 -270 -51720
rect -130 -51755 0 -51720
rect -800 -51760 0 -51755
rect 150200 -52410 150300 -50985
rect 150000 -52485 150300 -52410
rect -1000 -52590 0 -52515
rect -1000 -54015 -900 -52590
rect -800 -53220 0 -53215
rect -800 -53255 -790 -53220
rect -590 -53255 -270 -53220
rect -130 -53255 0 -53220
rect -800 -53260 0 -53255
rect 150200 -53910 150300 -52485
rect 150000 -53985 150300 -53910
rect -1000 -54090 0 -54015
rect -1000 -55515 -900 -54090
rect -800 -54720 0 -54715
rect -800 -54755 -790 -54720
rect -590 -54755 -270 -54720
rect -130 -54755 0 -54720
rect -800 -54760 0 -54755
rect 150200 -55410 150300 -53985
rect 150000 -55485 150300 -55410
rect -1000 -55590 0 -55515
rect -1000 -57015 -900 -55590
rect -800 -56220 0 -56215
rect -800 -56255 -790 -56220
rect -590 -56255 -270 -56220
rect -130 -56255 0 -56220
rect -800 -56260 0 -56255
rect 150200 -56910 150300 -55485
rect 150000 -56985 150300 -56910
rect -1000 -57090 0 -57015
rect -1000 -58515 -900 -57090
rect -800 -57720 0 -57715
rect -800 -57755 -790 -57720
rect -590 -57755 -270 -57720
rect -130 -57755 0 -57720
rect -800 -57760 0 -57755
rect 150200 -58410 150300 -56985
rect 150000 -58485 150300 -58410
rect -1000 -58590 0 -58515
rect -1000 -60015 -900 -58590
rect -800 -59220 0 -59215
rect -800 -59255 -790 -59220
rect -590 -59255 -270 -59220
rect -130 -59255 0 -59220
rect -800 -59260 0 -59255
rect 150200 -59910 150300 -58485
rect 150000 -59985 150300 -59910
rect -1000 -60090 0 -60015
rect -1000 -61515 -900 -60090
rect -800 -60720 0 -60715
rect -800 -60755 -790 -60720
rect -590 -60755 -270 -60720
rect -130 -60755 0 -60720
rect -800 -60760 0 -60755
rect 150200 -61410 150300 -59985
rect 150000 -61485 150300 -61410
rect -1000 -61590 0 -61515
rect -1000 -63015 -900 -61590
rect -800 -62220 0 -62215
rect -800 -62255 -790 -62220
rect -590 -62255 -270 -62220
rect -130 -62255 0 -62220
rect -800 -62260 0 -62255
rect 150200 -62910 150300 -61485
rect 150000 -62985 150300 -62910
rect -1000 -63090 0 -63015
rect -1000 -64515 -900 -63090
rect -800 -63720 0 -63715
rect -800 -63755 -790 -63720
rect -590 -63755 -270 -63720
rect -130 -63755 0 -63720
rect -800 -63760 0 -63755
rect 150200 -64410 150300 -62985
rect 150000 -64485 150300 -64410
rect -1000 -64590 0 -64515
rect -1000 -66015 -900 -64590
rect -800 -65220 0 -65215
rect -800 -65255 -790 -65220
rect -590 -65255 -270 -65220
rect -130 -65255 0 -65220
rect -800 -65260 0 -65255
rect 150200 -65910 150300 -64485
rect 150000 -65985 150300 -65910
rect -1000 -66090 0 -66015
rect -1000 -67515 -900 -66090
rect -800 -66720 0 -66715
rect -800 -66755 -790 -66720
rect -590 -66755 -270 -66720
rect -130 -66755 0 -66720
rect -800 -66760 0 -66755
rect 150200 -67410 150300 -65985
rect 150000 -67485 150300 -67410
rect -1000 -67590 0 -67515
rect -1000 -69015 -900 -67590
rect -800 -68220 0 -68215
rect -800 -68255 -790 -68220
rect -590 -68255 -270 -68220
rect -130 -68255 0 -68220
rect -800 -68260 0 -68255
rect 150200 -68910 150300 -67485
rect 150000 -68985 150300 -68910
rect -1000 -69090 0 -69015
rect -1000 -70515 -900 -69090
rect -800 -69720 0 -69715
rect -800 -69755 -790 -69720
rect -590 -69755 -270 -69720
rect -130 -69755 0 -69720
rect -800 -69760 0 -69755
rect 150200 -70410 150300 -68985
rect 150000 -70485 150300 -70410
rect -1000 -70590 0 -70515
rect -1000 -72015 -900 -70590
rect -800 -71220 0 -71215
rect -800 -71255 -790 -71220
rect -590 -71255 -270 -71220
rect -130 -71255 0 -71220
rect -800 -71260 0 -71255
rect 150200 -71910 150300 -70485
rect 150000 -71985 150300 -71910
rect -1000 -72090 0 -72015
rect -1000 -73515 -900 -72090
rect -800 -72720 0 -72715
rect -800 -72755 -790 -72720
rect -590 -72755 -270 -72720
rect -130 -72755 0 -72720
rect -800 -72760 0 -72755
rect 150200 -73410 150300 -71985
rect 150000 -73485 150300 -73410
rect -1000 -73590 0 -73515
rect -1000 -75015 -900 -73590
rect -800 -74220 0 -74215
rect -800 -74255 -790 -74220
rect -590 -74255 -270 -74220
rect -130 -74255 0 -74220
rect -800 -74260 0 -74255
rect 150200 -74910 150300 -73485
rect 150000 -74985 150300 -74910
rect -1000 -75090 0 -75015
rect -1000 -76515 -900 -75090
rect -800 -75720 0 -75715
rect -800 -75755 -790 -75720
rect -590 -75755 -270 -75720
rect -130 -75755 0 -75720
rect -800 -75760 0 -75755
rect 150200 -76410 150300 -74985
rect 150000 -76485 150300 -76410
rect -1000 -76590 0 -76515
rect -1000 -78015 -900 -76590
rect -800 -77220 0 -77215
rect -800 -77255 -790 -77220
rect -590 -77255 -270 -77220
rect -130 -77255 0 -77220
rect -800 -77260 0 -77255
rect 150200 -77910 150300 -76485
rect 150000 -77985 150300 -77910
rect -1000 -78090 0 -78015
rect -1000 -79515 -900 -78090
rect -800 -78720 0 -78715
rect -800 -78755 -790 -78720
rect -590 -78755 -270 -78720
rect -130 -78755 0 -78720
rect -800 -78760 0 -78755
rect 150200 -79410 150300 -77985
rect 150000 -79485 150300 -79410
rect -1000 -79590 0 -79515
rect -1000 -81015 -900 -79590
rect -800 -80220 0 -80215
rect -800 -80255 -790 -80220
rect -590 -80255 -270 -80220
rect -130 -80255 0 -80220
rect -800 -80260 0 -80255
rect 150200 -80910 150300 -79485
rect 150000 -80985 150300 -80910
rect -1000 -81090 0 -81015
rect -1000 -82515 -900 -81090
rect -800 -81720 0 -81715
rect -800 -81755 -790 -81720
rect -590 -81755 -270 -81720
rect -130 -81755 0 -81720
rect -800 -81760 0 -81755
rect 150200 -82410 150300 -80985
rect 150000 -82485 150300 -82410
rect -1000 -82590 0 -82515
rect -1000 -84015 -900 -82590
rect -800 -83220 0 -83215
rect -800 -83255 -790 -83220
rect -590 -83255 -270 -83220
rect -130 -83255 0 -83220
rect -800 -83260 0 -83255
rect 150200 -83910 150300 -82485
rect 150000 -83985 150300 -83910
rect -1000 -84090 0 -84015
rect -1000 -85515 -900 -84090
rect -800 -84720 0 -84715
rect -800 -84755 -790 -84720
rect -590 -84755 -270 -84720
rect -130 -84755 0 -84720
rect -800 -84760 0 -84755
rect 150200 -85410 150300 -83985
rect 150000 -85485 150300 -85410
rect -1000 -85590 0 -85515
rect -1000 -87015 -900 -85590
rect -800 -86220 0 -86215
rect -800 -86255 -790 -86220
rect -590 -86255 -270 -86220
rect -130 -86255 0 -86220
rect -800 -86260 0 -86255
rect 150200 -86910 150300 -85485
rect 150000 -86985 150300 -86910
rect -1000 -87090 0 -87015
rect -1000 -88515 -900 -87090
rect -800 -87720 0 -87715
rect -800 -87755 -790 -87720
rect -590 -87755 -270 -87720
rect -130 -87755 0 -87720
rect -800 -87760 0 -87755
rect 150200 -88410 150300 -86985
rect 150000 -88485 150300 -88410
rect -1000 -88590 0 -88515
rect -1000 -90015 -900 -88590
rect -800 -89220 0 -89215
rect -800 -89255 -790 -89220
rect -590 -89255 -270 -89220
rect -130 -89255 0 -89220
rect -800 -89260 0 -89255
rect 150200 -89910 150300 -88485
rect 150000 -89985 150300 -89910
rect -1000 -90090 0 -90015
rect -1000 -91515 -900 -90090
rect -800 -90720 0 -90715
rect -800 -90755 -790 -90720
rect -590 -90755 -270 -90720
rect -130 -90755 0 -90720
rect -800 -90760 0 -90755
rect 150200 -91410 150300 -89985
rect 150000 -91485 150300 -91410
rect -1000 -91590 0 -91515
rect -1000 -93015 -900 -91590
rect -800 -92220 0 -92215
rect -800 -92255 -790 -92220
rect -590 -92255 -270 -92220
rect -130 -92255 0 -92220
rect -800 -92260 0 -92255
rect 150200 -92910 150300 -91485
rect 150000 -92985 150300 -92910
rect -1000 -93090 0 -93015
rect -1000 -94515 -900 -93090
rect -800 -93720 0 -93715
rect -800 -93755 -790 -93720
rect -590 -93755 -270 -93720
rect -130 -93755 0 -93720
rect -800 -93760 0 -93755
rect 150200 -94410 150300 -92985
rect 150000 -94485 150300 -94410
rect -1000 -94590 0 -94515
rect -1000 -96015 -900 -94590
rect -800 -95220 0 -95215
rect -800 -95255 -790 -95220
rect -590 -95255 -270 -95220
rect -130 -95255 0 -95220
rect -800 -95260 0 -95255
rect 150200 -95910 150300 -94485
rect 150000 -95985 150300 -95910
rect -1000 -96090 0 -96015
rect -1000 -97515 -900 -96090
rect -800 -96720 0 -96715
rect -800 -96755 -790 -96720
rect -590 -96755 -270 -96720
rect -130 -96755 0 -96720
rect -800 -96760 0 -96755
rect 150200 -97410 150300 -95985
rect 150000 -97485 150300 -97410
rect -1000 -97590 0 -97515
rect -1000 -99015 -900 -97590
rect -800 -98220 0 -98215
rect -800 -98255 -790 -98220
rect -590 -98255 -270 -98220
rect -130 -98255 0 -98220
rect -800 -98260 0 -98255
rect 150200 -98910 150300 -97485
rect 150000 -98985 150300 -98910
rect -1000 -99090 0 -99015
rect -1000 -100515 -900 -99090
rect -800 -99720 0 -99715
rect -800 -99755 -790 -99720
rect -590 -99755 -270 -99720
rect -130 -99755 0 -99720
rect -800 -99760 0 -99755
rect 150200 -100410 150300 -98985
rect 150000 -100485 150300 -100410
rect -1000 -100590 0 -100515
rect -1000 -102015 -900 -100590
rect -800 -101220 0 -101215
rect -800 -101255 -790 -101220
rect -590 -101255 -270 -101220
rect -130 -101255 0 -101220
rect -800 -101260 0 -101255
rect 150200 -101910 150300 -100485
rect 150000 -101985 150300 -101910
rect -1000 -102090 0 -102015
rect -1000 -103515 -900 -102090
rect -800 -102720 0 -102715
rect -800 -102755 -790 -102720
rect -590 -102755 -270 -102720
rect -130 -102755 0 -102720
rect -800 -102760 0 -102755
rect 150200 -103410 150300 -101985
rect 150000 -103485 150300 -103410
rect -1000 -103590 0 -103515
rect -1000 -105015 -900 -103590
rect -800 -104220 0 -104215
rect -800 -104255 -790 -104220
rect -590 -104255 -270 -104220
rect -130 -104255 0 -104220
rect -800 -104260 0 -104255
rect 150200 -104910 150300 -103485
rect 150000 -104985 150300 -104910
rect -1000 -105090 0 -105015
rect -1000 -106515 -900 -105090
rect -800 -105720 0 -105715
rect -800 -105755 -790 -105720
rect -590 -105755 -270 -105720
rect -130 -105755 0 -105720
rect -800 -105760 0 -105755
rect 150200 -106410 150300 -104985
rect 150000 -106485 150300 -106410
rect -1000 -106590 0 -106515
rect -1000 -108015 -900 -106590
rect -800 -107220 0 -107215
rect -800 -107255 -790 -107220
rect -590 -107255 -270 -107220
rect -130 -107255 0 -107220
rect -800 -107260 0 -107255
rect 150200 -107910 150300 -106485
rect 150000 -107985 150300 -107910
rect -1000 -108090 0 -108015
rect -1000 -109515 -900 -108090
rect -800 -108720 0 -108715
rect -800 -108755 -790 -108720
rect -590 -108755 -270 -108720
rect -130 -108755 0 -108720
rect -800 -108760 0 -108755
rect 150200 -109410 150300 -107985
rect 150000 -109485 150300 -109410
rect -1000 -109590 0 -109515
rect -1000 -111015 -900 -109590
rect -800 -110220 0 -110215
rect -800 -110255 -790 -110220
rect -590 -110255 -270 -110220
rect -130 -110255 0 -110220
rect -800 -110260 0 -110255
rect 150200 -110910 150300 -109485
rect 150000 -110985 150300 -110910
rect -1000 -111090 0 -111015
rect -1000 -112515 -900 -111090
rect -800 -111720 0 -111715
rect -800 -111755 -790 -111720
rect -590 -111755 -270 -111720
rect -130 -111755 0 -111720
rect -800 -111760 0 -111755
rect 150200 -112410 150300 -110985
rect 150000 -112485 150300 -112410
rect -1000 -112590 0 -112515
rect -1000 -114015 -900 -112590
rect -800 -113220 0 -113215
rect -800 -113255 -790 -113220
rect -590 -113255 -270 -113220
rect -130 -113255 0 -113220
rect -800 -113260 0 -113255
rect 150200 -113910 150300 -112485
rect 150000 -113985 150300 -113910
rect -1000 -114090 0 -114015
rect -1000 -115515 -900 -114090
rect -800 -114720 0 -114715
rect -800 -114755 -790 -114720
rect -590 -114755 -270 -114720
rect -130 -114755 0 -114720
rect -800 -114760 0 -114755
rect 150200 -115410 150300 -113985
rect 150000 -115485 150300 -115410
rect -1000 -115590 0 -115515
rect -1000 -117015 -900 -115590
rect -800 -116220 0 -116215
rect -800 -116255 -790 -116220
rect -590 -116255 -270 -116220
rect -130 -116255 0 -116220
rect -800 -116260 0 -116255
rect 150200 -116910 150300 -115485
rect 150000 -116985 150300 -116910
rect -1000 -117090 0 -117015
rect -1000 -118515 -900 -117090
rect -800 -117720 0 -117715
rect -800 -117755 -790 -117720
rect -590 -117755 -270 -117720
rect -130 -117755 0 -117720
rect -800 -117760 0 -117755
rect 150200 -118410 150300 -116985
rect 150000 -118485 150300 -118410
rect -1000 -118590 0 -118515
rect -1000 -120015 -900 -118590
rect -800 -119220 0 -119215
rect -800 -119255 -790 -119220
rect -590 -119255 -270 -119220
rect -130 -119255 0 -119220
rect -800 -119260 0 -119255
rect 150200 -119910 150300 -118485
rect 150000 -119985 150300 -119910
rect -1000 -120090 0 -120015
rect -1000 -121515 -900 -120090
rect -800 -120720 0 -120715
rect -800 -120755 -790 -120720
rect -590 -120755 -270 -120720
rect -130 -120755 0 -120720
rect -800 -120760 0 -120755
rect 150200 -121410 150300 -119985
rect 150000 -121485 150300 -121410
rect -1000 -121590 0 -121515
rect -1000 -123015 -900 -121590
rect -800 -122220 0 -122215
rect -800 -122255 -790 -122220
rect -590 -122255 -270 -122220
rect -130 -122255 0 -122220
rect -800 -122260 0 -122255
rect 150200 -122910 150300 -121485
rect 150000 -122985 150300 -122910
rect -1000 -123090 0 -123015
rect -1000 -124515 -900 -123090
rect -800 -123720 0 -123715
rect -800 -123755 -790 -123720
rect -590 -123755 -270 -123720
rect -130 -123755 0 -123720
rect -800 -123760 0 -123755
rect 150200 -124410 150300 -122985
rect 150000 -124485 150300 -124410
rect -1000 -124590 0 -124515
rect -1000 -126015 -900 -124590
rect -800 -125220 0 -125215
rect -800 -125255 -790 -125220
rect -590 -125255 -270 -125220
rect -130 -125255 0 -125220
rect -800 -125260 0 -125255
rect 150200 -125910 150300 -124485
rect 150000 -125985 150300 -125910
rect -1000 -126090 0 -126015
rect -1000 -127515 -900 -126090
rect -800 -126720 0 -126715
rect -800 -126755 -790 -126720
rect -590 -126755 -270 -126720
rect -130 -126755 0 -126720
rect -800 -126760 0 -126755
rect 150200 -127410 150300 -125985
rect 150000 -127485 150300 -127410
rect -1000 -127590 0 -127515
rect -1000 -129015 -900 -127590
rect -800 -128220 0 -128215
rect -800 -128255 -790 -128220
rect -590 -128255 -270 -128220
rect -130 -128255 0 -128220
rect -800 -128260 0 -128255
rect 150200 -128910 150300 -127485
rect 150000 -128985 150300 -128910
rect -1000 -129090 0 -129015
rect -1000 -130515 -900 -129090
rect -800 -129720 0 -129715
rect -800 -129755 -790 -129720
rect -590 -129755 -270 -129720
rect -130 -129755 0 -129720
rect -800 -129760 0 -129755
rect 150200 -130410 150300 -128985
rect 150000 -130485 150300 -130410
rect -1000 -130590 0 -130515
rect -1000 -132015 -900 -130590
rect -800 -131220 0 -131215
rect -800 -131255 -790 -131220
rect -590 -131255 -270 -131220
rect -130 -131255 0 -131220
rect -800 -131260 0 -131255
rect 150200 -131910 150300 -130485
rect 150000 -131985 150300 -131910
rect -1000 -132090 0 -132015
rect -1000 -133515 -900 -132090
rect -800 -132720 0 -132715
rect -800 -132755 -790 -132720
rect -590 -132755 -270 -132720
rect -130 -132755 0 -132720
rect -800 -132760 0 -132755
rect 150200 -133410 150300 -131985
rect 150000 -133485 150300 -133410
rect -1000 -133590 0 -133515
rect -1000 -135015 -900 -133590
rect -800 -134220 0 -134215
rect -800 -134255 -790 -134220
rect -590 -134255 -270 -134220
rect -130 -134255 0 -134220
rect -800 -134260 0 -134255
rect 150200 -134910 150300 -133485
rect 150000 -134985 150300 -134910
rect -1000 -135090 0 -135015
rect -1000 -136515 -900 -135090
rect -800 -135720 0 -135715
rect -800 -135755 -790 -135720
rect -590 -135755 -270 -135720
rect -130 -135755 0 -135720
rect -800 -135760 0 -135755
rect 150200 -136410 150300 -134985
rect 150000 -136485 150300 -136410
rect -1000 -136590 0 -136515
rect -1000 -138015 -900 -136590
rect -800 -137220 0 -137215
rect -800 -137255 -790 -137220
rect -590 -137255 -270 -137220
rect -130 -137255 0 -137220
rect -800 -137260 0 -137255
rect 150200 -137910 150300 -136485
rect 150000 -137985 150300 -137910
rect -1000 -138090 0 -138015
rect -1000 -139515 -900 -138090
rect -800 -138720 0 -138715
rect -800 -138755 -790 -138720
rect -590 -138755 -270 -138720
rect -130 -138755 0 -138720
rect -800 -138760 0 -138755
rect 150200 -139410 150300 -137985
rect 150000 -139485 150300 -139410
rect -1000 -139590 0 -139515
rect -1000 -141015 -900 -139590
rect -800 -140220 0 -140215
rect -800 -140255 -790 -140220
rect -590 -140255 -270 -140220
rect -130 -140255 0 -140220
rect -800 -140260 0 -140255
rect 150200 -140910 150300 -139485
rect 150000 -140985 150300 -140910
rect -1000 -141090 0 -141015
rect -1000 -142515 -900 -141090
rect -800 -141720 0 -141715
rect -800 -141755 -790 -141720
rect -590 -141755 -270 -141720
rect -130 -141755 0 -141720
rect -800 -141760 0 -141755
rect 150200 -142410 150300 -140985
rect 150000 -142485 150300 -142410
rect -1000 -142590 0 -142515
rect -1000 -144015 -900 -142590
rect -800 -143220 0 -143215
rect -800 -143255 -790 -143220
rect -590 -143255 -270 -143220
rect -130 -143255 0 -143220
rect -800 -143260 0 -143255
rect 150200 -143910 150300 -142485
rect 150000 -143985 150300 -143910
rect -1000 -144090 0 -144015
rect -1000 -145515 -900 -144090
rect -800 -144720 0 -144715
rect -800 -144755 -790 -144720
rect -590 -144755 -270 -144720
rect -130 -144755 0 -144720
rect -800 -144760 0 -144755
rect 150200 -145410 150300 -143985
rect 150000 -145485 150300 -145410
rect -1000 -145590 0 -145515
rect -1000 -147015 -900 -145590
rect -800 -146220 0 -146215
rect -800 -146255 -790 -146220
rect -590 -146255 -270 -146220
rect -130 -146255 0 -146220
rect -800 -146260 0 -146255
rect 150200 -146910 150300 -145485
rect 150000 -146985 150300 -146910
rect -1000 -147090 0 -147015
rect -1000 -148500 -900 -147090
rect -800 -147720 0 -147715
rect -800 -147755 -790 -147720
rect -590 -147755 -270 -147720
rect -130 -147755 0 -147720
rect -800 -147760 0 -147755
rect 150200 -148410 150300 -146985
rect 150000 -148485 150300 -148410
rect 270 -148600 280 -148565
rect 1060 -148600 1070 -148565
rect 270 -148615 1070 -148600
rect 270 -148645 280 -148615
rect 1060 -148645 1070 -148615
rect 270 -148650 1070 -148645
rect 1770 -148600 1780 -148565
rect 2560 -148600 2570 -148565
rect 1770 -148615 2570 -148600
rect 1770 -148645 1780 -148615
rect 2560 -148645 2570 -148615
rect 1770 -148650 2570 -148645
rect 3270 -148600 3280 -148565
rect 4060 -148600 4070 -148565
rect 3270 -148615 4070 -148600
rect 3270 -148645 3280 -148615
rect 4060 -148645 4070 -148615
rect 3270 -148650 4070 -148645
rect 4770 -148600 4780 -148565
rect 5560 -148600 5570 -148565
rect 4770 -148615 5570 -148600
rect 4770 -148645 4780 -148615
rect 5560 -148645 5570 -148615
rect 4770 -148650 5570 -148645
rect 6270 -148600 6280 -148565
rect 7060 -148600 7070 -148565
rect 6270 -148615 7070 -148600
rect 6270 -148645 6280 -148615
rect 7060 -148645 7070 -148615
rect 6270 -148650 7070 -148645
rect 7770 -148600 7780 -148565
rect 8560 -148600 8570 -148565
rect 7770 -148615 8570 -148600
rect 7770 -148645 7780 -148615
rect 8560 -148645 8570 -148615
rect 7770 -148650 8570 -148645
rect 9270 -148600 9280 -148565
rect 10060 -148600 10070 -148565
rect 9270 -148615 10070 -148600
rect 9270 -148645 9280 -148615
rect 10060 -148645 10070 -148615
rect 9270 -148650 10070 -148645
rect 10770 -148600 10780 -148565
rect 11560 -148600 11570 -148565
rect 10770 -148615 11570 -148600
rect 10770 -148645 10780 -148615
rect 11560 -148645 11570 -148615
rect 10770 -148650 11570 -148645
rect 12270 -148600 12280 -148565
rect 13060 -148600 13070 -148565
rect 12270 -148615 13070 -148600
rect 12270 -148645 12280 -148615
rect 13060 -148645 13070 -148615
rect 12270 -148650 13070 -148645
rect 13770 -148600 13780 -148565
rect 14560 -148600 14570 -148565
rect 13770 -148615 14570 -148600
rect 13770 -148645 13780 -148615
rect 14560 -148645 14570 -148615
rect 13770 -148650 14570 -148645
rect 15270 -148600 15280 -148565
rect 16060 -148600 16070 -148565
rect 15270 -148615 16070 -148600
rect 15270 -148645 15280 -148615
rect 16060 -148645 16070 -148615
rect 15270 -148650 16070 -148645
rect 16770 -148600 16780 -148565
rect 17560 -148600 17570 -148565
rect 16770 -148615 17570 -148600
rect 16770 -148645 16780 -148615
rect 17560 -148645 17570 -148615
rect 16770 -148650 17570 -148645
rect 18270 -148600 18280 -148565
rect 19060 -148600 19070 -148565
rect 18270 -148615 19070 -148600
rect 18270 -148645 18280 -148615
rect 19060 -148645 19070 -148615
rect 18270 -148650 19070 -148645
rect 19770 -148600 19780 -148565
rect 20560 -148600 20570 -148565
rect 19770 -148615 20570 -148600
rect 19770 -148645 19780 -148615
rect 20560 -148645 20570 -148615
rect 19770 -148650 20570 -148645
rect 21270 -148600 21280 -148565
rect 22060 -148600 22070 -148565
rect 21270 -148615 22070 -148600
rect 21270 -148645 21280 -148615
rect 22060 -148645 22070 -148615
rect 21270 -148650 22070 -148645
rect 22770 -148600 22780 -148565
rect 23560 -148600 23570 -148565
rect 22770 -148615 23570 -148600
rect 22770 -148645 22780 -148615
rect 23560 -148645 23570 -148615
rect 22770 -148650 23570 -148645
rect 24270 -148600 24280 -148565
rect 25060 -148600 25070 -148565
rect 24270 -148615 25070 -148600
rect 24270 -148645 24280 -148615
rect 25060 -148645 25070 -148615
rect 24270 -148650 25070 -148645
rect 25770 -148600 25780 -148565
rect 26560 -148600 26570 -148565
rect 25770 -148615 26570 -148600
rect 25770 -148645 25780 -148615
rect 26560 -148645 26570 -148615
rect 25770 -148650 26570 -148645
rect 27270 -148600 27280 -148565
rect 28060 -148600 28070 -148565
rect 27270 -148615 28070 -148600
rect 27270 -148645 27280 -148615
rect 28060 -148645 28070 -148615
rect 27270 -148650 28070 -148645
rect 28770 -148600 28780 -148565
rect 29560 -148600 29570 -148565
rect 28770 -148615 29570 -148600
rect 28770 -148645 28780 -148615
rect 29560 -148645 29570 -148615
rect 28770 -148650 29570 -148645
rect 30270 -148600 30280 -148565
rect 31060 -148600 31070 -148565
rect 30270 -148615 31070 -148600
rect 30270 -148645 30280 -148615
rect 31060 -148645 31070 -148615
rect 30270 -148650 31070 -148645
rect 31770 -148600 31780 -148565
rect 32560 -148600 32570 -148565
rect 31770 -148615 32570 -148600
rect 31770 -148645 31780 -148615
rect 32560 -148645 32570 -148615
rect 31770 -148650 32570 -148645
rect 33270 -148600 33280 -148565
rect 34060 -148600 34070 -148565
rect 33270 -148615 34070 -148600
rect 33270 -148645 33280 -148615
rect 34060 -148645 34070 -148615
rect 33270 -148650 34070 -148645
rect 34770 -148600 34780 -148565
rect 35560 -148600 35570 -148565
rect 34770 -148615 35570 -148600
rect 34770 -148645 34780 -148615
rect 35560 -148645 35570 -148615
rect 34770 -148650 35570 -148645
rect 36270 -148600 36280 -148565
rect 37060 -148600 37070 -148565
rect 36270 -148615 37070 -148600
rect 36270 -148645 36280 -148615
rect 37060 -148645 37070 -148615
rect 36270 -148650 37070 -148645
rect 37770 -148600 37780 -148565
rect 38560 -148600 38570 -148565
rect 37770 -148615 38570 -148600
rect 37770 -148645 37780 -148615
rect 38560 -148645 38570 -148615
rect 37770 -148650 38570 -148645
rect 39270 -148600 39280 -148565
rect 40060 -148600 40070 -148565
rect 39270 -148615 40070 -148600
rect 39270 -148645 39280 -148615
rect 40060 -148645 40070 -148615
rect 39270 -148650 40070 -148645
rect 40770 -148600 40780 -148565
rect 41560 -148600 41570 -148565
rect 40770 -148615 41570 -148600
rect 40770 -148645 40780 -148615
rect 41560 -148645 41570 -148615
rect 40770 -148650 41570 -148645
rect 42270 -148600 42280 -148565
rect 43060 -148600 43070 -148565
rect 42270 -148615 43070 -148600
rect 42270 -148645 42280 -148615
rect 43060 -148645 43070 -148615
rect 42270 -148650 43070 -148645
rect 43770 -148600 43780 -148565
rect 44560 -148600 44570 -148565
rect 43770 -148615 44570 -148600
rect 43770 -148645 43780 -148615
rect 44560 -148645 44570 -148615
rect 43770 -148650 44570 -148645
rect 45270 -148600 45280 -148565
rect 46060 -148600 46070 -148565
rect 45270 -148615 46070 -148600
rect 45270 -148645 45280 -148615
rect 46060 -148645 46070 -148615
rect 45270 -148650 46070 -148645
rect 46770 -148600 46780 -148565
rect 47560 -148600 47570 -148565
rect 46770 -148615 47570 -148600
rect 46770 -148645 46780 -148615
rect 47560 -148645 47570 -148615
rect 46770 -148650 47570 -148645
rect 48270 -148600 48280 -148565
rect 49060 -148600 49070 -148565
rect 48270 -148615 49070 -148600
rect 48270 -148645 48280 -148615
rect 49060 -148645 49070 -148615
rect 48270 -148650 49070 -148645
rect 49770 -148600 49780 -148565
rect 50560 -148600 50570 -148565
rect 49770 -148615 50570 -148600
rect 49770 -148645 49780 -148615
rect 50560 -148645 50570 -148615
rect 49770 -148650 50570 -148645
rect 51270 -148600 51280 -148565
rect 52060 -148600 52070 -148565
rect 51270 -148615 52070 -148600
rect 51270 -148645 51280 -148615
rect 52060 -148645 52070 -148615
rect 51270 -148650 52070 -148645
rect 52770 -148600 52780 -148565
rect 53560 -148600 53570 -148565
rect 52770 -148615 53570 -148600
rect 52770 -148645 52780 -148615
rect 53560 -148645 53570 -148615
rect 52770 -148650 53570 -148645
rect 54270 -148600 54280 -148565
rect 55060 -148600 55070 -148565
rect 54270 -148615 55070 -148600
rect 54270 -148645 54280 -148615
rect 55060 -148645 55070 -148615
rect 54270 -148650 55070 -148645
rect 55770 -148600 55780 -148565
rect 56560 -148600 56570 -148565
rect 55770 -148615 56570 -148600
rect 55770 -148645 55780 -148615
rect 56560 -148645 56570 -148615
rect 55770 -148650 56570 -148645
rect 57270 -148600 57280 -148565
rect 58060 -148600 58070 -148565
rect 57270 -148615 58070 -148600
rect 57270 -148645 57280 -148615
rect 58060 -148645 58070 -148615
rect 57270 -148650 58070 -148645
rect 58770 -148600 58780 -148565
rect 59560 -148600 59570 -148565
rect 58770 -148615 59570 -148600
rect 58770 -148645 58780 -148615
rect 59560 -148645 59570 -148615
rect 58770 -148650 59570 -148645
rect 60270 -148600 60280 -148565
rect 61060 -148600 61070 -148565
rect 60270 -148615 61070 -148600
rect 60270 -148645 60280 -148615
rect 61060 -148645 61070 -148615
rect 60270 -148650 61070 -148645
rect 61770 -148600 61780 -148565
rect 62560 -148600 62570 -148565
rect 61770 -148615 62570 -148600
rect 61770 -148645 61780 -148615
rect 62560 -148645 62570 -148615
rect 61770 -148650 62570 -148645
rect 63270 -148600 63280 -148565
rect 64060 -148600 64070 -148565
rect 63270 -148615 64070 -148600
rect 63270 -148645 63280 -148615
rect 64060 -148645 64070 -148615
rect 63270 -148650 64070 -148645
rect 64770 -148600 64780 -148565
rect 65560 -148600 65570 -148565
rect 64770 -148615 65570 -148600
rect 64770 -148645 64780 -148615
rect 65560 -148645 65570 -148615
rect 64770 -148650 65570 -148645
rect 66270 -148600 66280 -148565
rect 67060 -148600 67070 -148565
rect 66270 -148615 67070 -148600
rect 66270 -148645 66280 -148615
rect 67060 -148645 67070 -148615
rect 66270 -148650 67070 -148645
rect 67770 -148600 67780 -148565
rect 68560 -148600 68570 -148565
rect 67770 -148615 68570 -148600
rect 67770 -148645 67780 -148615
rect 68560 -148645 68570 -148615
rect 67770 -148650 68570 -148645
rect 69270 -148600 69280 -148565
rect 70060 -148600 70070 -148565
rect 69270 -148615 70070 -148600
rect 69270 -148645 69280 -148615
rect 70060 -148645 70070 -148615
rect 69270 -148650 70070 -148645
rect 70770 -148600 70780 -148565
rect 71560 -148600 71570 -148565
rect 70770 -148615 71570 -148600
rect 70770 -148645 70780 -148615
rect 71560 -148645 71570 -148615
rect 70770 -148650 71570 -148645
rect 72270 -148600 72280 -148565
rect 73060 -148600 73070 -148565
rect 72270 -148615 73070 -148600
rect 72270 -148645 72280 -148615
rect 73060 -148645 73070 -148615
rect 72270 -148650 73070 -148645
rect 73770 -148600 73780 -148565
rect 74560 -148600 74570 -148565
rect 73770 -148615 74570 -148600
rect 73770 -148645 73780 -148615
rect 74560 -148645 74570 -148615
rect 73770 -148650 74570 -148645
rect 75270 -148600 75280 -148565
rect 76060 -148600 76070 -148565
rect 75270 -148615 76070 -148600
rect 75270 -148645 75280 -148615
rect 76060 -148645 76070 -148615
rect 75270 -148650 76070 -148645
rect 76770 -148600 76780 -148565
rect 77560 -148600 77570 -148565
rect 76770 -148615 77570 -148600
rect 76770 -148645 76780 -148615
rect 77560 -148645 77570 -148615
rect 76770 -148650 77570 -148645
rect 78270 -148600 78280 -148565
rect 79060 -148600 79070 -148565
rect 78270 -148615 79070 -148600
rect 78270 -148645 78280 -148615
rect 79060 -148645 79070 -148615
rect 78270 -148650 79070 -148645
rect 79770 -148600 79780 -148565
rect 80560 -148600 80570 -148565
rect 79770 -148615 80570 -148600
rect 79770 -148645 79780 -148615
rect 80560 -148645 80570 -148615
rect 79770 -148650 80570 -148645
rect 81270 -148600 81280 -148565
rect 82060 -148600 82070 -148565
rect 81270 -148615 82070 -148600
rect 81270 -148645 81280 -148615
rect 82060 -148645 82070 -148615
rect 81270 -148650 82070 -148645
rect 82770 -148600 82780 -148565
rect 83560 -148600 83570 -148565
rect 82770 -148615 83570 -148600
rect 82770 -148645 82780 -148615
rect 83560 -148645 83570 -148615
rect 82770 -148650 83570 -148645
rect 84270 -148600 84280 -148565
rect 85060 -148600 85070 -148565
rect 84270 -148615 85070 -148600
rect 84270 -148645 84280 -148615
rect 85060 -148645 85070 -148615
rect 84270 -148650 85070 -148645
rect 85770 -148600 85780 -148565
rect 86560 -148600 86570 -148565
rect 85770 -148615 86570 -148600
rect 85770 -148645 85780 -148615
rect 86560 -148645 86570 -148615
rect 85770 -148650 86570 -148645
rect 87270 -148600 87280 -148565
rect 88060 -148600 88070 -148565
rect 87270 -148615 88070 -148600
rect 87270 -148645 87280 -148615
rect 88060 -148645 88070 -148615
rect 87270 -148650 88070 -148645
rect 88770 -148600 88780 -148565
rect 89560 -148600 89570 -148565
rect 88770 -148615 89570 -148600
rect 88770 -148645 88780 -148615
rect 89560 -148645 89570 -148615
rect 88770 -148650 89570 -148645
rect 90270 -148600 90280 -148565
rect 91060 -148600 91070 -148565
rect 90270 -148615 91070 -148600
rect 90270 -148645 90280 -148615
rect 91060 -148645 91070 -148615
rect 90270 -148650 91070 -148645
rect 91770 -148600 91780 -148565
rect 92560 -148600 92570 -148565
rect 91770 -148615 92570 -148600
rect 91770 -148645 91780 -148615
rect 92560 -148645 92570 -148615
rect 91770 -148650 92570 -148645
rect 93270 -148600 93280 -148565
rect 94060 -148600 94070 -148565
rect 93270 -148615 94070 -148600
rect 93270 -148645 93280 -148615
rect 94060 -148645 94070 -148615
rect 93270 -148650 94070 -148645
rect 94770 -148600 94780 -148565
rect 95560 -148600 95570 -148565
rect 94770 -148615 95570 -148600
rect 94770 -148645 94780 -148615
rect 95560 -148645 95570 -148615
rect 94770 -148650 95570 -148645
rect 96270 -148600 96280 -148565
rect 97060 -148600 97070 -148565
rect 96270 -148615 97070 -148600
rect 96270 -148645 96280 -148615
rect 97060 -148645 97070 -148615
rect 96270 -148650 97070 -148645
rect 97770 -148600 97780 -148565
rect 98560 -148600 98570 -148565
rect 97770 -148615 98570 -148600
rect 97770 -148645 97780 -148615
rect 98560 -148645 98570 -148615
rect 97770 -148650 98570 -148645
rect 99270 -148600 99280 -148565
rect 100060 -148600 100070 -148565
rect 99270 -148615 100070 -148600
rect 99270 -148645 99280 -148615
rect 100060 -148645 100070 -148615
rect 99270 -148650 100070 -148645
rect 100770 -148600 100780 -148565
rect 101560 -148600 101570 -148565
rect 100770 -148615 101570 -148600
rect 100770 -148645 100780 -148615
rect 101560 -148645 101570 -148615
rect 100770 -148650 101570 -148645
rect 102270 -148600 102280 -148565
rect 103060 -148600 103070 -148565
rect 102270 -148615 103070 -148600
rect 102270 -148645 102280 -148615
rect 103060 -148645 103070 -148615
rect 102270 -148650 103070 -148645
rect 103770 -148600 103780 -148565
rect 104560 -148600 104570 -148565
rect 103770 -148615 104570 -148600
rect 103770 -148645 103780 -148615
rect 104560 -148645 104570 -148615
rect 103770 -148650 104570 -148645
rect 105270 -148600 105280 -148565
rect 106060 -148600 106070 -148565
rect 105270 -148615 106070 -148600
rect 105270 -148645 105280 -148615
rect 106060 -148645 106070 -148615
rect 105270 -148650 106070 -148645
rect 106770 -148600 106780 -148565
rect 107560 -148600 107570 -148565
rect 106770 -148615 107570 -148600
rect 106770 -148645 106780 -148615
rect 107560 -148645 107570 -148615
rect 106770 -148650 107570 -148645
rect 108270 -148600 108280 -148565
rect 109060 -148600 109070 -148565
rect 108270 -148615 109070 -148600
rect 108270 -148645 108280 -148615
rect 109060 -148645 109070 -148615
rect 108270 -148650 109070 -148645
rect 109770 -148600 109780 -148565
rect 110560 -148600 110570 -148565
rect 109770 -148615 110570 -148600
rect 109770 -148645 109780 -148615
rect 110560 -148645 110570 -148615
rect 109770 -148650 110570 -148645
rect 111270 -148600 111280 -148565
rect 112060 -148600 112070 -148565
rect 111270 -148615 112070 -148600
rect 111270 -148645 111280 -148615
rect 112060 -148645 112070 -148615
rect 111270 -148650 112070 -148645
rect 112770 -148600 112780 -148565
rect 113560 -148600 113570 -148565
rect 112770 -148615 113570 -148600
rect 112770 -148645 112780 -148615
rect 113560 -148645 113570 -148615
rect 112770 -148650 113570 -148645
rect 114270 -148600 114280 -148565
rect 115060 -148600 115070 -148565
rect 114270 -148615 115070 -148600
rect 114270 -148645 114280 -148615
rect 115060 -148645 115070 -148615
rect 114270 -148650 115070 -148645
rect 115770 -148600 115780 -148565
rect 116560 -148600 116570 -148565
rect 115770 -148615 116570 -148600
rect 115770 -148645 115780 -148615
rect 116560 -148645 116570 -148615
rect 115770 -148650 116570 -148645
rect 117270 -148600 117280 -148565
rect 118060 -148600 118070 -148565
rect 117270 -148615 118070 -148600
rect 117270 -148645 117280 -148615
rect 118060 -148645 118070 -148615
rect 117270 -148650 118070 -148645
rect 118770 -148600 118780 -148565
rect 119560 -148600 119570 -148565
rect 118770 -148615 119570 -148600
rect 118770 -148645 118780 -148615
rect 119560 -148645 119570 -148615
rect 118770 -148650 119570 -148645
rect 120270 -148600 120280 -148565
rect 121060 -148600 121070 -148565
rect 120270 -148615 121070 -148600
rect 120270 -148645 120280 -148615
rect 121060 -148645 121070 -148615
rect 120270 -148650 121070 -148645
rect 121770 -148600 121780 -148565
rect 122560 -148600 122570 -148565
rect 121770 -148615 122570 -148600
rect 121770 -148645 121780 -148615
rect 122560 -148645 122570 -148615
rect 121770 -148650 122570 -148645
rect 123270 -148600 123280 -148565
rect 124060 -148600 124070 -148565
rect 123270 -148615 124070 -148600
rect 123270 -148645 123280 -148615
rect 124060 -148645 124070 -148615
rect 123270 -148650 124070 -148645
rect 124770 -148600 124780 -148565
rect 125560 -148600 125570 -148565
rect 124770 -148615 125570 -148600
rect 124770 -148645 124780 -148615
rect 125560 -148645 125570 -148615
rect 124770 -148650 125570 -148645
rect 126270 -148600 126280 -148565
rect 127060 -148600 127070 -148565
rect 126270 -148615 127070 -148600
rect 126270 -148645 126280 -148615
rect 127060 -148645 127070 -148615
rect 126270 -148650 127070 -148645
rect 127770 -148600 127780 -148565
rect 128560 -148600 128570 -148565
rect 127770 -148615 128570 -148600
rect 127770 -148645 127780 -148615
rect 128560 -148645 128570 -148615
rect 127770 -148650 128570 -148645
rect 129270 -148600 129280 -148565
rect 130060 -148600 130070 -148565
rect 129270 -148615 130070 -148600
rect 129270 -148645 129280 -148615
rect 130060 -148645 130070 -148615
rect 129270 -148650 130070 -148645
rect 130770 -148600 130780 -148565
rect 131560 -148600 131570 -148565
rect 130770 -148615 131570 -148600
rect 130770 -148645 130780 -148615
rect 131560 -148645 131570 -148615
rect 130770 -148650 131570 -148645
rect 132270 -148600 132280 -148565
rect 133060 -148600 133070 -148565
rect 132270 -148615 133070 -148600
rect 132270 -148645 132280 -148615
rect 133060 -148645 133070 -148615
rect 132270 -148650 133070 -148645
rect 133770 -148600 133780 -148565
rect 134560 -148600 134570 -148565
rect 133770 -148615 134570 -148600
rect 133770 -148645 133780 -148615
rect 134560 -148645 134570 -148615
rect 133770 -148650 134570 -148645
rect 135270 -148600 135280 -148565
rect 136060 -148600 136070 -148565
rect 135270 -148615 136070 -148600
rect 135270 -148645 135280 -148615
rect 136060 -148645 136070 -148615
rect 135270 -148650 136070 -148645
rect 136770 -148600 136780 -148565
rect 137560 -148600 137570 -148565
rect 136770 -148615 137570 -148600
rect 136770 -148645 136780 -148615
rect 137560 -148645 137570 -148615
rect 136770 -148650 137570 -148645
rect 138270 -148600 138280 -148565
rect 139060 -148600 139070 -148565
rect 138270 -148615 139070 -148600
rect 138270 -148645 138280 -148615
rect 139060 -148645 139070 -148615
rect 138270 -148650 139070 -148645
rect 139770 -148600 139780 -148565
rect 140560 -148600 140570 -148565
rect 139770 -148615 140570 -148600
rect 139770 -148645 139780 -148615
rect 140560 -148645 140570 -148615
rect 139770 -148650 140570 -148645
rect 141270 -148600 141280 -148565
rect 142060 -148600 142070 -148565
rect 141270 -148615 142070 -148600
rect 141270 -148645 141280 -148615
rect 142060 -148645 142070 -148615
rect 141270 -148650 142070 -148645
rect 142770 -148600 142780 -148565
rect 143560 -148600 143570 -148565
rect 142770 -148615 143570 -148600
rect 142770 -148645 142780 -148615
rect 143560 -148645 143570 -148615
rect 142770 -148650 143570 -148645
rect 144270 -148600 144280 -148565
rect 145060 -148600 145070 -148565
rect 144270 -148615 145070 -148600
rect 144270 -148645 144280 -148615
rect 145060 -148645 145070 -148615
rect 144270 -148650 145070 -148645
rect 145770 -148600 145780 -148565
rect 146560 -148600 146570 -148565
rect 145770 -148615 146570 -148600
rect 145770 -148645 145780 -148615
rect 146560 -148645 146570 -148615
rect 145770 -148650 146570 -148645
rect 147270 -148600 147280 -148565
rect 148060 -148600 148070 -148565
rect 147270 -148615 148070 -148600
rect 147270 -148645 147280 -148615
rect 148060 -148645 148070 -148615
rect 147270 -148650 148070 -148645
rect 148770 -148600 148780 -148565
rect 149560 -148600 149570 -148565
rect 148770 -148615 149570 -148600
rect 148770 -148645 148780 -148615
rect 149560 -148645 149570 -148615
rect 148770 -148650 149570 -148645
rect 110 -148750 220 -148745
rect 110 -148850 120 -148750
rect 210 -148850 220 -148750
rect 110 -148855 220 -148850
rect 1610 -148750 1720 -148745
rect 1610 -148850 1620 -148750
rect 1710 -148850 1720 -148750
rect 1610 -148855 1720 -148850
rect 3110 -148750 3220 -148745
rect 3110 -148850 3120 -148750
rect 3210 -148850 3220 -148750
rect 3110 -148855 3220 -148850
rect 4610 -148750 4720 -148745
rect 4610 -148850 4620 -148750
rect 4710 -148850 4720 -148750
rect 4610 -148855 4720 -148850
rect 6110 -148750 6220 -148745
rect 6110 -148850 6120 -148750
rect 6210 -148850 6220 -148750
rect 6110 -148855 6220 -148850
rect 7610 -148750 7720 -148745
rect 7610 -148850 7620 -148750
rect 7710 -148850 7720 -148750
rect 7610 -148855 7720 -148850
rect 9110 -148750 9220 -148745
rect 9110 -148850 9120 -148750
rect 9210 -148850 9220 -148750
rect 9110 -148855 9220 -148850
rect 10610 -148750 10720 -148745
rect 10610 -148850 10620 -148750
rect 10710 -148850 10720 -148750
rect 10610 -148855 10720 -148850
rect 12110 -148750 12220 -148745
rect 12110 -148850 12120 -148750
rect 12210 -148850 12220 -148750
rect 12110 -148855 12220 -148850
rect 13610 -148750 13720 -148745
rect 13610 -148850 13620 -148750
rect 13710 -148850 13720 -148750
rect 13610 -148855 13720 -148850
rect 15110 -148750 15220 -148745
rect 15110 -148850 15120 -148750
rect 15210 -148850 15220 -148750
rect 15110 -148855 15220 -148850
rect 16610 -148750 16720 -148745
rect 16610 -148850 16620 -148750
rect 16710 -148850 16720 -148750
rect 16610 -148855 16720 -148850
rect 18110 -148750 18220 -148745
rect 18110 -148850 18120 -148750
rect 18210 -148850 18220 -148750
rect 18110 -148855 18220 -148850
rect 19610 -148750 19720 -148745
rect 19610 -148850 19620 -148750
rect 19710 -148850 19720 -148750
rect 19610 -148855 19720 -148850
rect 21110 -148750 21220 -148745
rect 21110 -148850 21120 -148750
rect 21210 -148850 21220 -148750
rect 21110 -148855 21220 -148850
rect 22610 -148750 22720 -148745
rect 22610 -148850 22620 -148750
rect 22710 -148850 22720 -148750
rect 22610 -148855 22720 -148850
rect 24110 -148750 24220 -148745
rect 24110 -148850 24120 -148750
rect 24210 -148850 24220 -148750
rect 24110 -148855 24220 -148850
rect 25610 -148750 25720 -148745
rect 25610 -148850 25620 -148750
rect 25710 -148850 25720 -148750
rect 25610 -148855 25720 -148850
rect 27110 -148750 27220 -148745
rect 27110 -148850 27120 -148750
rect 27210 -148850 27220 -148750
rect 27110 -148855 27220 -148850
rect 28610 -148750 28720 -148745
rect 28610 -148850 28620 -148750
rect 28710 -148850 28720 -148750
rect 28610 -148855 28720 -148850
rect 30110 -148750 30220 -148745
rect 30110 -148850 30120 -148750
rect 30210 -148850 30220 -148750
rect 30110 -148855 30220 -148850
rect 31610 -148750 31720 -148745
rect 31610 -148850 31620 -148750
rect 31710 -148850 31720 -148750
rect 31610 -148855 31720 -148850
rect 33110 -148750 33220 -148745
rect 33110 -148850 33120 -148750
rect 33210 -148850 33220 -148750
rect 33110 -148855 33220 -148850
rect 34610 -148750 34720 -148745
rect 34610 -148850 34620 -148750
rect 34710 -148850 34720 -148750
rect 34610 -148855 34720 -148850
rect 36110 -148750 36220 -148745
rect 36110 -148850 36120 -148750
rect 36210 -148850 36220 -148750
rect 36110 -148855 36220 -148850
rect 37610 -148750 37720 -148745
rect 37610 -148850 37620 -148750
rect 37710 -148850 37720 -148750
rect 37610 -148855 37720 -148850
rect 39110 -148750 39220 -148745
rect 39110 -148850 39120 -148750
rect 39210 -148850 39220 -148750
rect 39110 -148855 39220 -148850
rect 40610 -148750 40720 -148745
rect 40610 -148850 40620 -148750
rect 40710 -148850 40720 -148750
rect 40610 -148855 40720 -148850
rect 42110 -148750 42220 -148745
rect 42110 -148850 42120 -148750
rect 42210 -148850 42220 -148750
rect 42110 -148855 42220 -148850
rect 43610 -148750 43720 -148745
rect 43610 -148850 43620 -148750
rect 43710 -148850 43720 -148750
rect 43610 -148855 43720 -148850
rect 45110 -148750 45220 -148745
rect 45110 -148850 45120 -148750
rect 45210 -148850 45220 -148750
rect 45110 -148855 45220 -148850
rect 46610 -148750 46720 -148745
rect 46610 -148850 46620 -148750
rect 46710 -148850 46720 -148750
rect 46610 -148855 46720 -148850
rect 48110 -148750 48220 -148745
rect 48110 -148850 48120 -148750
rect 48210 -148850 48220 -148750
rect 48110 -148855 48220 -148850
rect 49610 -148750 49720 -148745
rect 49610 -148850 49620 -148750
rect 49710 -148850 49720 -148750
rect 49610 -148855 49720 -148850
rect 51110 -148750 51220 -148745
rect 51110 -148850 51120 -148750
rect 51210 -148850 51220 -148750
rect 51110 -148855 51220 -148850
rect 52610 -148750 52720 -148745
rect 52610 -148850 52620 -148750
rect 52710 -148850 52720 -148750
rect 52610 -148855 52720 -148850
rect 54110 -148750 54220 -148745
rect 54110 -148850 54120 -148750
rect 54210 -148850 54220 -148750
rect 54110 -148855 54220 -148850
rect 55610 -148750 55720 -148745
rect 55610 -148850 55620 -148750
rect 55710 -148850 55720 -148750
rect 55610 -148855 55720 -148850
rect 57110 -148750 57220 -148745
rect 57110 -148850 57120 -148750
rect 57210 -148850 57220 -148750
rect 57110 -148855 57220 -148850
rect 58610 -148750 58720 -148745
rect 58610 -148850 58620 -148750
rect 58710 -148850 58720 -148750
rect 58610 -148855 58720 -148850
rect 60110 -148750 60220 -148745
rect 60110 -148850 60120 -148750
rect 60210 -148850 60220 -148750
rect 60110 -148855 60220 -148850
rect 61610 -148750 61720 -148745
rect 61610 -148850 61620 -148750
rect 61710 -148850 61720 -148750
rect 61610 -148855 61720 -148850
rect 63110 -148750 63220 -148745
rect 63110 -148850 63120 -148750
rect 63210 -148850 63220 -148750
rect 63110 -148855 63220 -148850
rect 64610 -148750 64720 -148745
rect 64610 -148850 64620 -148750
rect 64710 -148850 64720 -148750
rect 64610 -148855 64720 -148850
rect 66110 -148750 66220 -148745
rect 66110 -148850 66120 -148750
rect 66210 -148850 66220 -148750
rect 66110 -148855 66220 -148850
rect 67610 -148750 67720 -148745
rect 67610 -148850 67620 -148750
rect 67710 -148850 67720 -148750
rect 67610 -148855 67720 -148850
rect 69110 -148750 69220 -148745
rect 69110 -148850 69120 -148750
rect 69210 -148850 69220 -148750
rect 69110 -148855 69220 -148850
rect 70610 -148750 70720 -148745
rect 70610 -148850 70620 -148750
rect 70710 -148850 70720 -148750
rect 70610 -148855 70720 -148850
rect 72110 -148750 72220 -148745
rect 72110 -148850 72120 -148750
rect 72210 -148850 72220 -148750
rect 72110 -148855 72220 -148850
rect 73610 -148750 73720 -148745
rect 73610 -148850 73620 -148750
rect 73710 -148850 73720 -148750
rect 73610 -148855 73720 -148850
rect 75110 -148750 75220 -148745
rect 75110 -148850 75120 -148750
rect 75210 -148850 75220 -148750
rect 75110 -148855 75220 -148850
rect 76610 -148750 76720 -148745
rect 76610 -148850 76620 -148750
rect 76710 -148850 76720 -148750
rect 76610 -148855 76720 -148850
rect 78110 -148750 78220 -148745
rect 78110 -148850 78120 -148750
rect 78210 -148850 78220 -148750
rect 78110 -148855 78220 -148850
rect 79610 -148750 79720 -148745
rect 79610 -148850 79620 -148750
rect 79710 -148850 79720 -148750
rect 79610 -148855 79720 -148850
rect 81110 -148750 81220 -148745
rect 81110 -148850 81120 -148750
rect 81210 -148850 81220 -148750
rect 81110 -148855 81220 -148850
rect 82610 -148750 82720 -148745
rect 82610 -148850 82620 -148750
rect 82710 -148850 82720 -148750
rect 82610 -148855 82720 -148850
rect 84110 -148750 84220 -148745
rect 84110 -148850 84120 -148750
rect 84210 -148850 84220 -148750
rect 84110 -148855 84220 -148850
rect 85610 -148750 85720 -148745
rect 85610 -148850 85620 -148750
rect 85710 -148850 85720 -148750
rect 85610 -148855 85720 -148850
rect 87110 -148750 87220 -148745
rect 87110 -148850 87120 -148750
rect 87210 -148850 87220 -148750
rect 87110 -148855 87220 -148850
rect 88610 -148750 88720 -148745
rect 88610 -148850 88620 -148750
rect 88710 -148850 88720 -148750
rect 88610 -148855 88720 -148850
rect 90110 -148750 90220 -148745
rect 90110 -148850 90120 -148750
rect 90210 -148850 90220 -148750
rect 90110 -148855 90220 -148850
rect 91610 -148750 91720 -148745
rect 91610 -148850 91620 -148750
rect 91710 -148850 91720 -148750
rect 91610 -148855 91720 -148850
rect 93110 -148750 93220 -148745
rect 93110 -148850 93120 -148750
rect 93210 -148850 93220 -148750
rect 93110 -148855 93220 -148850
rect 94610 -148750 94720 -148745
rect 94610 -148850 94620 -148750
rect 94710 -148850 94720 -148750
rect 94610 -148855 94720 -148850
rect 96110 -148750 96220 -148745
rect 96110 -148850 96120 -148750
rect 96210 -148850 96220 -148750
rect 96110 -148855 96220 -148850
rect 97610 -148750 97720 -148745
rect 97610 -148850 97620 -148750
rect 97710 -148850 97720 -148750
rect 97610 -148855 97720 -148850
rect 99110 -148750 99220 -148745
rect 99110 -148850 99120 -148750
rect 99210 -148850 99220 -148750
rect 99110 -148855 99220 -148850
rect 100610 -148750 100720 -148745
rect 100610 -148850 100620 -148750
rect 100710 -148850 100720 -148750
rect 100610 -148855 100720 -148850
rect 102110 -148750 102220 -148745
rect 102110 -148850 102120 -148750
rect 102210 -148850 102220 -148750
rect 102110 -148855 102220 -148850
rect 103610 -148750 103720 -148745
rect 103610 -148850 103620 -148750
rect 103710 -148850 103720 -148750
rect 103610 -148855 103720 -148850
rect 105110 -148750 105220 -148745
rect 105110 -148850 105120 -148750
rect 105210 -148850 105220 -148750
rect 105110 -148855 105220 -148850
rect 106610 -148750 106720 -148745
rect 106610 -148850 106620 -148750
rect 106710 -148850 106720 -148750
rect 106610 -148855 106720 -148850
rect 108110 -148750 108220 -148745
rect 108110 -148850 108120 -148750
rect 108210 -148850 108220 -148750
rect 108110 -148855 108220 -148850
rect 109610 -148750 109720 -148745
rect 109610 -148850 109620 -148750
rect 109710 -148850 109720 -148750
rect 109610 -148855 109720 -148850
rect 111110 -148750 111220 -148745
rect 111110 -148850 111120 -148750
rect 111210 -148850 111220 -148750
rect 111110 -148855 111220 -148850
rect 112610 -148750 112720 -148745
rect 112610 -148850 112620 -148750
rect 112710 -148850 112720 -148750
rect 112610 -148855 112720 -148850
rect 114110 -148750 114220 -148745
rect 114110 -148850 114120 -148750
rect 114210 -148850 114220 -148750
rect 114110 -148855 114220 -148850
rect 115610 -148750 115720 -148745
rect 115610 -148850 115620 -148750
rect 115710 -148850 115720 -148750
rect 115610 -148855 115720 -148850
rect 117110 -148750 117220 -148745
rect 117110 -148850 117120 -148750
rect 117210 -148850 117220 -148750
rect 117110 -148855 117220 -148850
rect 118610 -148750 118720 -148745
rect 118610 -148850 118620 -148750
rect 118710 -148850 118720 -148750
rect 118610 -148855 118720 -148850
rect 120110 -148750 120220 -148745
rect 120110 -148850 120120 -148750
rect 120210 -148850 120220 -148750
rect 120110 -148855 120220 -148850
rect 121610 -148750 121720 -148745
rect 121610 -148850 121620 -148750
rect 121710 -148850 121720 -148750
rect 121610 -148855 121720 -148850
rect 123110 -148750 123220 -148745
rect 123110 -148850 123120 -148750
rect 123210 -148850 123220 -148750
rect 123110 -148855 123220 -148850
rect 124610 -148750 124720 -148745
rect 124610 -148850 124620 -148750
rect 124710 -148850 124720 -148750
rect 124610 -148855 124720 -148850
rect 126110 -148750 126220 -148745
rect 126110 -148850 126120 -148750
rect 126210 -148850 126220 -148750
rect 126110 -148855 126220 -148850
rect 127610 -148750 127720 -148745
rect 127610 -148850 127620 -148750
rect 127710 -148850 127720 -148750
rect 127610 -148855 127720 -148850
rect 129110 -148750 129220 -148745
rect 129110 -148850 129120 -148750
rect 129210 -148850 129220 -148750
rect 129110 -148855 129220 -148850
rect 130610 -148750 130720 -148745
rect 130610 -148850 130620 -148750
rect 130710 -148850 130720 -148750
rect 130610 -148855 130720 -148850
rect 132110 -148750 132220 -148745
rect 132110 -148850 132120 -148750
rect 132210 -148850 132220 -148750
rect 132110 -148855 132220 -148850
rect 133610 -148750 133720 -148745
rect 133610 -148850 133620 -148750
rect 133710 -148850 133720 -148750
rect 133610 -148855 133720 -148850
rect 135110 -148750 135220 -148745
rect 135110 -148850 135120 -148750
rect 135210 -148850 135220 -148750
rect 135110 -148855 135220 -148850
rect 136610 -148750 136720 -148745
rect 136610 -148850 136620 -148750
rect 136710 -148850 136720 -148750
rect 136610 -148855 136720 -148850
rect 138110 -148750 138220 -148745
rect 138110 -148850 138120 -148750
rect 138210 -148850 138220 -148750
rect 138110 -148855 138220 -148850
rect 139610 -148750 139720 -148745
rect 139610 -148850 139620 -148750
rect 139710 -148850 139720 -148750
rect 139610 -148855 139720 -148850
rect 141110 -148750 141220 -148745
rect 141110 -148850 141120 -148750
rect 141210 -148850 141220 -148750
rect 141110 -148855 141220 -148850
rect 142610 -148750 142720 -148745
rect 142610 -148850 142620 -148750
rect 142710 -148850 142720 -148750
rect 142610 -148855 142720 -148850
rect 144110 -148750 144220 -148745
rect 144110 -148850 144120 -148750
rect 144210 -148850 144220 -148750
rect 144110 -148855 144220 -148850
rect 145610 -148750 145720 -148745
rect 145610 -148850 145620 -148750
rect 145710 -148850 145720 -148750
rect 145610 -148855 145720 -148850
rect 147110 -148750 147220 -148745
rect 147110 -148850 147120 -148750
rect 147210 -148850 147220 -148750
rect 147110 -148855 147220 -148850
rect 148610 -148750 148720 -148745
rect 148610 -148850 148620 -148750
rect 148710 -148850 148720 -148750
rect 148610 -148855 148720 -148850
rect 270 -148960 150370 -148950
rect 270 -149040 280 -148960
rect 270 -149050 150370 -149040
<< via1 >>
rect -960 1680 -450 1725
rect 25 1680 70 1725
rect 1525 1680 1570 1725
rect 3025 1680 3070 1725
rect 4525 1680 4570 1725
rect 6025 1680 6070 1725
rect 7525 1680 7570 1725
rect 9025 1680 9070 1725
rect 10525 1680 10570 1725
rect 12025 1680 12070 1725
rect 13525 1680 13570 1725
rect 15025 1680 15070 1725
rect 16525 1680 16570 1725
rect 18025 1680 18070 1725
rect 19525 1680 19570 1725
rect 21025 1680 21070 1725
rect 22525 1680 22570 1725
rect 24025 1680 24070 1725
rect 25525 1680 25570 1725
rect 27025 1680 27070 1725
rect 28525 1680 28570 1725
rect 30025 1680 30070 1725
rect 31525 1680 31570 1725
rect 33025 1680 33070 1725
rect 34525 1680 34570 1725
rect 36025 1680 36070 1725
rect 37525 1680 37570 1725
rect 39025 1680 39070 1725
rect 40525 1680 40570 1725
rect 42025 1680 42070 1725
rect 43525 1680 43570 1725
rect 45025 1680 45070 1725
rect 46525 1680 46570 1725
rect 48025 1680 48070 1725
rect 49525 1680 49570 1725
rect 51025 1680 51070 1725
rect 52525 1680 52570 1725
rect 54025 1680 54070 1725
rect 55525 1680 55570 1725
rect 57025 1680 57070 1725
rect 58525 1680 58570 1725
rect 60025 1680 60070 1725
rect 61525 1680 61570 1725
rect 63025 1680 63070 1725
rect 64525 1680 64570 1725
rect 66025 1680 66070 1725
rect 67525 1680 67570 1725
rect 69025 1680 69070 1725
rect 70525 1680 70570 1725
rect 72025 1680 72070 1725
rect 73525 1680 73570 1725
rect 75025 1680 75070 1725
rect 76525 1680 76570 1725
rect 78025 1680 78070 1725
rect 79525 1680 79570 1725
rect 81025 1680 81070 1725
rect 82525 1680 82570 1725
rect 84025 1680 84070 1725
rect 85525 1680 85570 1725
rect 87025 1680 87070 1725
rect 88525 1680 88570 1725
rect 90025 1680 90070 1725
rect 91525 1680 91570 1725
rect 93025 1680 93070 1725
rect 94525 1680 94570 1725
rect 96025 1680 96070 1725
rect 97525 1680 97570 1725
rect 99025 1680 99070 1725
rect 100525 1680 100570 1725
rect 102025 1680 102070 1725
rect 103525 1680 103570 1725
rect 105025 1680 105070 1725
rect 106525 1680 106570 1725
rect 108025 1680 108070 1725
rect 109525 1680 109570 1725
rect 111025 1680 111070 1725
rect 112525 1680 112570 1725
rect 114025 1680 114070 1725
rect 115525 1680 115570 1725
rect 117025 1680 117070 1725
rect 118525 1680 118570 1725
rect 120025 1680 120070 1725
rect 121525 1680 121570 1725
rect 123025 1680 123070 1725
rect 124525 1680 124570 1725
rect 126025 1680 126070 1725
rect 127525 1680 127570 1725
rect 129025 1680 129070 1725
rect 130525 1680 130570 1725
rect 132025 1680 132070 1725
rect 133525 1680 133570 1725
rect 135025 1680 135070 1725
rect 136525 1680 136570 1725
rect 138025 1680 138070 1725
rect 139525 1680 139570 1725
rect 141025 1680 141070 1725
rect 142525 1680 142570 1725
rect 144025 1680 144070 1725
rect 145525 1680 145570 1725
rect 147025 1680 147070 1725
rect 148525 1680 148570 1725
rect -790 745 -590 780
rect -270 745 -130 780
rect -790 -755 -590 -720
rect -270 -755 -130 -720
rect -790 -2255 -590 -2220
rect -270 -2255 -130 -2220
rect -790 -3755 -590 -3720
rect -270 -3755 -130 -3720
rect -790 -5255 -590 -5220
rect -270 -5255 -130 -5220
rect -790 -6755 -590 -6720
rect -270 -6755 -130 -6720
rect -790 -8255 -590 -8220
rect -270 -8255 -130 -8220
rect -790 -9755 -590 -9720
rect -270 -9755 -130 -9720
rect -790 -11255 -590 -11220
rect -270 -11255 -130 -11220
rect -790 -12755 -590 -12720
rect -270 -12755 -130 -12720
rect -790 -14255 -590 -14220
rect -270 -14255 -130 -14220
rect -790 -15755 -590 -15720
rect -270 -15755 -130 -15720
rect -790 -17255 -590 -17220
rect -270 -17255 -130 -17220
rect -790 -18755 -590 -18720
rect -270 -18755 -130 -18720
rect -790 -20255 -590 -20220
rect -270 -20255 -130 -20220
rect -790 -21755 -590 -21720
rect -270 -21755 -130 -21720
rect -790 -23255 -590 -23220
rect -270 -23255 -130 -23220
rect -790 -24755 -590 -24720
rect -270 -24755 -130 -24720
rect -790 -26255 -590 -26220
rect -270 -26255 -130 -26220
rect -790 -27755 -590 -27720
rect -270 -27755 -130 -27720
rect -790 -29255 -590 -29220
rect -270 -29255 -130 -29220
rect -790 -30755 -590 -30720
rect -270 -30755 -130 -30720
rect -790 -32255 -590 -32220
rect -270 -32255 -130 -32220
rect -790 -33755 -590 -33720
rect -270 -33755 -130 -33720
rect -790 -35255 -590 -35220
rect -270 -35255 -130 -35220
rect -790 -36755 -590 -36720
rect -270 -36755 -130 -36720
rect -790 -38255 -590 -38220
rect -270 -38255 -130 -38220
rect -790 -39755 -590 -39720
rect -270 -39755 -130 -39720
rect -790 -41255 -590 -41220
rect -270 -41255 -130 -41220
rect -790 -42755 -590 -42720
rect -270 -42755 -130 -42720
rect -790 -44255 -590 -44220
rect -270 -44255 -130 -44220
rect -790 -45755 -590 -45720
rect -270 -45755 -130 -45720
rect -790 -47255 -590 -47220
rect -270 -47255 -130 -47220
rect -790 -48755 -590 -48720
rect -270 -48755 -130 -48720
rect -790 -50255 -590 -50220
rect -270 -50255 -130 -50220
rect -790 -51755 -590 -51720
rect -270 -51755 -130 -51720
rect -790 -53255 -590 -53220
rect -270 -53255 -130 -53220
rect -790 -54755 -590 -54720
rect -270 -54755 -130 -54720
rect -790 -56255 -590 -56220
rect -270 -56255 -130 -56220
rect -790 -57755 -590 -57720
rect -270 -57755 -130 -57720
rect -790 -59255 -590 -59220
rect -270 -59255 -130 -59220
rect -790 -60755 -590 -60720
rect -270 -60755 -130 -60720
rect -790 -62255 -590 -62220
rect -270 -62255 -130 -62220
rect -790 -63755 -590 -63720
rect -270 -63755 -130 -63720
rect -790 -65255 -590 -65220
rect -270 -65255 -130 -65220
rect -790 -66755 -590 -66720
rect -270 -66755 -130 -66720
rect -790 -68255 -590 -68220
rect -270 -68255 -130 -68220
rect -790 -69755 -590 -69720
rect -270 -69755 -130 -69720
rect -790 -71255 -590 -71220
rect -270 -71255 -130 -71220
rect -790 -72755 -590 -72720
rect -270 -72755 -130 -72720
rect -790 -74255 -590 -74220
rect -270 -74255 -130 -74220
rect -790 -75755 -590 -75720
rect -270 -75755 -130 -75720
rect -790 -77255 -590 -77220
rect -270 -77255 -130 -77220
rect -790 -78755 -590 -78720
rect -270 -78755 -130 -78720
rect -790 -80255 -590 -80220
rect -270 -80255 -130 -80220
rect -790 -81755 -590 -81720
rect -270 -81755 -130 -81720
rect -790 -83255 -590 -83220
rect -270 -83255 -130 -83220
rect -790 -84755 -590 -84720
rect -270 -84755 -130 -84720
rect -790 -86255 -590 -86220
rect -270 -86255 -130 -86220
rect -790 -87755 -590 -87720
rect -270 -87755 -130 -87720
rect -790 -89255 -590 -89220
rect -270 -89255 -130 -89220
rect -790 -90755 -590 -90720
rect -270 -90755 -130 -90720
rect -790 -92255 -590 -92220
rect -270 -92255 -130 -92220
rect -790 -93755 -590 -93720
rect -270 -93755 -130 -93720
rect -790 -95255 -590 -95220
rect -270 -95255 -130 -95220
rect -790 -96755 -590 -96720
rect -270 -96755 -130 -96720
rect -790 -98255 -590 -98220
rect -270 -98255 -130 -98220
rect -790 -99755 -590 -99720
rect -270 -99755 -130 -99720
rect -790 -101255 -590 -101220
rect -270 -101255 -130 -101220
rect -790 -102755 -590 -102720
rect -270 -102755 -130 -102720
rect -790 -104255 -590 -104220
rect -270 -104255 -130 -104220
rect -790 -105755 -590 -105720
rect -270 -105755 -130 -105720
rect -790 -107255 -590 -107220
rect -270 -107255 -130 -107220
rect -790 -108755 -590 -108720
rect -270 -108755 -130 -108720
rect -790 -110255 -590 -110220
rect -270 -110255 -130 -110220
rect -790 -111755 -590 -111720
rect -270 -111755 -130 -111720
rect -790 -113255 -590 -113220
rect -270 -113255 -130 -113220
rect -790 -114755 -590 -114720
rect -270 -114755 -130 -114720
rect -790 -116255 -590 -116220
rect -270 -116255 -130 -116220
rect -790 -117755 -590 -117720
rect -270 -117755 -130 -117720
rect -790 -119255 -590 -119220
rect -270 -119255 -130 -119220
rect -790 -120755 -590 -120720
rect -270 -120755 -130 -120720
rect -790 -122255 -590 -122220
rect -270 -122255 -130 -122220
rect -790 -123755 -590 -123720
rect -270 -123755 -130 -123720
rect -790 -125255 -590 -125220
rect -270 -125255 -130 -125220
rect -790 -126755 -590 -126720
rect -270 -126755 -130 -126720
rect -790 -128255 -590 -128220
rect -270 -128255 -130 -128220
rect -790 -129755 -590 -129720
rect -270 -129755 -130 -129720
rect -790 -131255 -590 -131220
rect -270 -131255 -130 -131220
rect -790 -132755 -590 -132720
rect -270 -132755 -130 -132720
rect -790 -134255 -590 -134220
rect -270 -134255 -130 -134220
rect -790 -135755 -590 -135720
rect -270 -135755 -130 -135720
rect -790 -137255 -590 -137220
rect -270 -137255 -130 -137220
rect -790 -138755 -590 -138720
rect -270 -138755 -130 -138720
rect -790 -140255 -590 -140220
rect -270 -140255 -130 -140220
rect -790 -141755 -590 -141720
rect -270 -141755 -130 -141720
rect -790 -143255 -590 -143220
rect -270 -143255 -130 -143220
rect -790 -144755 -590 -144720
rect -270 -144755 -130 -144720
rect -790 -146255 -590 -146220
rect -270 -146255 -130 -146220
rect -790 -147755 -590 -147720
rect -270 -147755 -130 -147720
rect 280 -148600 1060 -148565
rect 1780 -148600 2560 -148565
rect 3280 -148600 4060 -148565
rect 4780 -148600 5560 -148565
rect 6280 -148600 7060 -148565
rect 7780 -148600 8560 -148565
rect 9280 -148600 10060 -148565
rect 10780 -148600 11560 -148565
rect 12280 -148600 13060 -148565
rect 13780 -148600 14560 -148565
rect 15280 -148600 16060 -148565
rect 16780 -148600 17560 -148565
rect 18280 -148600 19060 -148565
rect 19780 -148600 20560 -148565
rect 21280 -148600 22060 -148565
rect 22780 -148600 23560 -148565
rect 24280 -148600 25060 -148565
rect 25780 -148600 26560 -148565
rect 27280 -148600 28060 -148565
rect 28780 -148600 29560 -148565
rect 30280 -148600 31060 -148565
rect 31780 -148600 32560 -148565
rect 33280 -148600 34060 -148565
rect 34780 -148600 35560 -148565
rect 36280 -148600 37060 -148565
rect 37780 -148600 38560 -148565
rect 39280 -148600 40060 -148565
rect 40780 -148600 41560 -148565
rect 42280 -148600 43060 -148565
rect 43780 -148600 44560 -148565
rect 45280 -148600 46060 -148565
rect 46780 -148600 47560 -148565
rect 48280 -148600 49060 -148565
rect 49780 -148600 50560 -148565
rect 51280 -148600 52060 -148565
rect 52780 -148600 53560 -148565
rect 54280 -148600 55060 -148565
rect 55780 -148600 56560 -148565
rect 57280 -148600 58060 -148565
rect 58780 -148600 59560 -148565
rect 60280 -148600 61060 -148565
rect 61780 -148600 62560 -148565
rect 63280 -148600 64060 -148565
rect 64780 -148600 65560 -148565
rect 66280 -148600 67060 -148565
rect 67780 -148600 68560 -148565
rect 69280 -148600 70060 -148565
rect 70780 -148600 71560 -148565
rect 72280 -148600 73060 -148565
rect 73780 -148600 74560 -148565
rect 75280 -148600 76060 -148565
rect 76780 -148600 77560 -148565
rect 78280 -148600 79060 -148565
rect 79780 -148600 80560 -148565
rect 81280 -148600 82060 -148565
rect 82780 -148600 83560 -148565
rect 84280 -148600 85060 -148565
rect 85780 -148600 86560 -148565
rect 87280 -148600 88060 -148565
rect 88780 -148600 89560 -148565
rect 90280 -148600 91060 -148565
rect 91780 -148600 92560 -148565
rect 93280 -148600 94060 -148565
rect 94780 -148600 95560 -148565
rect 96280 -148600 97060 -148565
rect 97780 -148600 98560 -148565
rect 99280 -148600 100060 -148565
rect 100780 -148600 101560 -148565
rect 102280 -148600 103060 -148565
rect 103780 -148600 104560 -148565
rect 105280 -148600 106060 -148565
rect 106780 -148600 107560 -148565
rect 108280 -148600 109060 -148565
rect 109780 -148600 110560 -148565
rect 111280 -148600 112060 -148565
rect 112780 -148600 113560 -148565
rect 114280 -148600 115060 -148565
rect 115780 -148600 116560 -148565
rect 117280 -148600 118060 -148565
rect 118780 -148600 119560 -148565
rect 120280 -148600 121060 -148565
rect 121780 -148600 122560 -148565
rect 123280 -148600 124060 -148565
rect 124780 -148600 125560 -148565
rect 126280 -148600 127060 -148565
rect 127780 -148600 128560 -148565
rect 129280 -148600 130060 -148565
rect 130780 -148600 131560 -148565
rect 132280 -148600 133060 -148565
rect 133780 -148600 134560 -148565
rect 135280 -148600 136060 -148565
rect 136780 -148600 137560 -148565
rect 138280 -148600 139060 -148565
rect 139780 -148600 140560 -148565
rect 141280 -148600 142060 -148565
rect 142780 -148600 143560 -148565
rect 144280 -148600 145060 -148565
rect 145780 -148600 146560 -148565
rect 147280 -148600 148060 -148565
rect 148780 -148600 149560 -148565
rect 120 -148850 210 -148750
rect 1620 -148850 1710 -148750
rect 3120 -148850 3210 -148750
rect 4620 -148850 4710 -148750
rect 6120 -148850 6210 -148750
rect 7620 -148850 7710 -148750
rect 9120 -148850 9210 -148750
rect 10620 -148850 10710 -148750
rect 12120 -148850 12210 -148750
rect 13620 -148850 13710 -148750
rect 15120 -148850 15210 -148750
rect 16620 -148850 16710 -148750
rect 18120 -148850 18210 -148750
rect 19620 -148850 19710 -148750
rect 21120 -148850 21210 -148750
rect 22620 -148850 22710 -148750
rect 24120 -148850 24210 -148750
rect 25620 -148850 25710 -148750
rect 27120 -148850 27210 -148750
rect 28620 -148850 28710 -148750
rect 30120 -148850 30210 -148750
rect 31620 -148850 31710 -148750
rect 33120 -148850 33210 -148750
rect 34620 -148850 34710 -148750
rect 36120 -148850 36210 -148750
rect 37620 -148850 37710 -148750
rect 39120 -148850 39210 -148750
rect 40620 -148850 40710 -148750
rect 42120 -148850 42210 -148750
rect 43620 -148850 43710 -148750
rect 45120 -148850 45210 -148750
rect 46620 -148850 46710 -148750
rect 48120 -148850 48210 -148750
rect 49620 -148850 49710 -148750
rect 51120 -148850 51210 -148750
rect 52620 -148850 52710 -148750
rect 54120 -148850 54210 -148750
rect 55620 -148850 55710 -148750
rect 57120 -148850 57210 -148750
rect 58620 -148850 58710 -148750
rect 60120 -148850 60210 -148750
rect 61620 -148850 61710 -148750
rect 63120 -148850 63210 -148750
rect 64620 -148850 64710 -148750
rect 66120 -148850 66210 -148750
rect 67620 -148850 67710 -148750
rect 69120 -148850 69210 -148750
rect 70620 -148850 70710 -148750
rect 72120 -148850 72210 -148750
rect 73620 -148850 73710 -148750
rect 75120 -148850 75210 -148750
rect 76620 -148850 76710 -148750
rect 78120 -148850 78210 -148750
rect 79620 -148850 79710 -148750
rect 81120 -148850 81210 -148750
rect 82620 -148850 82710 -148750
rect 84120 -148850 84210 -148750
rect 85620 -148850 85710 -148750
rect 87120 -148850 87210 -148750
rect 88620 -148850 88710 -148750
rect 90120 -148850 90210 -148750
rect 91620 -148850 91710 -148750
rect 93120 -148850 93210 -148750
rect 94620 -148850 94710 -148750
rect 96120 -148850 96210 -148750
rect 97620 -148850 97710 -148750
rect 99120 -148850 99210 -148750
rect 100620 -148850 100710 -148750
rect 102120 -148850 102210 -148750
rect 103620 -148850 103710 -148750
rect 105120 -148850 105210 -148750
rect 106620 -148850 106710 -148750
rect 108120 -148850 108210 -148750
rect 109620 -148850 109710 -148750
rect 111120 -148850 111210 -148750
rect 112620 -148850 112710 -148750
rect 114120 -148850 114210 -148750
rect 115620 -148850 115710 -148750
rect 117120 -148850 117210 -148750
rect 118620 -148850 118710 -148750
rect 120120 -148850 120210 -148750
rect 121620 -148850 121710 -148750
rect 123120 -148850 123210 -148750
rect 124620 -148850 124710 -148750
rect 126120 -148850 126210 -148750
rect 127620 -148850 127710 -148750
rect 129120 -148850 129210 -148750
rect 130620 -148850 130710 -148750
rect 132120 -148850 132210 -148750
rect 133620 -148850 133710 -148750
rect 135120 -148850 135210 -148750
rect 136620 -148850 136710 -148750
rect 138120 -148850 138210 -148750
rect 139620 -148850 139710 -148750
rect 141120 -148850 141210 -148750
rect 142620 -148850 142710 -148750
rect 144120 -148850 144210 -148750
rect 145620 -148850 145710 -148750
rect 147120 -148850 147210 -148750
rect 148620 -148850 148710 -148750
rect 280 -148990 1060 -148960
rect 1060 -148990 1780 -148960
rect 1780 -148990 2560 -148960
rect 2560 -148990 3280 -148960
rect 3280 -148990 4060 -148960
rect 4060 -148990 4780 -148960
rect 4780 -148990 5560 -148960
rect 5560 -148990 6280 -148960
rect 6280 -148990 7060 -148960
rect 7060 -148990 7780 -148960
rect 7780 -148990 8560 -148960
rect 8560 -148990 9280 -148960
rect 9280 -148990 10060 -148960
rect 10060 -148990 10780 -148960
rect 10780 -148990 11560 -148960
rect 11560 -148990 12280 -148960
rect 12280 -148990 13060 -148960
rect 13060 -148990 13780 -148960
rect 13780 -148990 14560 -148960
rect 14560 -148990 15280 -148960
rect 15280 -148990 16060 -148960
rect 16060 -148990 16780 -148960
rect 16780 -148990 17560 -148960
rect 17560 -148990 18280 -148960
rect 18280 -148990 19060 -148960
rect 19060 -148990 19780 -148960
rect 19780 -148990 20560 -148960
rect 20560 -148990 21280 -148960
rect 21280 -148990 22060 -148960
rect 22060 -148990 22780 -148960
rect 22780 -148990 23560 -148960
rect 23560 -148990 24280 -148960
rect 24280 -148990 25060 -148960
rect 25060 -148990 25780 -148960
rect 25780 -148990 26560 -148960
rect 26560 -148990 27280 -148960
rect 27280 -148990 28060 -148960
rect 28060 -148990 28780 -148960
rect 28780 -148990 29560 -148960
rect 29560 -148990 30280 -148960
rect 30280 -148990 31060 -148960
rect 31060 -148990 31780 -148960
rect 31780 -148990 32560 -148960
rect 32560 -148990 33280 -148960
rect 33280 -148990 34060 -148960
rect 34060 -148990 34780 -148960
rect 34780 -148990 35560 -148960
rect 35560 -148990 36280 -148960
rect 36280 -148990 37060 -148960
rect 37060 -148990 37780 -148960
rect 37780 -148990 38560 -148960
rect 38560 -148990 39280 -148960
rect 39280 -148990 40060 -148960
rect 40060 -148990 40780 -148960
rect 40780 -148990 41560 -148960
rect 41560 -148990 42280 -148960
rect 42280 -148990 43060 -148960
rect 43060 -148990 43780 -148960
rect 43780 -148990 44560 -148960
rect 44560 -148990 45280 -148960
rect 45280 -148990 46060 -148960
rect 46060 -148990 46780 -148960
rect 46780 -148990 47560 -148960
rect 47560 -148990 48280 -148960
rect 48280 -148990 49060 -148960
rect 49060 -148990 49780 -148960
rect 49780 -148990 50560 -148960
rect 50560 -148990 51280 -148960
rect 51280 -148990 52060 -148960
rect 52060 -148990 52780 -148960
rect 52780 -148990 53560 -148960
rect 53560 -148990 54280 -148960
rect 54280 -148990 55060 -148960
rect 55060 -148990 55780 -148960
rect 55780 -148990 56560 -148960
rect 56560 -148990 57280 -148960
rect 57280 -148990 58060 -148960
rect 58060 -148990 58780 -148960
rect 58780 -148990 59560 -148960
rect 59560 -148990 60280 -148960
rect 60280 -148990 61060 -148960
rect 61060 -148990 61780 -148960
rect 61780 -148990 62560 -148960
rect 62560 -148990 63280 -148960
rect 63280 -148990 64060 -148960
rect 64060 -148990 64780 -148960
rect 64780 -148990 65560 -148960
rect 65560 -148990 66280 -148960
rect 66280 -148990 67060 -148960
rect 67060 -148990 67780 -148960
rect 67780 -148990 68560 -148960
rect 68560 -148990 69280 -148960
rect 69280 -148990 70060 -148960
rect 70060 -148990 70780 -148960
rect 70780 -148990 71560 -148960
rect 71560 -148990 72280 -148960
rect 72280 -148990 73060 -148960
rect 73060 -148990 73780 -148960
rect 73780 -148990 74560 -148960
rect 74560 -148990 75280 -148960
rect 75280 -148990 76060 -148960
rect 76060 -148990 76780 -148960
rect 76780 -148990 77560 -148960
rect 77560 -148990 78280 -148960
rect 78280 -148990 79060 -148960
rect 79060 -148990 79780 -148960
rect 79780 -148990 80560 -148960
rect 80560 -148990 81280 -148960
rect 81280 -148990 82060 -148960
rect 82060 -148990 82780 -148960
rect 82780 -148990 83560 -148960
rect 83560 -148990 84280 -148960
rect 84280 -148990 85060 -148960
rect 85060 -148990 85780 -148960
rect 85780 -148990 86560 -148960
rect 86560 -148990 87280 -148960
rect 87280 -148990 88060 -148960
rect 88060 -148990 88780 -148960
rect 88780 -148990 89560 -148960
rect 89560 -148990 90280 -148960
rect 90280 -148990 91060 -148960
rect 91060 -148990 91780 -148960
rect 91780 -148990 92560 -148960
rect 92560 -148990 93280 -148960
rect 93280 -148990 94060 -148960
rect 94060 -148990 94780 -148960
rect 94780 -148990 95560 -148960
rect 95560 -148990 96280 -148960
rect 96280 -148990 97060 -148960
rect 97060 -148990 97780 -148960
rect 97780 -148990 98560 -148960
rect 98560 -148990 99280 -148960
rect 99280 -148990 100060 -148960
rect 100060 -148990 100780 -148960
rect 100780 -148990 101560 -148960
rect 101560 -148990 102280 -148960
rect 102280 -148990 103060 -148960
rect 103060 -148990 103780 -148960
rect 103780 -148990 104560 -148960
rect 104560 -148990 105280 -148960
rect 105280 -148990 106060 -148960
rect 106060 -148990 106780 -148960
rect 106780 -148990 107560 -148960
rect 107560 -148990 108280 -148960
rect 108280 -148990 109060 -148960
rect 109060 -148990 109780 -148960
rect 109780 -148990 110560 -148960
rect 110560 -148990 111280 -148960
rect 111280 -148990 112060 -148960
rect 112060 -148990 112780 -148960
rect 112780 -148990 113560 -148960
rect 113560 -148990 114280 -148960
rect 114280 -148990 115060 -148960
rect 115060 -148990 115780 -148960
rect 115780 -148990 116560 -148960
rect 116560 -148990 117280 -148960
rect 117280 -148990 118060 -148960
rect 118060 -148990 118780 -148960
rect 118780 -148990 119560 -148960
rect 119560 -148990 120280 -148960
rect 120280 -148990 121060 -148960
rect 121060 -148990 121780 -148960
rect 121780 -148990 122560 -148960
rect 122560 -148990 123280 -148960
rect 123280 -148990 124060 -148960
rect 124060 -148990 124780 -148960
rect 124780 -148990 125560 -148960
rect 125560 -148990 126280 -148960
rect 126280 -148990 127060 -148960
rect 127060 -148990 127780 -148960
rect 127780 -148990 128560 -148960
rect 128560 -148990 129280 -148960
rect 129280 -148990 130060 -148960
rect 130060 -148990 130780 -148960
rect 130780 -148990 131560 -148960
rect 131560 -148990 132280 -148960
rect 132280 -148990 133060 -148960
rect 133060 -148990 133780 -148960
rect 133780 -148990 134560 -148960
rect 134560 -148990 135280 -148960
rect 135280 -148990 136060 -148960
rect 136060 -148990 136780 -148960
rect 136780 -148990 137560 -148960
rect 137560 -148990 138280 -148960
rect 138280 -148990 139060 -148960
rect 139060 -148990 139780 -148960
rect 139780 -148990 140560 -148960
rect 140560 -148990 141280 -148960
rect 141280 -148990 142060 -148960
rect 142060 -148990 142780 -148960
rect 142780 -148990 143560 -148960
rect 143560 -148990 144280 -148960
rect 144280 -148990 145060 -148960
rect 145060 -148990 145780 -148960
rect 145780 -148990 146560 -148960
rect 146560 -148990 147280 -148960
rect 147280 -148990 148060 -148960
rect 148060 -148990 148780 -148960
rect 148780 -148990 149560 -148960
rect 149560 -148990 150370 -148960
rect 280 -149040 150370 -148990
<< metal2 >>
rect 0 2020 150000 2075
rect -1500 1725 -445 1730
rect -1500 1680 -960 1725
rect -450 1680 -445 1725
rect -1500 1675 -445 1680
rect -1500 780 -500 785
rect -1500 745 -790 780
rect -590 745 -500 780
rect -1500 740 -500 745
rect -375 115 -320 2000
rect 240 1825 295 1830
rect 240 1780 245 1825
rect 290 1780 295 1825
rect 240 1775 295 1780
rect 20 1725 75 1730
rect 20 1680 25 1725
rect 70 1680 75 1725
rect 20 1675 75 1680
rect 30 1500 65 1675
rect 250 1500 285 1775
rect 510 1500 545 2020
rect 1740 1825 1795 1830
rect 1740 1780 1745 1825
rect 1790 1780 1795 1825
rect 1740 1775 1795 1780
rect 1520 1725 1575 1730
rect 1520 1680 1525 1725
rect 1570 1680 1575 1725
rect 1520 1675 1575 1680
rect 1530 1500 1565 1675
rect 1750 1500 1785 1775
rect 2010 1500 2045 2020
rect 3240 1825 3295 1830
rect 3240 1780 3245 1825
rect 3290 1780 3295 1825
rect 3240 1775 3295 1780
rect 3020 1725 3075 1730
rect 3020 1680 3025 1725
rect 3070 1680 3075 1725
rect 3020 1675 3075 1680
rect 3030 1500 3065 1675
rect 3250 1500 3285 1775
rect 3510 1500 3545 2020
rect 4740 1825 4795 1830
rect 4740 1780 4745 1825
rect 4790 1780 4795 1825
rect 4740 1775 4795 1780
rect 4520 1725 4575 1730
rect 4520 1680 4525 1725
rect 4570 1680 4575 1725
rect 4520 1675 4575 1680
rect 4530 1500 4565 1675
rect 4750 1500 4785 1775
rect 5010 1500 5045 2020
rect 6240 1825 6295 1830
rect 6240 1780 6245 1825
rect 6290 1780 6295 1825
rect 6240 1775 6295 1780
rect 6020 1725 6075 1730
rect 6020 1680 6025 1725
rect 6070 1680 6075 1725
rect 6020 1675 6075 1680
rect 6030 1500 6065 1675
rect 6250 1500 6285 1775
rect 6510 1500 6545 2020
rect 7740 1825 7795 1830
rect 7740 1780 7745 1825
rect 7790 1780 7795 1825
rect 7740 1775 7795 1780
rect 7520 1725 7575 1730
rect 7520 1680 7525 1725
rect 7570 1680 7575 1725
rect 7520 1675 7575 1680
rect 7530 1500 7565 1675
rect 7750 1500 7785 1775
rect 8010 1500 8045 2020
rect 9240 1825 9295 1830
rect 9240 1780 9245 1825
rect 9290 1780 9295 1825
rect 9240 1775 9295 1780
rect 9020 1725 9075 1730
rect 9020 1680 9025 1725
rect 9070 1680 9075 1725
rect 9020 1675 9075 1680
rect 9030 1500 9065 1675
rect 9250 1500 9285 1775
rect 9510 1500 9545 2020
rect 10740 1825 10795 1830
rect 10740 1780 10745 1825
rect 10790 1780 10795 1825
rect 10740 1775 10795 1780
rect 10520 1725 10575 1730
rect 10520 1680 10525 1725
rect 10570 1680 10575 1725
rect 10520 1675 10575 1680
rect 10530 1500 10565 1675
rect 10750 1500 10785 1775
rect 11010 1500 11045 2020
rect 12240 1825 12295 1830
rect 12240 1780 12245 1825
rect 12290 1780 12295 1825
rect 12240 1775 12295 1780
rect 12020 1725 12075 1730
rect 12020 1680 12025 1725
rect 12070 1680 12075 1725
rect 12020 1675 12075 1680
rect 12030 1500 12065 1675
rect 12250 1500 12285 1775
rect 12510 1500 12545 2020
rect 13740 1825 13795 1830
rect 13740 1780 13745 1825
rect 13790 1780 13795 1825
rect 13740 1775 13795 1780
rect 13520 1725 13575 1730
rect 13520 1680 13525 1725
rect 13570 1680 13575 1725
rect 13520 1675 13575 1680
rect 13530 1500 13565 1675
rect 13750 1500 13785 1775
rect 14010 1500 14045 2020
rect 15240 1825 15295 1830
rect 15240 1780 15245 1825
rect 15290 1780 15295 1825
rect 15240 1775 15295 1780
rect 15020 1725 15075 1730
rect 15020 1680 15025 1725
rect 15070 1680 15075 1725
rect 15020 1675 15075 1680
rect 15030 1500 15065 1675
rect 15250 1500 15285 1775
rect 15510 1500 15545 2020
rect 16740 1825 16795 1830
rect 16740 1780 16745 1825
rect 16790 1780 16795 1825
rect 16740 1775 16795 1780
rect 16520 1725 16575 1730
rect 16520 1680 16525 1725
rect 16570 1680 16575 1725
rect 16520 1675 16575 1680
rect 16530 1500 16565 1675
rect 16750 1500 16785 1775
rect 17010 1500 17045 2020
rect 18240 1825 18295 1830
rect 18240 1780 18245 1825
rect 18290 1780 18295 1825
rect 18240 1775 18295 1780
rect 18020 1725 18075 1730
rect 18020 1680 18025 1725
rect 18070 1680 18075 1725
rect 18020 1675 18075 1680
rect 18030 1500 18065 1675
rect 18250 1500 18285 1775
rect 18510 1500 18545 2020
rect 19740 1825 19795 1830
rect 19740 1780 19745 1825
rect 19790 1780 19795 1825
rect 19740 1775 19795 1780
rect 19520 1725 19575 1730
rect 19520 1680 19525 1725
rect 19570 1680 19575 1725
rect 19520 1675 19575 1680
rect 19530 1500 19565 1675
rect 19750 1500 19785 1775
rect 20010 1500 20045 2020
rect 21240 1825 21295 1830
rect 21240 1780 21245 1825
rect 21290 1780 21295 1825
rect 21240 1775 21295 1780
rect 21020 1725 21075 1730
rect 21020 1680 21025 1725
rect 21070 1680 21075 1725
rect 21020 1675 21075 1680
rect 21030 1500 21065 1675
rect 21250 1500 21285 1775
rect 21510 1500 21545 2020
rect 22740 1825 22795 1830
rect 22740 1780 22745 1825
rect 22790 1780 22795 1825
rect 22740 1775 22795 1780
rect 22520 1725 22575 1730
rect 22520 1680 22525 1725
rect 22570 1680 22575 1725
rect 22520 1675 22575 1680
rect 22530 1500 22565 1675
rect 22750 1500 22785 1775
rect 23010 1500 23045 2020
rect 24240 1825 24295 1830
rect 24240 1780 24245 1825
rect 24290 1780 24295 1825
rect 24240 1775 24295 1780
rect 24020 1725 24075 1730
rect 24020 1680 24025 1725
rect 24070 1680 24075 1725
rect 24020 1675 24075 1680
rect 24030 1500 24065 1675
rect 24250 1500 24285 1775
rect 24510 1500 24545 2020
rect 25740 1825 25795 1830
rect 25740 1780 25745 1825
rect 25790 1780 25795 1825
rect 25740 1775 25795 1780
rect 25520 1725 25575 1730
rect 25520 1680 25525 1725
rect 25570 1680 25575 1725
rect 25520 1675 25575 1680
rect 25530 1500 25565 1675
rect 25750 1500 25785 1775
rect 26010 1500 26045 2020
rect 27240 1825 27295 1830
rect 27240 1780 27245 1825
rect 27290 1780 27295 1825
rect 27240 1775 27295 1780
rect 27020 1725 27075 1730
rect 27020 1680 27025 1725
rect 27070 1680 27075 1725
rect 27020 1675 27075 1680
rect 27030 1500 27065 1675
rect 27250 1500 27285 1775
rect 27510 1500 27545 2020
rect 28740 1825 28795 1830
rect 28740 1780 28745 1825
rect 28790 1780 28795 1825
rect 28740 1775 28795 1780
rect 28520 1725 28575 1730
rect 28520 1680 28525 1725
rect 28570 1680 28575 1725
rect 28520 1675 28575 1680
rect 28530 1500 28565 1675
rect 28750 1500 28785 1775
rect 29010 1500 29045 2020
rect 30240 1825 30295 1830
rect 30240 1780 30245 1825
rect 30290 1780 30295 1825
rect 30240 1775 30295 1780
rect 30020 1725 30075 1730
rect 30020 1680 30025 1725
rect 30070 1680 30075 1725
rect 30020 1675 30075 1680
rect 30030 1500 30065 1675
rect 30250 1500 30285 1775
rect 30510 1500 30545 2020
rect 31740 1825 31795 1830
rect 31740 1780 31745 1825
rect 31790 1780 31795 1825
rect 31740 1775 31795 1780
rect 31520 1725 31575 1730
rect 31520 1680 31525 1725
rect 31570 1680 31575 1725
rect 31520 1675 31575 1680
rect 31530 1500 31565 1675
rect 31750 1500 31785 1775
rect 32010 1500 32045 2020
rect 33240 1825 33295 1830
rect 33240 1780 33245 1825
rect 33290 1780 33295 1825
rect 33240 1775 33295 1780
rect 33020 1725 33075 1730
rect 33020 1680 33025 1725
rect 33070 1680 33075 1725
rect 33020 1675 33075 1680
rect 33030 1500 33065 1675
rect 33250 1500 33285 1775
rect 33510 1500 33545 2020
rect 34740 1825 34795 1830
rect 34740 1780 34745 1825
rect 34790 1780 34795 1825
rect 34740 1775 34795 1780
rect 34520 1725 34575 1730
rect 34520 1680 34525 1725
rect 34570 1680 34575 1725
rect 34520 1675 34575 1680
rect 34530 1500 34565 1675
rect 34750 1500 34785 1775
rect 35010 1500 35045 2020
rect 36240 1825 36295 1830
rect 36240 1780 36245 1825
rect 36290 1780 36295 1825
rect 36240 1775 36295 1780
rect 36020 1725 36075 1730
rect 36020 1680 36025 1725
rect 36070 1680 36075 1725
rect 36020 1675 36075 1680
rect 36030 1500 36065 1675
rect 36250 1500 36285 1775
rect 36510 1500 36545 2020
rect 37740 1825 37795 1830
rect 37740 1780 37745 1825
rect 37790 1780 37795 1825
rect 37740 1775 37795 1780
rect 37520 1725 37575 1730
rect 37520 1680 37525 1725
rect 37570 1680 37575 1725
rect 37520 1675 37575 1680
rect 37530 1500 37565 1675
rect 37750 1500 37785 1775
rect 38010 1500 38045 2020
rect 39240 1825 39295 1830
rect 39240 1780 39245 1825
rect 39290 1780 39295 1825
rect 39240 1775 39295 1780
rect 39020 1725 39075 1730
rect 39020 1680 39025 1725
rect 39070 1680 39075 1725
rect 39020 1675 39075 1680
rect 39030 1500 39065 1675
rect 39250 1500 39285 1775
rect 39510 1500 39545 2020
rect 40740 1825 40795 1830
rect 40740 1780 40745 1825
rect 40790 1780 40795 1825
rect 40740 1775 40795 1780
rect 40520 1725 40575 1730
rect 40520 1680 40525 1725
rect 40570 1680 40575 1725
rect 40520 1675 40575 1680
rect 40530 1500 40565 1675
rect 40750 1500 40785 1775
rect 41010 1500 41045 2020
rect 42240 1825 42295 1830
rect 42240 1780 42245 1825
rect 42290 1780 42295 1825
rect 42240 1775 42295 1780
rect 42020 1725 42075 1730
rect 42020 1680 42025 1725
rect 42070 1680 42075 1725
rect 42020 1675 42075 1680
rect 42030 1500 42065 1675
rect 42250 1500 42285 1775
rect 42510 1500 42545 2020
rect 43740 1825 43795 1830
rect 43740 1780 43745 1825
rect 43790 1780 43795 1825
rect 43740 1775 43795 1780
rect 43520 1725 43575 1730
rect 43520 1680 43525 1725
rect 43570 1680 43575 1725
rect 43520 1675 43575 1680
rect 43530 1500 43565 1675
rect 43750 1500 43785 1775
rect 44010 1500 44045 2020
rect 45240 1825 45295 1830
rect 45240 1780 45245 1825
rect 45290 1780 45295 1825
rect 45240 1775 45295 1780
rect 45020 1725 45075 1730
rect 45020 1680 45025 1725
rect 45070 1680 45075 1725
rect 45020 1675 45075 1680
rect 45030 1500 45065 1675
rect 45250 1500 45285 1775
rect 45510 1500 45545 2020
rect 46740 1825 46795 1830
rect 46740 1780 46745 1825
rect 46790 1780 46795 1825
rect 46740 1775 46795 1780
rect 46520 1725 46575 1730
rect 46520 1680 46525 1725
rect 46570 1680 46575 1725
rect 46520 1675 46575 1680
rect 46530 1500 46565 1675
rect 46750 1500 46785 1775
rect 47010 1500 47045 2020
rect 48240 1825 48295 1830
rect 48240 1780 48245 1825
rect 48290 1780 48295 1825
rect 48240 1775 48295 1780
rect 48020 1725 48075 1730
rect 48020 1680 48025 1725
rect 48070 1680 48075 1725
rect 48020 1675 48075 1680
rect 48030 1500 48065 1675
rect 48250 1500 48285 1775
rect 48510 1500 48545 2020
rect 49740 1825 49795 1830
rect 49740 1780 49745 1825
rect 49790 1780 49795 1825
rect 49740 1775 49795 1780
rect 49520 1725 49575 1730
rect 49520 1680 49525 1725
rect 49570 1680 49575 1725
rect 49520 1675 49575 1680
rect 49530 1500 49565 1675
rect 49750 1500 49785 1775
rect 50010 1500 50045 2020
rect 51240 1825 51295 1830
rect 51240 1780 51245 1825
rect 51290 1780 51295 1825
rect 51240 1775 51295 1780
rect 51020 1725 51075 1730
rect 51020 1680 51025 1725
rect 51070 1680 51075 1725
rect 51020 1675 51075 1680
rect 51030 1500 51065 1675
rect 51250 1500 51285 1775
rect 51510 1500 51545 2020
rect 52740 1825 52795 1830
rect 52740 1780 52745 1825
rect 52790 1780 52795 1825
rect 52740 1775 52795 1780
rect 52520 1725 52575 1730
rect 52520 1680 52525 1725
rect 52570 1680 52575 1725
rect 52520 1675 52575 1680
rect 52530 1500 52565 1675
rect 52750 1500 52785 1775
rect 53010 1500 53045 2020
rect 54240 1825 54295 1830
rect 54240 1780 54245 1825
rect 54290 1780 54295 1825
rect 54240 1775 54295 1780
rect 54020 1725 54075 1730
rect 54020 1680 54025 1725
rect 54070 1680 54075 1725
rect 54020 1675 54075 1680
rect 54030 1500 54065 1675
rect 54250 1500 54285 1775
rect 54510 1500 54545 2020
rect 55740 1825 55795 1830
rect 55740 1780 55745 1825
rect 55790 1780 55795 1825
rect 55740 1775 55795 1780
rect 55520 1725 55575 1730
rect 55520 1680 55525 1725
rect 55570 1680 55575 1725
rect 55520 1675 55575 1680
rect 55530 1500 55565 1675
rect 55750 1500 55785 1775
rect 56010 1500 56045 2020
rect 57240 1825 57295 1830
rect 57240 1780 57245 1825
rect 57290 1780 57295 1825
rect 57240 1775 57295 1780
rect 57020 1725 57075 1730
rect 57020 1680 57025 1725
rect 57070 1680 57075 1725
rect 57020 1675 57075 1680
rect 57030 1500 57065 1675
rect 57250 1500 57285 1775
rect 57510 1500 57545 2020
rect 58740 1825 58795 1830
rect 58740 1780 58745 1825
rect 58790 1780 58795 1825
rect 58740 1775 58795 1780
rect 58520 1725 58575 1730
rect 58520 1680 58525 1725
rect 58570 1680 58575 1725
rect 58520 1675 58575 1680
rect 58530 1500 58565 1675
rect 58750 1500 58785 1775
rect 59010 1500 59045 2020
rect 60240 1825 60295 1830
rect 60240 1780 60245 1825
rect 60290 1780 60295 1825
rect 60240 1775 60295 1780
rect 60020 1725 60075 1730
rect 60020 1680 60025 1725
rect 60070 1680 60075 1725
rect 60020 1675 60075 1680
rect 60030 1500 60065 1675
rect 60250 1500 60285 1775
rect 60510 1500 60545 2020
rect 61740 1825 61795 1830
rect 61740 1780 61745 1825
rect 61790 1780 61795 1825
rect 61740 1775 61795 1780
rect 61520 1725 61575 1730
rect 61520 1680 61525 1725
rect 61570 1680 61575 1725
rect 61520 1675 61575 1680
rect 61530 1500 61565 1675
rect 61750 1500 61785 1775
rect 62010 1500 62045 2020
rect 63240 1825 63295 1830
rect 63240 1780 63245 1825
rect 63290 1780 63295 1825
rect 63240 1775 63295 1780
rect 63020 1725 63075 1730
rect 63020 1680 63025 1725
rect 63070 1680 63075 1725
rect 63020 1675 63075 1680
rect 63030 1500 63065 1675
rect 63250 1500 63285 1775
rect 63510 1500 63545 2020
rect 64740 1825 64795 1830
rect 64740 1780 64745 1825
rect 64790 1780 64795 1825
rect 64740 1775 64795 1780
rect 64520 1725 64575 1730
rect 64520 1680 64525 1725
rect 64570 1680 64575 1725
rect 64520 1675 64575 1680
rect 64530 1500 64565 1675
rect 64750 1500 64785 1775
rect 65010 1500 65045 2020
rect 66240 1825 66295 1830
rect 66240 1780 66245 1825
rect 66290 1780 66295 1825
rect 66240 1775 66295 1780
rect 66020 1725 66075 1730
rect 66020 1680 66025 1725
rect 66070 1680 66075 1725
rect 66020 1675 66075 1680
rect 66030 1500 66065 1675
rect 66250 1500 66285 1775
rect 66510 1500 66545 2020
rect 67740 1825 67795 1830
rect 67740 1780 67745 1825
rect 67790 1780 67795 1825
rect 67740 1775 67795 1780
rect 67520 1725 67575 1730
rect 67520 1680 67525 1725
rect 67570 1680 67575 1725
rect 67520 1675 67575 1680
rect 67530 1500 67565 1675
rect 67750 1500 67785 1775
rect 68010 1500 68045 2020
rect 69240 1825 69295 1830
rect 69240 1780 69245 1825
rect 69290 1780 69295 1825
rect 69240 1775 69295 1780
rect 69020 1725 69075 1730
rect 69020 1680 69025 1725
rect 69070 1680 69075 1725
rect 69020 1675 69075 1680
rect 69030 1500 69065 1675
rect 69250 1500 69285 1775
rect 69510 1500 69545 2020
rect 70740 1825 70795 1830
rect 70740 1780 70745 1825
rect 70790 1780 70795 1825
rect 70740 1775 70795 1780
rect 70520 1725 70575 1730
rect 70520 1680 70525 1725
rect 70570 1680 70575 1725
rect 70520 1675 70575 1680
rect 70530 1500 70565 1675
rect 70750 1500 70785 1775
rect 71010 1500 71045 2020
rect 72240 1825 72295 1830
rect 72240 1780 72245 1825
rect 72290 1780 72295 1825
rect 72240 1775 72295 1780
rect 72020 1725 72075 1730
rect 72020 1680 72025 1725
rect 72070 1680 72075 1725
rect 72020 1675 72075 1680
rect 72030 1500 72065 1675
rect 72250 1500 72285 1775
rect 72510 1500 72545 2020
rect 73740 1825 73795 1830
rect 73740 1780 73745 1825
rect 73790 1780 73795 1825
rect 73740 1775 73795 1780
rect 73520 1725 73575 1730
rect 73520 1680 73525 1725
rect 73570 1680 73575 1725
rect 73520 1675 73575 1680
rect 73530 1500 73565 1675
rect 73750 1500 73785 1775
rect 74010 1500 74045 2020
rect 75240 1825 75295 1830
rect 75240 1780 75245 1825
rect 75290 1780 75295 1825
rect 75240 1775 75295 1780
rect 75020 1725 75075 1730
rect 75020 1680 75025 1725
rect 75070 1680 75075 1725
rect 75020 1675 75075 1680
rect 75030 1500 75065 1675
rect 75250 1500 75285 1775
rect 75510 1500 75545 2020
rect 76740 1825 76795 1830
rect 76740 1780 76745 1825
rect 76790 1780 76795 1825
rect 76740 1775 76795 1780
rect 76520 1725 76575 1730
rect 76520 1680 76525 1725
rect 76570 1680 76575 1725
rect 76520 1675 76575 1680
rect 76530 1500 76565 1675
rect 76750 1500 76785 1775
rect 77010 1500 77045 2020
rect 78240 1825 78295 1830
rect 78240 1780 78245 1825
rect 78290 1780 78295 1825
rect 78240 1775 78295 1780
rect 78020 1725 78075 1730
rect 78020 1680 78025 1725
rect 78070 1680 78075 1725
rect 78020 1675 78075 1680
rect 78030 1500 78065 1675
rect 78250 1500 78285 1775
rect 78510 1500 78545 2020
rect 79740 1825 79795 1830
rect 79740 1780 79745 1825
rect 79790 1780 79795 1825
rect 79740 1775 79795 1780
rect 79520 1725 79575 1730
rect 79520 1680 79525 1725
rect 79570 1680 79575 1725
rect 79520 1675 79575 1680
rect 79530 1500 79565 1675
rect 79750 1500 79785 1775
rect 80010 1500 80045 2020
rect 81240 1825 81295 1830
rect 81240 1780 81245 1825
rect 81290 1780 81295 1825
rect 81240 1775 81295 1780
rect 81020 1725 81075 1730
rect 81020 1680 81025 1725
rect 81070 1680 81075 1725
rect 81020 1675 81075 1680
rect 81030 1500 81065 1675
rect 81250 1500 81285 1775
rect 81510 1500 81545 2020
rect 82740 1825 82795 1830
rect 82740 1780 82745 1825
rect 82790 1780 82795 1825
rect 82740 1775 82795 1780
rect 82520 1725 82575 1730
rect 82520 1680 82525 1725
rect 82570 1680 82575 1725
rect 82520 1675 82575 1680
rect 82530 1500 82565 1675
rect 82750 1500 82785 1775
rect 83010 1500 83045 2020
rect 84240 1825 84295 1830
rect 84240 1780 84245 1825
rect 84290 1780 84295 1825
rect 84240 1775 84295 1780
rect 84020 1725 84075 1730
rect 84020 1680 84025 1725
rect 84070 1680 84075 1725
rect 84020 1675 84075 1680
rect 84030 1500 84065 1675
rect 84250 1500 84285 1775
rect 84510 1500 84545 2020
rect 85740 1825 85795 1830
rect 85740 1780 85745 1825
rect 85790 1780 85795 1825
rect 85740 1775 85795 1780
rect 85520 1725 85575 1730
rect 85520 1680 85525 1725
rect 85570 1680 85575 1725
rect 85520 1675 85575 1680
rect 85530 1500 85565 1675
rect 85750 1500 85785 1775
rect 86010 1500 86045 2020
rect 87240 1825 87295 1830
rect 87240 1780 87245 1825
rect 87290 1780 87295 1825
rect 87240 1775 87295 1780
rect 87020 1725 87075 1730
rect 87020 1680 87025 1725
rect 87070 1680 87075 1725
rect 87020 1675 87075 1680
rect 87030 1500 87065 1675
rect 87250 1500 87285 1775
rect 87510 1500 87545 2020
rect 88740 1825 88795 1830
rect 88740 1780 88745 1825
rect 88790 1780 88795 1825
rect 88740 1775 88795 1780
rect 88520 1725 88575 1730
rect 88520 1680 88525 1725
rect 88570 1680 88575 1725
rect 88520 1675 88575 1680
rect 88530 1500 88565 1675
rect 88750 1500 88785 1775
rect 89010 1500 89045 2020
rect 90240 1825 90295 1830
rect 90240 1780 90245 1825
rect 90290 1780 90295 1825
rect 90240 1775 90295 1780
rect 90020 1725 90075 1730
rect 90020 1680 90025 1725
rect 90070 1680 90075 1725
rect 90020 1675 90075 1680
rect 90030 1500 90065 1675
rect 90250 1500 90285 1775
rect 90510 1500 90545 2020
rect 91740 1825 91795 1830
rect 91740 1780 91745 1825
rect 91790 1780 91795 1825
rect 91740 1775 91795 1780
rect 91520 1725 91575 1730
rect 91520 1680 91525 1725
rect 91570 1680 91575 1725
rect 91520 1675 91575 1680
rect 91530 1500 91565 1675
rect 91750 1500 91785 1775
rect 92010 1500 92045 2020
rect 93240 1825 93295 1830
rect 93240 1780 93245 1825
rect 93290 1780 93295 1825
rect 93240 1775 93295 1780
rect 93020 1725 93075 1730
rect 93020 1680 93025 1725
rect 93070 1680 93075 1725
rect 93020 1675 93075 1680
rect 93030 1500 93065 1675
rect 93250 1500 93285 1775
rect 93510 1500 93545 2020
rect 94740 1825 94795 1830
rect 94740 1780 94745 1825
rect 94790 1780 94795 1825
rect 94740 1775 94795 1780
rect 94520 1725 94575 1730
rect 94520 1680 94525 1725
rect 94570 1680 94575 1725
rect 94520 1675 94575 1680
rect 94530 1500 94565 1675
rect 94750 1500 94785 1775
rect 95010 1500 95045 2020
rect 96240 1825 96295 1830
rect 96240 1780 96245 1825
rect 96290 1780 96295 1825
rect 96240 1775 96295 1780
rect 96020 1725 96075 1730
rect 96020 1680 96025 1725
rect 96070 1680 96075 1725
rect 96020 1675 96075 1680
rect 96030 1500 96065 1675
rect 96250 1500 96285 1775
rect 96510 1500 96545 2020
rect 97740 1825 97795 1830
rect 97740 1780 97745 1825
rect 97790 1780 97795 1825
rect 97740 1775 97795 1780
rect 97520 1725 97575 1730
rect 97520 1680 97525 1725
rect 97570 1680 97575 1725
rect 97520 1675 97575 1680
rect 97530 1500 97565 1675
rect 97750 1500 97785 1775
rect 98010 1500 98045 2020
rect 99240 1825 99295 1830
rect 99240 1780 99245 1825
rect 99290 1780 99295 1825
rect 99240 1775 99295 1780
rect 99020 1725 99075 1730
rect 99020 1680 99025 1725
rect 99070 1680 99075 1725
rect 99020 1675 99075 1680
rect 99030 1500 99065 1675
rect 99250 1500 99285 1775
rect 99510 1500 99545 2020
rect 100740 1825 100795 1830
rect 100740 1780 100745 1825
rect 100790 1780 100795 1825
rect 100740 1775 100795 1780
rect 100520 1725 100575 1730
rect 100520 1680 100525 1725
rect 100570 1680 100575 1725
rect 100520 1675 100575 1680
rect 100530 1500 100565 1675
rect 100750 1500 100785 1775
rect 101010 1500 101045 2020
rect 102240 1825 102295 1830
rect 102240 1780 102245 1825
rect 102290 1780 102295 1825
rect 102240 1775 102295 1780
rect 102020 1725 102075 1730
rect 102020 1680 102025 1725
rect 102070 1680 102075 1725
rect 102020 1675 102075 1680
rect 102030 1500 102065 1675
rect 102250 1500 102285 1775
rect 102510 1500 102545 2020
rect 103740 1825 103795 1830
rect 103740 1780 103745 1825
rect 103790 1780 103795 1825
rect 103740 1775 103795 1780
rect 103520 1725 103575 1730
rect 103520 1680 103525 1725
rect 103570 1680 103575 1725
rect 103520 1675 103575 1680
rect 103530 1500 103565 1675
rect 103750 1500 103785 1775
rect 104010 1500 104045 2020
rect 105240 1825 105295 1830
rect 105240 1780 105245 1825
rect 105290 1780 105295 1825
rect 105240 1775 105295 1780
rect 105020 1725 105075 1730
rect 105020 1680 105025 1725
rect 105070 1680 105075 1725
rect 105020 1675 105075 1680
rect 105030 1500 105065 1675
rect 105250 1500 105285 1775
rect 105510 1500 105545 2020
rect 106740 1825 106795 1830
rect 106740 1780 106745 1825
rect 106790 1780 106795 1825
rect 106740 1775 106795 1780
rect 106520 1725 106575 1730
rect 106520 1680 106525 1725
rect 106570 1680 106575 1725
rect 106520 1675 106575 1680
rect 106530 1500 106565 1675
rect 106750 1500 106785 1775
rect 107010 1500 107045 2020
rect 108240 1825 108295 1830
rect 108240 1780 108245 1825
rect 108290 1780 108295 1825
rect 108240 1775 108295 1780
rect 108020 1725 108075 1730
rect 108020 1680 108025 1725
rect 108070 1680 108075 1725
rect 108020 1675 108075 1680
rect 108030 1500 108065 1675
rect 108250 1500 108285 1775
rect 108510 1500 108545 2020
rect 109740 1825 109795 1830
rect 109740 1780 109745 1825
rect 109790 1780 109795 1825
rect 109740 1775 109795 1780
rect 109520 1725 109575 1730
rect 109520 1680 109525 1725
rect 109570 1680 109575 1725
rect 109520 1675 109575 1680
rect 109530 1500 109565 1675
rect 109750 1500 109785 1775
rect 110010 1500 110045 2020
rect 111240 1825 111295 1830
rect 111240 1780 111245 1825
rect 111290 1780 111295 1825
rect 111240 1775 111295 1780
rect 111020 1725 111075 1730
rect 111020 1680 111025 1725
rect 111070 1680 111075 1725
rect 111020 1675 111075 1680
rect 111030 1500 111065 1675
rect 111250 1500 111285 1775
rect 111510 1500 111545 2020
rect 112740 1825 112795 1830
rect 112740 1780 112745 1825
rect 112790 1780 112795 1825
rect 112740 1775 112795 1780
rect 112520 1725 112575 1730
rect 112520 1680 112525 1725
rect 112570 1680 112575 1725
rect 112520 1675 112575 1680
rect 112530 1500 112565 1675
rect 112750 1500 112785 1775
rect 113010 1500 113045 2020
rect 114240 1825 114295 1830
rect 114240 1780 114245 1825
rect 114290 1780 114295 1825
rect 114240 1775 114295 1780
rect 114020 1725 114075 1730
rect 114020 1680 114025 1725
rect 114070 1680 114075 1725
rect 114020 1675 114075 1680
rect 114030 1500 114065 1675
rect 114250 1500 114285 1775
rect 114510 1500 114545 2020
rect 115740 1825 115795 1830
rect 115740 1780 115745 1825
rect 115790 1780 115795 1825
rect 115740 1775 115795 1780
rect 115520 1725 115575 1730
rect 115520 1680 115525 1725
rect 115570 1680 115575 1725
rect 115520 1675 115575 1680
rect 115530 1500 115565 1675
rect 115750 1500 115785 1775
rect 116010 1500 116045 2020
rect 117240 1825 117295 1830
rect 117240 1780 117245 1825
rect 117290 1780 117295 1825
rect 117240 1775 117295 1780
rect 117020 1725 117075 1730
rect 117020 1680 117025 1725
rect 117070 1680 117075 1725
rect 117020 1675 117075 1680
rect 117030 1500 117065 1675
rect 117250 1500 117285 1775
rect 117510 1500 117545 2020
rect 118740 1825 118795 1830
rect 118740 1780 118745 1825
rect 118790 1780 118795 1825
rect 118740 1775 118795 1780
rect 118520 1725 118575 1730
rect 118520 1680 118525 1725
rect 118570 1680 118575 1725
rect 118520 1675 118575 1680
rect 118530 1500 118565 1675
rect 118750 1500 118785 1775
rect 119010 1500 119045 2020
rect 120240 1825 120295 1830
rect 120240 1780 120245 1825
rect 120290 1780 120295 1825
rect 120240 1775 120295 1780
rect 120020 1725 120075 1730
rect 120020 1680 120025 1725
rect 120070 1680 120075 1725
rect 120020 1675 120075 1680
rect 120030 1500 120065 1675
rect 120250 1500 120285 1775
rect 120510 1500 120545 2020
rect 121740 1825 121795 1830
rect 121740 1780 121745 1825
rect 121790 1780 121795 1825
rect 121740 1775 121795 1780
rect 121520 1725 121575 1730
rect 121520 1680 121525 1725
rect 121570 1680 121575 1725
rect 121520 1675 121575 1680
rect 121530 1500 121565 1675
rect 121750 1500 121785 1775
rect 122010 1500 122045 2020
rect 123240 1825 123295 1830
rect 123240 1780 123245 1825
rect 123290 1780 123295 1825
rect 123240 1775 123295 1780
rect 123020 1725 123075 1730
rect 123020 1680 123025 1725
rect 123070 1680 123075 1725
rect 123020 1675 123075 1680
rect 123030 1500 123065 1675
rect 123250 1500 123285 1775
rect 123510 1500 123545 2020
rect 124740 1825 124795 1830
rect 124740 1780 124745 1825
rect 124790 1780 124795 1825
rect 124740 1775 124795 1780
rect 124520 1725 124575 1730
rect 124520 1680 124525 1725
rect 124570 1680 124575 1725
rect 124520 1675 124575 1680
rect 124530 1500 124565 1675
rect 124750 1500 124785 1775
rect 125010 1500 125045 2020
rect 126240 1825 126295 1830
rect 126240 1780 126245 1825
rect 126290 1780 126295 1825
rect 126240 1775 126295 1780
rect 126020 1725 126075 1730
rect 126020 1680 126025 1725
rect 126070 1680 126075 1725
rect 126020 1675 126075 1680
rect 126030 1500 126065 1675
rect 126250 1500 126285 1775
rect 126510 1500 126545 2020
rect 127740 1825 127795 1830
rect 127740 1780 127745 1825
rect 127790 1780 127795 1825
rect 127740 1775 127795 1780
rect 127520 1725 127575 1730
rect 127520 1680 127525 1725
rect 127570 1680 127575 1725
rect 127520 1675 127575 1680
rect 127530 1500 127565 1675
rect 127750 1500 127785 1775
rect 128010 1500 128045 2020
rect 129240 1825 129295 1830
rect 129240 1780 129245 1825
rect 129290 1780 129295 1825
rect 129240 1775 129295 1780
rect 129020 1725 129075 1730
rect 129020 1680 129025 1725
rect 129070 1680 129075 1725
rect 129020 1675 129075 1680
rect 129030 1500 129065 1675
rect 129250 1500 129285 1775
rect 129510 1500 129545 2020
rect 130740 1825 130795 1830
rect 130740 1780 130745 1825
rect 130790 1780 130795 1825
rect 130740 1775 130795 1780
rect 130520 1725 130575 1730
rect 130520 1680 130525 1725
rect 130570 1680 130575 1725
rect 130520 1675 130575 1680
rect 130530 1500 130565 1675
rect 130750 1500 130785 1775
rect 131010 1500 131045 2020
rect 132240 1825 132295 1830
rect 132240 1780 132245 1825
rect 132290 1780 132295 1825
rect 132240 1775 132295 1780
rect 132020 1725 132075 1730
rect 132020 1680 132025 1725
rect 132070 1680 132075 1725
rect 132020 1675 132075 1680
rect 132030 1500 132065 1675
rect 132250 1500 132285 1775
rect 132510 1500 132545 2020
rect 133740 1825 133795 1830
rect 133740 1780 133745 1825
rect 133790 1780 133795 1825
rect 133740 1775 133795 1780
rect 133520 1725 133575 1730
rect 133520 1680 133525 1725
rect 133570 1680 133575 1725
rect 133520 1675 133575 1680
rect 133530 1500 133565 1675
rect 133750 1500 133785 1775
rect 134010 1500 134045 2020
rect 135240 1825 135295 1830
rect 135240 1780 135245 1825
rect 135290 1780 135295 1825
rect 135240 1775 135295 1780
rect 135020 1725 135075 1730
rect 135020 1680 135025 1725
rect 135070 1680 135075 1725
rect 135020 1675 135075 1680
rect 135030 1500 135065 1675
rect 135250 1500 135285 1775
rect 135510 1500 135545 2020
rect 136740 1825 136795 1830
rect 136740 1780 136745 1825
rect 136790 1780 136795 1825
rect 136740 1775 136795 1780
rect 136520 1725 136575 1730
rect 136520 1680 136525 1725
rect 136570 1680 136575 1725
rect 136520 1675 136575 1680
rect 136530 1500 136565 1675
rect 136750 1500 136785 1775
rect 137010 1500 137045 2020
rect 138240 1825 138295 1830
rect 138240 1780 138245 1825
rect 138290 1780 138295 1825
rect 138240 1775 138295 1780
rect 138020 1725 138075 1730
rect 138020 1680 138025 1725
rect 138070 1680 138075 1725
rect 138020 1675 138075 1680
rect 138030 1500 138065 1675
rect 138250 1500 138285 1775
rect 138510 1500 138545 2020
rect 139740 1825 139795 1830
rect 139740 1780 139745 1825
rect 139790 1780 139795 1825
rect 139740 1775 139795 1780
rect 139520 1725 139575 1730
rect 139520 1680 139525 1725
rect 139570 1680 139575 1725
rect 139520 1675 139575 1680
rect 139530 1500 139565 1675
rect 139750 1500 139785 1775
rect 140010 1500 140045 2020
rect 141240 1825 141295 1830
rect 141240 1780 141245 1825
rect 141290 1780 141295 1825
rect 141240 1775 141295 1780
rect 141020 1725 141075 1730
rect 141020 1680 141025 1725
rect 141070 1680 141075 1725
rect 141020 1675 141075 1680
rect 141030 1500 141065 1675
rect 141250 1500 141285 1775
rect 141510 1500 141545 2020
rect 142740 1825 142795 1830
rect 142740 1780 142745 1825
rect 142790 1780 142795 1825
rect 142740 1775 142795 1780
rect 142520 1725 142575 1730
rect 142520 1680 142525 1725
rect 142570 1680 142575 1725
rect 142520 1675 142575 1680
rect 142530 1500 142565 1675
rect 142750 1500 142785 1775
rect 143010 1500 143045 2020
rect 144240 1825 144295 1830
rect 144240 1780 144245 1825
rect 144290 1780 144295 1825
rect 144240 1775 144295 1780
rect 144020 1725 144075 1730
rect 144020 1680 144025 1725
rect 144070 1680 144075 1725
rect 144020 1675 144075 1680
rect 144030 1500 144065 1675
rect 144250 1500 144285 1775
rect 144510 1500 144545 2020
rect 145740 1825 145795 1830
rect 145740 1780 145745 1825
rect 145790 1780 145795 1825
rect 145740 1775 145795 1780
rect 145520 1725 145575 1730
rect 145520 1680 145525 1725
rect 145570 1680 145575 1725
rect 145520 1675 145575 1680
rect 145530 1500 145565 1675
rect 145750 1500 145785 1775
rect 146010 1500 146045 2020
rect 147240 1825 147295 1830
rect 147240 1780 147245 1825
rect 147290 1780 147295 1825
rect 147240 1775 147295 1780
rect 147020 1725 147075 1730
rect 147020 1680 147025 1725
rect 147070 1680 147075 1725
rect 147020 1675 147075 1680
rect 147030 1500 147065 1675
rect 147250 1500 147285 1775
rect 147510 1500 147545 2020
rect 148740 1825 148795 1830
rect 148740 1780 148745 1825
rect 148790 1780 148795 1825
rect 148740 1775 148795 1780
rect 148520 1725 148575 1730
rect 148520 1680 148525 1725
rect 148570 1680 148575 1725
rect 148520 1675 148575 1680
rect 148530 1500 148565 1675
rect 148750 1500 148785 1775
rect 149010 1500 149045 2020
rect -280 780 -130 785
rect -280 745 -270 780
rect -280 740 -130 745
rect -375 80 -370 115
rect -325 80 -320 115
rect -1500 -720 -500 -715
rect -1500 -755 -790 -720
rect -590 -755 -500 -720
rect -1500 -760 -500 -755
rect -375 -1385 -320 80
rect -280 -720 -130 -715
rect -280 -755 -270 -720
rect -280 -760 -130 -755
rect -375 -1420 -370 -1385
rect -325 -1420 -320 -1385
rect -1500 -2220 -500 -2215
rect -1500 -2255 -790 -2220
rect -590 -2255 -500 -2220
rect -1500 -2260 -500 -2255
rect -375 -2885 -320 -1420
rect -280 -2220 -130 -2215
rect -280 -2255 -270 -2220
rect -280 -2260 -130 -2255
rect -375 -2920 -370 -2885
rect -325 -2920 -320 -2885
rect -1500 -3720 -500 -3715
rect -1500 -3755 -790 -3720
rect -590 -3755 -500 -3720
rect -1500 -3760 -500 -3755
rect -375 -4385 -320 -2920
rect -280 -3720 -130 -3715
rect -280 -3755 -270 -3720
rect -280 -3760 -130 -3755
rect -375 -4420 -370 -4385
rect -325 -4420 -320 -4385
rect -1500 -5220 -500 -5215
rect -1500 -5255 -790 -5220
rect -590 -5255 -500 -5220
rect -1500 -5260 -500 -5255
rect -375 -5885 -320 -4420
rect -280 -5220 -130 -5215
rect -280 -5255 -270 -5220
rect -280 -5260 -130 -5255
rect -375 -5920 -370 -5885
rect -325 -5920 -320 -5885
rect -1500 -6720 -500 -6715
rect -1500 -6755 -790 -6720
rect -590 -6755 -500 -6720
rect -1500 -6760 -500 -6755
rect -375 -7385 -320 -5920
rect -280 -6720 -130 -6715
rect -280 -6755 -270 -6720
rect -280 -6760 -130 -6755
rect -375 -7420 -370 -7385
rect -325 -7420 -320 -7385
rect -1500 -8220 -500 -8215
rect -1500 -8255 -790 -8220
rect -590 -8255 -500 -8220
rect -1500 -8260 -500 -8255
rect -375 -8885 -320 -7420
rect -280 -8220 -130 -8215
rect -280 -8255 -270 -8220
rect -280 -8260 -130 -8255
rect -375 -8920 -370 -8885
rect -325 -8920 -320 -8885
rect -1500 -9720 -500 -9715
rect -1500 -9755 -790 -9720
rect -590 -9755 -500 -9720
rect -1500 -9760 -500 -9755
rect -375 -10385 -320 -8920
rect -280 -9720 -130 -9715
rect -280 -9755 -270 -9720
rect -280 -9760 -130 -9755
rect -375 -10420 -370 -10385
rect -325 -10420 -320 -10385
rect -1500 -11220 -500 -11215
rect -1500 -11255 -790 -11220
rect -590 -11255 -500 -11220
rect -1500 -11260 -500 -11255
rect -375 -11885 -320 -10420
rect -280 -11220 -130 -11215
rect -280 -11255 -270 -11220
rect -280 -11260 -130 -11255
rect -375 -11920 -370 -11885
rect -325 -11920 -320 -11885
rect -1500 -12720 -500 -12715
rect -1500 -12755 -790 -12720
rect -590 -12755 -500 -12720
rect -1500 -12760 -500 -12755
rect -375 -13385 -320 -11920
rect -280 -12720 -130 -12715
rect -280 -12755 -270 -12720
rect -280 -12760 -130 -12755
rect -375 -13420 -370 -13385
rect -325 -13420 -320 -13385
rect -1500 -14220 -500 -14215
rect -1500 -14255 -790 -14220
rect -590 -14255 -500 -14220
rect -1500 -14260 -500 -14255
rect -375 -14885 -320 -13420
rect -280 -14220 -130 -14215
rect -280 -14255 -270 -14220
rect -280 -14260 -130 -14255
rect -375 -14920 -370 -14885
rect -325 -14920 -320 -14885
rect -1500 -15720 -500 -15715
rect -1500 -15755 -790 -15720
rect -590 -15755 -500 -15720
rect -1500 -15760 -500 -15755
rect -375 -16385 -320 -14920
rect -280 -15720 -130 -15715
rect -280 -15755 -270 -15720
rect -280 -15760 -130 -15755
rect -375 -16420 -370 -16385
rect -325 -16420 -320 -16385
rect -1500 -17220 -500 -17215
rect -1500 -17255 -790 -17220
rect -590 -17255 -500 -17220
rect -1500 -17260 -500 -17255
rect -375 -17885 -320 -16420
rect -280 -17220 -130 -17215
rect -280 -17255 -270 -17220
rect -280 -17260 -130 -17255
rect -375 -17920 -370 -17885
rect -325 -17920 -320 -17885
rect -1500 -18720 -500 -18715
rect -1500 -18755 -790 -18720
rect -590 -18755 -500 -18720
rect -1500 -18760 -500 -18755
rect -375 -19385 -320 -17920
rect -280 -18720 -130 -18715
rect -280 -18755 -270 -18720
rect -280 -18760 -130 -18755
rect -375 -19420 -370 -19385
rect -325 -19420 -320 -19385
rect -1500 -20220 -500 -20215
rect -1500 -20255 -790 -20220
rect -590 -20255 -500 -20220
rect -1500 -20260 -500 -20255
rect -375 -20885 -320 -19420
rect -280 -20220 -130 -20215
rect -280 -20255 -270 -20220
rect -280 -20260 -130 -20255
rect -375 -20920 -370 -20885
rect -325 -20920 -320 -20885
rect -1500 -21720 -500 -21715
rect -1500 -21755 -790 -21720
rect -590 -21755 -500 -21720
rect -1500 -21760 -500 -21755
rect -375 -22385 -320 -20920
rect -280 -21720 -130 -21715
rect -280 -21755 -270 -21720
rect -280 -21760 -130 -21755
rect -375 -22420 -370 -22385
rect -325 -22420 -320 -22385
rect -1500 -23220 -500 -23215
rect -1500 -23255 -790 -23220
rect -590 -23255 -500 -23220
rect -1500 -23260 -500 -23255
rect -375 -23885 -320 -22420
rect -280 -23220 -130 -23215
rect -280 -23255 -270 -23220
rect -280 -23260 -130 -23255
rect -375 -23920 -370 -23885
rect -325 -23920 -320 -23885
rect -1500 -24720 -500 -24715
rect -1500 -24755 -790 -24720
rect -590 -24755 -500 -24720
rect -1500 -24760 -500 -24755
rect -375 -25385 -320 -23920
rect -280 -24720 -130 -24715
rect -280 -24755 -270 -24720
rect -280 -24760 -130 -24755
rect -375 -25420 -370 -25385
rect -325 -25420 -320 -25385
rect -1500 -26220 -500 -26215
rect -1500 -26255 -790 -26220
rect -590 -26255 -500 -26220
rect -1500 -26260 -500 -26255
rect -375 -26885 -320 -25420
rect -280 -26220 -130 -26215
rect -280 -26255 -270 -26220
rect -280 -26260 -130 -26255
rect -375 -26920 -370 -26885
rect -325 -26920 -320 -26885
rect -1500 -27720 -500 -27715
rect -1500 -27755 -790 -27720
rect -590 -27755 -500 -27720
rect -1500 -27760 -500 -27755
rect -375 -28385 -320 -26920
rect -280 -27720 -130 -27715
rect -280 -27755 -270 -27720
rect -280 -27760 -130 -27755
rect -375 -28420 -370 -28385
rect -325 -28420 -320 -28385
rect -1500 -29220 -500 -29215
rect -1500 -29255 -790 -29220
rect -590 -29255 -500 -29220
rect -1500 -29260 -500 -29255
rect -375 -29885 -320 -28420
rect -280 -29220 -130 -29215
rect -280 -29255 -270 -29220
rect -280 -29260 -130 -29255
rect -375 -29920 -370 -29885
rect -325 -29920 -320 -29885
rect -1500 -30720 -500 -30715
rect -1500 -30755 -790 -30720
rect -590 -30755 -500 -30720
rect -1500 -30760 -500 -30755
rect -375 -31385 -320 -29920
rect -280 -30720 -130 -30715
rect -280 -30755 -270 -30720
rect -280 -30760 -130 -30755
rect -375 -31420 -370 -31385
rect -325 -31420 -320 -31385
rect -1500 -32220 -500 -32215
rect -1500 -32255 -790 -32220
rect -590 -32255 -500 -32220
rect -1500 -32260 -500 -32255
rect -375 -32885 -320 -31420
rect -280 -32220 -130 -32215
rect -280 -32255 -270 -32220
rect -280 -32260 -130 -32255
rect -375 -32920 -370 -32885
rect -325 -32920 -320 -32885
rect -1500 -33720 -500 -33715
rect -1500 -33755 -790 -33720
rect -590 -33755 -500 -33720
rect -1500 -33760 -500 -33755
rect -375 -34385 -320 -32920
rect -280 -33720 -130 -33715
rect -280 -33755 -270 -33720
rect -280 -33760 -130 -33755
rect -375 -34420 -370 -34385
rect -325 -34420 -320 -34385
rect -1500 -35220 -500 -35215
rect -1500 -35255 -790 -35220
rect -590 -35255 -500 -35220
rect -1500 -35260 -500 -35255
rect -375 -35885 -320 -34420
rect -280 -35220 -130 -35215
rect -280 -35255 -270 -35220
rect -280 -35260 -130 -35255
rect -375 -35920 -370 -35885
rect -325 -35920 -320 -35885
rect -1500 -36720 -500 -36715
rect -1500 -36755 -790 -36720
rect -590 -36755 -500 -36720
rect -1500 -36760 -500 -36755
rect -375 -37385 -320 -35920
rect -280 -36720 -130 -36715
rect -280 -36755 -270 -36720
rect -280 -36760 -130 -36755
rect -375 -37420 -370 -37385
rect -325 -37420 -320 -37385
rect -1500 -38220 -500 -38215
rect -1500 -38255 -790 -38220
rect -590 -38255 -500 -38220
rect -1500 -38260 -500 -38255
rect -375 -38885 -320 -37420
rect -280 -38220 -130 -38215
rect -280 -38255 -270 -38220
rect -280 -38260 -130 -38255
rect -375 -38920 -370 -38885
rect -325 -38920 -320 -38885
rect -1500 -39720 -500 -39715
rect -1500 -39755 -790 -39720
rect -590 -39755 -500 -39720
rect -1500 -39760 -500 -39755
rect -375 -40385 -320 -38920
rect -280 -39720 -130 -39715
rect -280 -39755 -270 -39720
rect -280 -39760 -130 -39755
rect -375 -40420 -370 -40385
rect -325 -40420 -320 -40385
rect -1500 -41220 -500 -41215
rect -1500 -41255 -790 -41220
rect -590 -41255 -500 -41220
rect -1500 -41260 -500 -41255
rect -375 -41885 -320 -40420
rect -280 -41220 -130 -41215
rect -280 -41255 -270 -41220
rect -280 -41260 -130 -41255
rect -375 -41920 -370 -41885
rect -325 -41920 -320 -41885
rect -1500 -42720 -500 -42715
rect -1500 -42755 -790 -42720
rect -590 -42755 -500 -42720
rect -1500 -42760 -500 -42755
rect -375 -43385 -320 -41920
rect -280 -42720 -130 -42715
rect -280 -42755 -270 -42720
rect -280 -42760 -130 -42755
rect -375 -43420 -370 -43385
rect -325 -43420 -320 -43385
rect -1500 -44220 -500 -44215
rect -1500 -44255 -790 -44220
rect -590 -44255 -500 -44220
rect -1500 -44260 -500 -44255
rect -375 -44885 -320 -43420
rect -280 -44220 -130 -44215
rect -280 -44255 -270 -44220
rect -280 -44260 -130 -44255
rect -375 -44920 -370 -44885
rect -325 -44920 -320 -44885
rect -1500 -45720 -500 -45715
rect -1500 -45755 -790 -45720
rect -590 -45755 -500 -45720
rect -1500 -45760 -500 -45755
rect -375 -46385 -320 -44920
rect -280 -45720 -130 -45715
rect -280 -45755 -270 -45720
rect -280 -45760 -130 -45755
rect -375 -46420 -370 -46385
rect -325 -46420 -320 -46385
rect -1500 -47220 -500 -47215
rect -1500 -47255 -790 -47220
rect -590 -47255 -500 -47220
rect -1500 -47260 -500 -47255
rect -375 -47885 -320 -46420
rect -280 -47220 -130 -47215
rect -280 -47255 -270 -47220
rect -280 -47260 -130 -47255
rect -375 -47920 -370 -47885
rect -325 -47920 -320 -47885
rect -1500 -48720 -500 -48715
rect -1500 -48755 -790 -48720
rect -590 -48755 -500 -48720
rect -1500 -48760 -500 -48755
rect -375 -49385 -320 -47920
rect -280 -48720 -130 -48715
rect -280 -48755 -270 -48720
rect -280 -48760 -130 -48755
rect -375 -49420 -370 -49385
rect -325 -49420 -320 -49385
rect -1500 -50220 -500 -50215
rect -1500 -50255 -790 -50220
rect -590 -50255 -500 -50220
rect -1500 -50260 -500 -50255
rect -375 -50885 -320 -49420
rect -280 -50220 -130 -50215
rect -280 -50255 -270 -50220
rect -280 -50260 -130 -50255
rect -375 -50920 -370 -50885
rect -325 -50920 -320 -50885
rect -1500 -51720 -500 -51715
rect -1500 -51755 -790 -51720
rect -590 -51755 -500 -51720
rect -1500 -51760 -500 -51755
rect -375 -52385 -320 -50920
rect -280 -51720 -130 -51715
rect -280 -51755 -270 -51720
rect -280 -51760 -130 -51755
rect -375 -52420 -370 -52385
rect -325 -52420 -320 -52385
rect -1500 -53220 -500 -53215
rect -1500 -53255 -790 -53220
rect -590 -53255 -500 -53220
rect -1500 -53260 -500 -53255
rect -375 -53885 -320 -52420
rect -280 -53220 -130 -53215
rect -280 -53255 -270 -53220
rect -280 -53260 -130 -53255
rect -375 -53920 -370 -53885
rect -325 -53920 -320 -53885
rect -1500 -54720 -500 -54715
rect -1500 -54755 -790 -54720
rect -590 -54755 -500 -54720
rect -1500 -54760 -500 -54755
rect -375 -55385 -320 -53920
rect -280 -54720 -130 -54715
rect -280 -54755 -270 -54720
rect -280 -54760 -130 -54755
rect -375 -55420 -370 -55385
rect -325 -55420 -320 -55385
rect -1500 -56220 -500 -56215
rect -1500 -56255 -790 -56220
rect -590 -56255 -500 -56220
rect -1500 -56260 -500 -56255
rect -375 -56885 -320 -55420
rect -280 -56220 -130 -56215
rect -280 -56255 -270 -56220
rect -280 -56260 -130 -56255
rect -375 -56920 -370 -56885
rect -325 -56920 -320 -56885
rect -1500 -57720 -500 -57715
rect -1500 -57755 -790 -57720
rect -590 -57755 -500 -57720
rect -1500 -57760 -500 -57755
rect -375 -58385 -320 -56920
rect -280 -57720 -130 -57715
rect -280 -57755 -270 -57720
rect -280 -57760 -130 -57755
rect -375 -58420 -370 -58385
rect -325 -58420 -320 -58385
rect -1500 -59220 -500 -59215
rect -1500 -59255 -790 -59220
rect -590 -59255 -500 -59220
rect -1500 -59260 -500 -59255
rect -375 -59885 -320 -58420
rect -280 -59220 -130 -59215
rect -280 -59255 -270 -59220
rect -280 -59260 -130 -59255
rect -375 -59920 -370 -59885
rect -325 -59920 -320 -59885
rect -1500 -60720 -500 -60715
rect -1500 -60755 -790 -60720
rect -590 -60755 -500 -60720
rect -1500 -60760 -500 -60755
rect -375 -61385 -320 -59920
rect -280 -60720 -130 -60715
rect -280 -60755 -270 -60720
rect -280 -60760 -130 -60755
rect -375 -61420 -370 -61385
rect -325 -61420 -320 -61385
rect -1500 -62220 -500 -62215
rect -1500 -62255 -790 -62220
rect -590 -62255 -500 -62220
rect -1500 -62260 -500 -62255
rect -375 -62885 -320 -61420
rect -280 -62220 -130 -62215
rect -280 -62255 -270 -62220
rect -280 -62260 -130 -62255
rect -375 -62920 -370 -62885
rect -325 -62920 -320 -62885
rect -1500 -63720 -500 -63715
rect -1500 -63755 -790 -63720
rect -590 -63755 -500 -63720
rect -1500 -63760 -500 -63755
rect -375 -64385 -320 -62920
rect -280 -63720 -130 -63715
rect -280 -63755 -270 -63720
rect -280 -63760 -130 -63755
rect -375 -64420 -370 -64385
rect -325 -64420 -320 -64385
rect -1500 -65220 -500 -65215
rect -1500 -65255 -790 -65220
rect -590 -65255 -500 -65220
rect -1500 -65260 -500 -65255
rect -375 -65885 -320 -64420
rect -280 -65220 -130 -65215
rect -280 -65255 -270 -65220
rect -280 -65260 -130 -65255
rect -375 -65920 -370 -65885
rect -325 -65920 -320 -65885
rect -1500 -66720 -500 -66715
rect -1500 -66755 -790 -66720
rect -590 -66755 -500 -66720
rect -1500 -66760 -500 -66755
rect -375 -67385 -320 -65920
rect -280 -66720 -130 -66715
rect -280 -66755 -270 -66720
rect -280 -66760 -130 -66755
rect -375 -67420 -370 -67385
rect -325 -67420 -320 -67385
rect -1500 -68220 -500 -68215
rect -1500 -68255 -790 -68220
rect -590 -68255 -500 -68220
rect -1500 -68260 -500 -68255
rect -375 -68885 -320 -67420
rect -280 -68220 -130 -68215
rect -280 -68255 -270 -68220
rect -280 -68260 -130 -68255
rect -375 -68920 -370 -68885
rect -325 -68920 -320 -68885
rect -1500 -69720 -500 -69715
rect -1500 -69755 -790 -69720
rect -590 -69755 -500 -69720
rect -1500 -69760 -500 -69755
rect -375 -70385 -320 -68920
rect -280 -69720 -130 -69715
rect -280 -69755 -270 -69720
rect -280 -69760 -130 -69755
rect -375 -70420 -370 -70385
rect -325 -70420 -320 -70385
rect -1500 -71220 -500 -71215
rect -1500 -71255 -790 -71220
rect -590 -71255 -500 -71220
rect -1500 -71260 -500 -71255
rect -375 -71885 -320 -70420
rect -280 -71220 -130 -71215
rect -280 -71255 -270 -71220
rect -280 -71260 -130 -71255
rect -375 -71920 -370 -71885
rect -325 -71920 -320 -71885
rect -1500 -72720 -500 -72715
rect -1500 -72755 -790 -72720
rect -590 -72755 -500 -72720
rect -1500 -72760 -500 -72755
rect -375 -73385 -320 -71920
rect -280 -72720 -130 -72715
rect -280 -72755 -270 -72720
rect -280 -72760 -130 -72755
rect -375 -73420 -370 -73385
rect -325 -73420 -320 -73385
rect -1500 -74220 -500 -74215
rect -1500 -74255 -790 -74220
rect -590 -74255 -500 -74220
rect -1500 -74260 -500 -74255
rect -375 -74885 -320 -73420
rect -280 -74220 -130 -74215
rect -280 -74255 -270 -74220
rect -280 -74260 -130 -74255
rect -375 -74920 -370 -74885
rect -325 -74920 -320 -74885
rect -1500 -75720 -500 -75715
rect -1500 -75755 -790 -75720
rect -590 -75755 -500 -75720
rect -1500 -75760 -500 -75755
rect -375 -76385 -320 -74920
rect -280 -75720 -130 -75715
rect -280 -75755 -270 -75720
rect -280 -75760 -130 -75755
rect -375 -76420 -370 -76385
rect -325 -76420 -320 -76385
rect -1500 -77220 -500 -77215
rect -1500 -77255 -790 -77220
rect -590 -77255 -500 -77220
rect -1500 -77260 -500 -77255
rect -375 -77885 -320 -76420
rect -280 -77220 -130 -77215
rect -280 -77255 -270 -77220
rect -280 -77260 -130 -77255
rect -375 -77920 -370 -77885
rect -325 -77920 -320 -77885
rect -1500 -78720 -500 -78715
rect -1500 -78755 -790 -78720
rect -590 -78755 -500 -78720
rect -1500 -78760 -500 -78755
rect -375 -79385 -320 -77920
rect -280 -78720 -130 -78715
rect -280 -78755 -270 -78720
rect -280 -78760 -130 -78755
rect -375 -79420 -370 -79385
rect -325 -79420 -320 -79385
rect -1500 -80220 -500 -80215
rect -1500 -80255 -790 -80220
rect -590 -80255 -500 -80220
rect -1500 -80260 -500 -80255
rect -375 -80885 -320 -79420
rect -280 -80220 -130 -80215
rect -280 -80255 -270 -80220
rect -280 -80260 -130 -80255
rect -375 -80920 -370 -80885
rect -325 -80920 -320 -80885
rect -1500 -81720 -500 -81715
rect -1500 -81755 -790 -81720
rect -590 -81755 -500 -81720
rect -1500 -81760 -500 -81755
rect -375 -82385 -320 -80920
rect -280 -81720 -130 -81715
rect -280 -81755 -270 -81720
rect -280 -81760 -130 -81755
rect -375 -82420 -370 -82385
rect -325 -82420 -320 -82385
rect -1500 -83220 -500 -83215
rect -1500 -83255 -790 -83220
rect -590 -83255 -500 -83220
rect -1500 -83260 -500 -83255
rect -375 -83885 -320 -82420
rect -280 -83220 -130 -83215
rect -280 -83255 -270 -83220
rect -280 -83260 -130 -83255
rect -375 -83920 -370 -83885
rect -325 -83920 -320 -83885
rect -1500 -84720 -500 -84715
rect -1500 -84755 -790 -84720
rect -590 -84755 -500 -84720
rect -1500 -84760 -500 -84755
rect -375 -85385 -320 -83920
rect -280 -84720 -130 -84715
rect -280 -84755 -270 -84720
rect -280 -84760 -130 -84755
rect -375 -85420 -370 -85385
rect -325 -85420 -320 -85385
rect -1500 -86220 -500 -86215
rect -1500 -86255 -790 -86220
rect -590 -86255 -500 -86220
rect -1500 -86260 -500 -86255
rect -375 -86885 -320 -85420
rect -280 -86220 -130 -86215
rect -280 -86255 -270 -86220
rect -280 -86260 -130 -86255
rect -375 -86920 -370 -86885
rect -325 -86920 -320 -86885
rect -1500 -87720 -500 -87715
rect -1500 -87755 -790 -87720
rect -590 -87755 -500 -87720
rect -1500 -87760 -500 -87755
rect -375 -88385 -320 -86920
rect -280 -87720 -130 -87715
rect -280 -87755 -270 -87720
rect -280 -87760 -130 -87755
rect -375 -88420 -370 -88385
rect -325 -88420 -320 -88385
rect -1500 -89220 -500 -89215
rect -1500 -89255 -790 -89220
rect -590 -89255 -500 -89220
rect -1500 -89260 -500 -89255
rect -375 -89885 -320 -88420
rect -280 -89220 -130 -89215
rect -280 -89255 -270 -89220
rect -280 -89260 -130 -89255
rect -375 -89920 -370 -89885
rect -325 -89920 -320 -89885
rect -1500 -90720 -500 -90715
rect -1500 -90755 -790 -90720
rect -590 -90755 -500 -90720
rect -1500 -90760 -500 -90755
rect -375 -91385 -320 -89920
rect -280 -90720 -130 -90715
rect -280 -90755 -270 -90720
rect -280 -90760 -130 -90755
rect -375 -91420 -370 -91385
rect -325 -91420 -320 -91385
rect -1500 -92220 -500 -92215
rect -1500 -92255 -790 -92220
rect -590 -92255 -500 -92220
rect -1500 -92260 -500 -92255
rect -375 -92885 -320 -91420
rect -280 -92220 -130 -92215
rect -280 -92255 -270 -92220
rect -280 -92260 -130 -92255
rect -375 -92920 -370 -92885
rect -325 -92920 -320 -92885
rect -1500 -93720 -500 -93715
rect -1500 -93755 -790 -93720
rect -590 -93755 -500 -93720
rect -1500 -93760 -500 -93755
rect -375 -94385 -320 -92920
rect -280 -93720 -130 -93715
rect -280 -93755 -270 -93720
rect -280 -93760 -130 -93755
rect -375 -94420 -370 -94385
rect -325 -94420 -320 -94385
rect -1500 -95220 -500 -95215
rect -1500 -95255 -790 -95220
rect -590 -95255 -500 -95220
rect -1500 -95260 -500 -95255
rect -375 -95885 -320 -94420
rect -280 -95220 -130 -95215
rect -280 -95255 -270 -95220
rect -280 -95260 -130 -95255
rect -375 -95920 -370 -95885
rect -325 -95920 -320 -95885
rect -1500 -96720 -500 -96715
rect -1500 -96755 -790 -96720
rect -590 -96755 -500 -96720
rect -1500 -96760 -500 -96755
rect -375 -97385 -320 -95920
rect -280 -96720 -130 -96715
rect -280 -96755 -270 -96720
rect -280 -96760 -130 -96755
rect -375 -97420 -370 -97385
rect -325 -97420 -320 -97385
rect -1500 -98220 -500 -98215
rect -1500 -98255 -790 -98220
rect -590 -98255 -500 -98220
rect -1500 -98260 -500 -98255
rect -375 -98885 -320 -97420
rect -280 -98220 -130 -98215
rect -280 -98255 -270 -98220
rect -280 -98260 -130 -98255
rect -375 -98920 -370 -98885
rect -325 -98920 -320 -98885
rect -1500 -99720 -500 -99715
rect -1500 -99755 -790 -99720
rect -590 -99755 -500 -99720
rect -1500 -99760 -500 -99755
rect -375 -100385 -320 -98920
rect -280 -99720 -130 -99715
rect -280 -99755 -270 -99720
rect -280 -99760 -130 -99755
rect -375 -100420 -370 -100385
rect -325 -100420 -320 -100385
rect -1500 -101220 -500 -101215
rect -1500 -101255 -790 -101220
rect -590 -101255 -500 -101220
rect -1500 -101260 -500 -101255
rect -375 -101885 -320 -100420
rect -280 -101220 -130 -101215
rect -280 -101255 -270 -101220
rect -280 -101260 -130 -101255
rect -375 -101920 -370 -101885
rect -325 -101920 -320 -101885
rect -1500 -102720 -500 -102715
rect -1500 -102755 -790 -102720
rect -590 -102755 -500 -102720
rect -1500 -102760 -500 -102755
rect -375 -103385 -320 -101920
rect -280 -102720 -130 -102715
rect -280 -102755 -270 -102720
rect -280 -102760 -130 -102755
rect -375 -103420 -370 -103385
rect -325 -103420 -320 -103385
rect -1500 -104220 -500 -104215
rect -1500 -104255 -790 -104220
rect -590 -104255 -500 -104220
rect -1500 -104260 -500 -104255
rect -375 -104885 -320 -103420
rect -280 -104220 -130 -104215
rect -280 -104255 -270 -104220
rect -280 -104260 -130 -104255
rect -375 -104920 -370 -104885
rect -325 -104920 -320 -104885
rect -1500 -105720 -500 -105715
rect -1500 -105755 -790 -105720
rect -590 -105755 -500 -105720
rect -1500 -105760 -500 -105755
rect -375 -106385 -320 -104920
rect -280 -105720 -130 -105715
rect -280 -105755 -270 -105720
rect -280 -105760 -130 -105755
rect -375 -106420 -370 -106385
rect -325 -106420 -320 -106385
rect -1500 -107220 -500 -107215
rect -1500 -107255 -790 -107220
rect -590 -107255 -500 -107220
rect -1500 -107260 -500 -107255
rect -375 -107885 -320 -106420
rect -280 -107220 -130 -107215
rect -280 -107255 -270 -107220
rect -280 -107260 -130 -107255
rect -375 -107920 -370 -107885
rect -325 -107920 -320 -107885
rect -1500 -108720 -500 -108715
rect -1500 -108755 -790 -108720
rect -590 -108755 -500 -108720
rect -1500 -108760 -500 -108755
rect -375 -109385 -320 -107920
rect -280 -108720 -130 -108715
rect -280 -108755 -270 -108720
rect -280 -108760 -130 -108755
rect -375 -109420 -370 -109385
rect -325 -109420 -320 -109385
rect -1500 -110220 -500 -110215
rect -1500 -110255 -790 -110220
rect -590 -110255 -500 -110220
rect -1500 -110260 -500 -110255
rect -375 -110885 -320 -109420
rect -280 -110220 -130 -110215
rect -280 -110255 -270 -110220
rect -280 -110260 -130 -110255
rect -375 -110920 -370 -110885
rect -325 -110920 -320 -110885
rect -1500 -111720 -500 -111715
rect -1500 -111755 -790 -111720
rect -590 -111755 -500 -111720
rect -1500 -111760 -500 -111755
rect -375 -112385 -320 -110920
rect -280 -111720 -130 -111715
rect -280 -111755 -270 -111720
rect -280 -111760 -130 -111755
rect -375 -112420 -370 -112385
rect -325 -112420 -320 -112385
rect -1500 -113220 -500 -113215
rect -1500 -113255 -790 -113220
rect -590 -113255 -500 -113220
rect -1500 -113260 -500 -113255
rect -375 -113885 -320 -112420
rect -280 -113220 -130 -113215
rect -280 -113255 -270 -113220
rect -280 -113260 -130 -113255
rect -375 -113920 -370 -113885
rect -325 -113920 -320 -113885
rect -1500 -114720 -500 -114715
rect -1500 -114755 -790 -114720
rect -590 -114755 -500 -114720
rect -1500 -114760 -500 -114755
rect -375 -115385 -320 -113920
rect -280 -114720 -130 -114715
rect -280 -114755 -270 -114720
rect -280 -114760 -130 -114755
rect -375 -115420 -370 -115385
rect -325 -115420 -320 -115385
rect -1500 -116220 -500 -116215
rect -1500 -116255 -790 -116220
rect -590 -116255 -500 -116220
rect -1500 -116260 -500 -116255
rect -375 -116885 -320 -115420
rect -280 -116220 -130 -116215
rect -280 -116255 -270 -116220
rect -280 -116260 -130 -116255
rect -375 -116920 -370 -116885
rect -325 -116920 -320 -116885
rect -1500 -117720 -500 -117715
rect -1500 -117755 -790 -117720
rect -590 -117755 -500 -117720
rect -1500 -117760 -500 -117755
rect -375 -118385 -320 -116920
rect -280 -117720 -130 -117715
rect -280 -117755 -270 -117720
rect -280 -117760 -130 -117755
rect -375 -118420 -370 -118385
rect -325 -118420 -320 -118385
rect -1500 -119220 -500 -119215
rect -1500 -119255 -790 -119220
rect -590 -119255 -500 -119220
rect -1500 -119260 -500 -119255
rect -375 -119885 -320 -118420
rect -280 -119220 -130 -119215
rect -280 -119255 -270 -119220
rect -280 -119260 -130 -119255
rect -375 -119920 -370 -119885
rect -325 -119920 -320 -119885
rect -1500 -120720 -500 -120715
rect -1500 -120755 -790 -120720
rect -590 -120755 -500 -120720
rect -1500 -120760 -500 -120755
rect -375 -121385 -320 -119920
rect -280 -120720 -130 -120715
rect -280 -120755 -270 -120720
rect -280 -120760 -130 -120755
rect -375 -121420 -370 -121385
rect -325 -121420 -320 -121385
rect -1500 -122220 -500 -122215
rect -1500 -122255 -790 -122220
rect -590 -122255 -500 -122220
rect -1500 -122260 -500 -122255
rect -375 -122885 -320 -121420
rect -280 -122220 -130 -122215
rect -280 -122255 -270 -122220
rect -280 -122260 -130 -122255
rect -375 -122920 -370 -122885
rect -325 -122920 -320 -122885
rect -1500 -123720 -500 -123715
rect -1500 -123755 -790 -123720
rect -590 -123755 -500 -123720
rect -1500 -123760 -500 -123755
rect -375 -124385 -320 -122920
rect -280 -123720 -130 -123715
rect -280 -123755 -270 -123720
rect -280 -123760 -130 -123755
rect -375 -124420 -370 -124385
rect -325 -124420 -320 -124385
rect -1500 -125220 -500 -125215
rect -1500 -125255 -790 -125220
rect -590 -125255 -500 -125220
rect -1500 -125260 -500 -125255
rect -375 -125885 -320 -124420
rect -280 -125220 -130 -125215
rect -280 -125255 -270 -125220
rect -280 -125260 -130 -125255
rect -375 -125920 -370 -125885
rect -325 -125920 -320 -125885
rect -1500 -126720 -500 -126715
rect -1500 -126755 -790 -126720
rect -590 -126755 -500 -126720
rect -1500 -126760 -500 -126755
rect -375 -127385 -320 -125920
rect -280 -126720 -130 -126715
rect -280 -126755 -270 -126720
rect -280 -126760 -130 -126755
rect -375 -127420 -370 -127385
rect -325 -127420 -320 -127385
rect -1500 -128220 -500 -128215
rect -1500 -128255 -790 -128220
rect -590 -128255 -500 -128220
rect -1500 -128260 -500 -128255
rect -375 -128885 -320 -127420
rect -280 -128220 -130 -128215
rect -280 -128255 -270 -128220
rect -280 -128260 -130 -128255
rect -375 -128920 -370 -128885
rect -325 -128920 -320 -128885
rect -1500 -129720 -500 -129715
rect -1500 -129755 -790 -129720
rect -590 -129755 -500 -129720
rect -1500 -129760 -500 -129755
rect -375 -130385 -320 -128920
rect -280 -129720 -130 -129715
rect -280 -129755 -270 -129720
rect -280 -129760 -130 -129755
rect -375 -130420 -370 -130385
rect -325 -130420 -320 -130385
rect -1500 -131220 -500 -131215
rect -1500 -131255 -790 -131220
rect -590 -131255 -500 -131220
rect -1500 -131260 -500 -131255
rect -375 -131885 -320 -130420
rect -280 -131220 -130 -131215
rect -280 -131255 -270 -131220
rect -280 -131260 -130 -131255
rect -375 -131920 -370 -131885
rect -325 -131920 -320 -131885
rect -1500 -132720 -500 -132715
rect -1500 -132755 -790 -132720
rect -590 -132755 -500 -132720
rect -1500 -132760 -500 -132755
rect -375 -133385 -320 -131920
rect -280 -132720 -130 -132715
rect -280 -132755 -270 -132720
rect -280 -132760 -130 -132755
rect -375 -133420 -370 -133385
rect -325 -133420 -320 -133385
rect -1500 -134220 -500 -134215
rect -1500 -134255 -790 -134220
rect -590 -134255 -500 -134220
rect -1500 -134260 -500 -134255
rect -375 -134885 -320 -133420
rect -280 -134220 -130 -134215
rect -280 -134255 -270 -134220
rect -280 -134260 -130 -134255
rect -375 -134920 -370 -134885
rect -325 -134920 -320 -134885
rect -1500 -135720 -500 -135715
rect -1500 -135755 -790 -135720
rect -590 -135755 -500 -135720
rect -1500 -135760 -500 -135755
rect -375 -136385 -320 -134920
rect -280 -135720 -130 -135715
rect -280 -135755 -270 -135720
rect -280 -135760 -130 -135755
rect -375 -136420 -370 -136385
rect -325 -136420 -320 -136385
rect -1500 -137220 -500 -137215
rect -1500 -137255 -790 -137220
rect -590 -137255 -500 -137220
rect -1500 -137260 -500 -137255
rect -375 -137885 -320 -136420
rect -280 -137220 -130 -137215
rect -280 -137255 -270 -137220
rect -280 -137260 -130 -137255
rect -375 -137920 -370 -137885
rect -325 -137920 -320 -137885
rect -1500 -138720 -500 -138715
rect -1500 -138755 -790 -138720
rect -590 -138755 -500 -138720
rect -1500 -138760 -500 -138755
rect -375 -139385 -320 -137920
rect -280 -138720 -130 -138715
rect -280 -138755 -270 -138720
rect -280 -138760 -130 -138755
rect -375 -139420 -370 -139385
rect -325 -139420 -320 -139385
rect -1500 -140220 -500 -140215
rect -1500 -140255 -790 -140220
rect -590 -140255 -500 -140220
rect -1500 -140260 -500 -140255
rect -375 -140885 -320 -139420
rect -280 -140220 -130 -140215
rect -280 -140255 -270 -140220
rect -280 -140260 -130 -140255
rect -375 -140920 -370 -140885
rect -325 -140920 -320 -140885
rect -1500 -141720 -500 -141715
rect -1500 -141755 -790 -141720
rect -590 -141755 -500 -141720
rect -1500 -141760 -500 -141755
rect -375 -142385 -320 -140920
rect -280 -141720 -130 -141715
rect -280 -141755 -270 -141720
rect -280 -141760 -130 -141755
rect -375 -142420 -370 -142385
rect -325 -142420 -320 -142385
rect -1500 -143220 -500 -143215
rect -1500 -143255 -790 -143220
rect -590 -143255 -500 -143220
rect -1500 -143260 -500 -143255
rect -375 -143885 -320 -142420
rect -280 -143220 -130 -143215
rect -280 -143255 -270 -143220
rect -280 -143260 -130 -143255
rect -375 -143920 -370 -143885
rect -325 -143920 -320 -143885
rect -1500 -144720 -500 -144715
rect -1500 -144755 -790 -144720
rect -590 -144755 -500 -144720
rect -1500 -144760 -500 -144755
rect -375 -145385 -320 -143920
rect -280 -144720 -130 -144715
rect -280 -144755 -270 -144720
rect -280 -144760 -130 -144755
rect -375 -145420 -370 -145385
rect -325 -145420 -320 -145385
rect -1500 -146220 -500 -146215
rect -1500 -146255 -790 -146220
rect -590 -146255 -500 -146220
rect -1500 -146260 -500 -146255
rect -375 -146885 -320 -145420
rect -280 -146220 -130 -146215
rect -280 -146255 -270 -146220
rect -280 -146260 -130 -146255
rect -375 -146920 -370 -146885
rect -325 -146920 -320 -146885
rect -1500 -147720 -500 -147715
rect -1500 -147755 -790 -147720
rect -590 -147755 -500 -147720
rect -1500 -147760 -500 -147755
rect -375 -148385 -320 -146920
rect -280 -147720 -130 -147715
rect -280 -147755 -270 -147720
rect -280 -147760 -130 -147755
rect -375 -148420 -370 -148385
rect -325 -148420 -320 -148385
rect -375 -148500 -320 -148420
rect 270 -148540 1390 -148530
rect 270 -148600 280 -148540
rect 1380 -148590 1390 -148540
rect 1060 -148600 1390 -148590
rect 1770 -148540 2890 -148530
rect 1770 -148600 1780 -148540
rect 2880 -148590 2890 -148540
rect 2560 -148600 2890 -148590
rect 3270 -148540 4390 -148530
rect 3270 -148600 3280 -148540
rect 4380 -148590 4390 -148540
rect 4060 -148600 4390 -148590
rect 4770 -148540 5890 -148530
rect 4770 -148600 4780 -148540
rect 5880 -148590 5890 -148540
rect 5560 -148600 5890 -148590
rect 6270 -148540 7390 -148530
rect 6270 -148600 6280 -148540
rect 7380 -148590 7390 -148540
rect 7060 -148600 7390 -148590
rect 7770 -148540 8890 -148530
rect 7770 -148600 7780 -148540
rect 8880 -148590 8890 -148540
rect 8560 -148600 8890 -148590
rect 9270 -148540 10390 -148530
rect 9270 -148600 9280 -148540
rect 10380 -148590 10390 -148540
rect 10060 -148600 10390 -148590
rect 10770 -148540 11890 -148530
rect 10770 -148600 10780 -148540
rect 11880 -148590 11890 -148540
rect 11560 -148600 11890 -148590
rect 12270 -148540 13390 -148530
rect 12270 -148600 12280 -148540
rect 13380 -148590 13390 -148540
rect 13060 -148600 13390 -148590
rect 13770 -148540 14890 -148530
rect 13770 -148600 13780 -148540
rect 14880 -148590 14890 -148540
rect 14560 -148600 14890 -148590
rect 15270 -148540 16390 -148530
rect 15270 -148600 15280 -148540
rect 16380 -148590 16390 -148540
rect 16060 -148600 16390 -148590
rect 16770 -148540 17890 -148530
rect 16770 -148600 16780 -148540
rect 17880 -148590 17890 -148540
rect 17560 -148600 17890 -148590
rect 18270 -148540 19390 -148530
rect 18270 -148600 18280 -148540
rect 19380 -148590 19390 -148540
rect 19060 -148600 19390 -148590
rect 19770 -148540 20890 -148530
rect 19770 -148600 19780 -148540
rect 20880 -148590 20890 -148540
rect 20560 -148600 20890 -148590
rect 21270 -148540 22390 -148530
rect 21270 -148600 21280 -148540
rect 22380 -148590 22390 -148540
rect 22060 -148600 22390 -148590
rect 22770 -148540 23890 -148530
rect 22770 -148600 22780 -148540
rect 23880 -148590 23890 -148540
rect 23560 -148600 23890 -148590
rect 24270 -148540 25390 -148530
rect 24270 -148600 24280 -148540
rect 25380 -148590 25390 -148540
rect 25060 -148600 25390 -148590
rect 25770 -148540 26890 -148530
rect 25770 -148600 25780 -148540
rect 26880 -148590 26890 -148540
rect 26560 -148600 26890 -148590
rect 27270 -148540 28390 -148530
rect 27270 -148600 27280 -148540
rect 28380 -148590 28390 -148540
rect 28060 -148600 28390 -148590
rect 28770 -148540 29890 -148530
rect 28770 -148600 28780 -148540
rect 29880 -148590 29890 -148540
rect 29560 -148600 29890 -148590
rect 30270 -148540 31390 -148530
rect 30270 -148600 30280 -148540
rect 31380 -148590 31390 -148540
rect 31060 -148600 31390 -148590
rect 31770 -148540 32890 -148530
rect 31770 -148600 31780 -148540
rect 32880 -148590 32890 -148540
rect 32560 -148600 32890 -148590
rect 33270 -148540 34390 -148530
rect 33270 -148600 33280 -148540
rect 34380 -148590 34390 -148540
rect 34060 -148600 34390 -148590
rect 34770 -148540 35890 -148530
rect 34770 -148600 34780 -148540
rect 35880 -148590 35890 -148540
rect 35560 -148600 35890 -148590
rect 36270 -148540 37390 -148530
rect 36270 -148600 36280 -148540
rect 37380 -148590 37390 -148540
rect 37060 -148600 37390 -148590
rect 37770 -148540 38890 -148530
rect 37770 -148600 37780 -148540
rect 38880 -148590 38890 -148540
rect 38560 -148600 38890 -148590
rect 39270 -148540 40390 -148530
rect 39270 -148600 39280 -148540
rect 40380 -148590 40390 -148540
rect 40060 -148600 40390 -148590
rect 40770 -148540 41890 -148530
rect 40770 -148600 40780 -148540
rect 41880 -148590 41890 -148540
rect 41560 -148600 41890 -148590
rect 42270 -148540 43390 -148530
rect 42270 -148600 42280 -148540
rect 43380 -148590 43390 -148540
rect 43060 -148600 43390 -148590
rect 43770 -148540 44890 -148530
rect 43770 -148600 43780 -148540
rect 44880 -148590 44890 -148540
rect 44560 -148600 44890 -148590
rect 45270 -148540 46390 -148530
rect 45270 -148600 45280 -148540
rect 46380 -148590 46390 -148540
rect 46060 -148600 46390 -148590
rect 46770 -148540 47890 -148530
rect 46770 -148600 46780 -148540
rect 47880 -148590 47890 -148540
rect 47560 -148600 47890 -148590
rect 48270 -148540 49390 -148530
rect 48270 -148600 48280 -148540
rect 49380 -148590 49390 -148540
rect 49060 -148600 49390 -148590
rect 49770 -148540 50890 -148530
rect 49770 -148600 49780 -148540
rect 50880 -148590 50890 -148540
rect 50560 -148600 50890 -148590
rect 51270 -148540 52390 -148530
rect 51270 -148600 51280 -148540
rect 52380 -148590 52390 -148540
rect 52060 -148600 52390 -148590
rect 52770 -148540 53890 -148530
rect 52770 -148600 52780 -148540
rect 53880 -148590 53890 -148540
rect 53560 -148600 53890 -148590
rect 54270 -148540 55390 -148530
rect 54270 -148600 54280 -148540
rect 55380 -148590 55390 -148540
rect 55060 -148600 55390 -148590
rect 55770 -148540 56890 -148530
rect 55770 -148600 55780 -148540
rect 56880 -148590 56890 -148540
rect 56560 -148600 56890 -148590
rect 57270 -148540 58390 -148530
rect 57270 -148600 57280 -148540
rect 58380 -148590 58390 -148540
rect 58060 -148600 58390 -148590
rect 58770 -148540 59890 -148530
rect 58770 -148600 58780 -148540
rect 59880 -148590 59890 -148540
rect 59560 -148600 59890 -148590
rect 60270 -148540 61390 -148530
rect 60270 -148600 60280 -148540
rect 61380 -148590 61390 -148540
rect 61060 -148600 61390 -148590
rect 61770 -148540 62890 -148530
rect 61770 -148600 61780 -148540
rect 62880 -148590 62890 -148540
rect 62560 -148600 62890 -148590
rect 63270 -148540 64390 -148530
rect 63270 -148600 63280 -148540
rect 64380 -148590 64390 -148540
rect 64060 -148600 64390 -148590
rect 64770 -148540 65890 -148530
rect 64770 -148600 64780 -148540
rect 65880 -148590 65890 -148540
rect 65560 -148600 65890 -148590
rect 66270 -148540 67390 -148530
rect 66270 -148600 66280 -148540
rect 67380 -148590 67390 -148540
rect 67060 -148600 67390 -148590
rect 67770 -148540 68890 -148530
rect 67770 -148600 67780 -148540
rect 68880 -148590 68890 -148540
rect 68560 -148600 68890 -148590
rect 69270 -148540 70390 -148530
rect 69270 -148600 69280 -148540
rect 70380 -148590 70390 -148540
rect 70060 -148600 70390 -148590
rect 70770 -148540 71890 -148530
rect 70770 -148600 70780 -148540
rect 71880 -148590 71890 -148540
rect 71560 -148600 71890 -148590
rect 72270 -148540 73390 -148530
rect 72270 -148600 72280 -148540
rect 73380 -148590 73390 -148540
rect 73060 -148600 73390 -148590
rect 73770 -148540 74890 -148530
rect 73770 -148600 73780 -148540
rect 74880 -148590 74890 -148540
rect 74560 -148600 74890 -148590
rect 75270 -148540 76390 -148530
rect 75270 -148600 75280 -148540
rect 76380 -148590 76390 -148540
rect 76060 -148600 76390 -148590
rect 76770 -148540 77890 -148530
rect 76770 -148600 76780 -148540
rect 77880 -148590 77890 -148540
rect 77560 -148600 77890 -148590
rect 78270 -148540 79390 -148530
rect 78270 -148600 78280 -148540
rect 79380 -148590 79390 -148540
rect 79060 -148600 79390 -148590
rect 79770 -148540 80890 -148530
rect 79770 -148600 79780 -148540
rect 80880 -148590 80890 -148540
rect 80560 -148600 80890 -148590
rect 81270 -148540 82390 -148530
rect 81270 -148600 81280 -148540
rect 82380 -148590 82390 -148540
rect 82060 -148600 82390 -148590
rect 82770 -148540 83890 -148530
rect 82770 -148600 82780 -148540
rect 83880 -148590 83890 -148540
rect 83560 -148600 83890 -148590
rect 84270 -148540 85390 -148530
rect 84270 -148600 84280 -148540
rect 85380 -148590 85390 -148540
rect 85060 -148600 85390 -148590
rect 85770 -148540 86890 -148530
rect 85770 -148600 85780 -148540
rect 86880 -148590 86890 -148540
rect 86560 -148600 86890 -148590
rect 87270 -148540 88390 -148530
rect 87270 -148600 87280 -148540
rect 88380 -148590 88390 -148540
rect 88060 -148600 88390 -148590
rect 88770 -148540 89890 -148530
rect 88770 -148600 88780 -148540
rect 89880 -148590 89890 -148540
rect 89560 -148600 89890 -148590
rect 90270 -148540 91390 -148530
rect 90270 -148600 90280 -148540
rect 91380 -148590 91390 -148540
rect 91060 -148600 91390 -148590
rect 91770 -148540 92890 -148530
rect 91770 -148600 91780 -148540
rect 92880 -148590 92890 -148540
rect 92560 -148600 92890 -148590
rect 93270 -148540 94390 -148530
rect 93270 -148600 93280 -148540
rect 94380 -148590 94390 -148540
rect 94060 -148600 94390 -148590
rect 94770 -148540 95890 -148530
rect 94770 -148600 94780 -148540
rect 95880 -148590 95890 -148540
rect 95560 -148600 95890 -148590
rect 96270 -148540 97390 -148530
rect 96270 -148600 96280 -148540
rect 97380 -148590 97390 -148540
rect 97060 -148600 97390 -148590
rect 97770 -148540 98890 -148530
rect 97770 -148600 97780 -148540
rect 98880 -148590 98890 -148540
rect 98560 -148600 98890 -148590
rect 99270 -148540 100390 -148530
rect 99270 -148600 99280 -148540
rect 100380 -148590 100390 -148540
rect 100060 -148600 100390 -148590
rect 100770 -148540 101890 -148530
rect 100770 -148600 100780 -148540
rect 101880 -148590 101890 -148540
rect 101560 -148600 101890 -148590
rect 102270 -148540 103390 -148530
rect 102270 -148600 102280 -148540
rect 103380 -148590 103390 -148540
rect 103060 -148600 103390 -148590
rect 103770 -148540 104890 -148530
rect 103770 -148600 103780 -148540
rect 104880 -148590 104890 -148540
rect 104560 -148600 104890 -148590
rect 105270 -148540 106390 -148530
rect 105270 -148600 105280 -148540
rect 106380 -148590 106390 -148540
rect 106060 -148600 106390 -148590
rect 106770 -148540 107890 -148530
rect 106770 -148600 106780 -148540
rect 107880 -148590 107890 -148540
rect 107560 -148600 107890 -148590
rect 108270 -148540 109390 -148530
rect 108270 -148600 108280 -148540
rect 109380 -148590 109390 -148540
rect 109060 -148600 109390 -148590
rect 109770 -148540 110890 -148530
rect 109770 -148600 109780 -148540
rect 110880 -148590 110890 -148540
rect 110560 -148600 110890 -148590
rect 111270 -148540 112390 -148530
rect 111270 -148600 111280 -148540
rect 112380 -148590 112390 -148540
rect 112060 -148600 112390 -148590
rect 112770 -148540 113890 -148530
rect 112770 -148600 112780 -148540
rect 113880 -148590 113890 -148540
rect 113560 -148600 113890 -148590
rect 114270 -148540 115390 -148530
rect 114270 -148600 114280 -148540
rect 115380 -148590 115390 -148540
rect 115060 -148600 115390 -148590
rect 115770 -148540 116890 -148530
rect 115770 -148600 115780 -148540
rect 116880 -148590 116890 -148540
rect 116560 -148600 116890 -148590
rect 117270 -148540 118390 -148530
rect 117270 -148600 117280 -148540
rect 118380 -148590 118390 -148540
rect 118060 -148600 118390 -148590
rect 118770 -148540 119890 -148530
rect 118770 -148600 118780 -148540
rect 119880 -148590 119890 -148540
rect 119560 -148600 119890 -148590
rect 120270 -148540 121390 -148530
rect 120270 -148600 120280 -148540
rect 121380 -148590 121390 -148540
rect 121060 -148600 121390 -148590
rect 121770 -148540 122890 -148530
rect 121770 -148600 121780 -148540
rect 122880 -148590 122890 -148540
rect 122560 -148600 122890 -148590
rect 123270 -148540 124390 -148530
rect 123270 -148600 123280 -148540
rect 124380 -148590 124390 -148540
rect 124060 -148600 124390 -148590
rect 124770 -148540 125890 -148530
rect 124770 -148600 124780 -148540
rect 125880 -148590 125890 -148540
rect 125560 -148600 125890 -148590
rect 126270 -148540 127390 -148530
rect 126270 -148600 126280 -148540
rect 127380 -148590 127390 -148540
rect 127060 -148600 127390 -148590
rect 127770 -148540 128890 -148530
rect 127770 -148600 127780 -148540
rect 128880 -148590 128890 -148540
rect 128560 -148600 128890 -148590
rect 129270 -148540 130390 -148530
rect 129270 -148600 129280 -148540
rect 130380 -148590 130390 -148540
rect 130060 -148600 130390 -148590
rect 130770 -148540 131890 -148530
rect 130770 -148600 130780 -148540
rect 131880 -148590 131890 -148540
rect 131560 -148600 131890 -148590
rect 132270 -148540 133390 -148530
rect 132270 -148600 132280 -148540
rect 133380 -148590 133390 -148540
rect 133060 -148600 133390 -148590
rect 133770 -148540 134890 -148530
rect 133770 -148600 133780 -148540
rect 134880 -148590 134890 -148540
rect 134560 -148600 134890 -148590
rect 135270 -148540 136390 -148530
rect 135270 -148600 135280 -148540
rect 136380 -148590 136390 -148540
rect 136060 -148600 136390 -148590
rect 136770 -148540 137890 -148530
rect 136770 -148600 136780 -148540
rect 137880 -148590 137890 -148540
rect 137560 -148600 137890 -148590
rect 138270 -148540 139390 -148530
rect 138270 -148600 138280 -148540
rect 139380 -148590 139390 -148540
rect 139060 -148600 139390 -148590
rect 139770 -148540 140890 -148530
rect 139770 -148600 139780 -148540
rect 140880 -148590 140890 -148540
rect 140560 -148600 140890 -148590
rect 141270 -148540 142390 -148530
rect 141270 -148600 141280 -148540
rect 142380 -148590 142390 -148540
rect 142060 -148600 142390 -148590
rect 142770 -148540 143890 -148530
rect 142770 -148600 142780 -148540
rect 143880 -148590 143890 -148540
rect 143560 -148600 143890 -148590
rect 144270 -148540 145390 -148530
rect 144270 -148600 144280 -148540
rect 145380 -148590 145390 -148540
rect 145060 -148600 145390 -148590
rect 145770 -148540 146890 -148530
rect 145770 -148600 145780 -148540
rect 146880 -148590 146890 -148540
rect 146560 -148600 146890 -148590
rect 147270 -148540 148390 -148530
rect 147270 -148600 147280 -148540
rect 148380 -148590 148390 -148540
rect 148060 -148600 148390 -148590
rect 148770 -148540 149890 -148530
rect 148770 -148600 148780 -148540
rect 149880 -148590 149890 -148540
rect 149560 -148600 149890 -148590
rect 110 -148750 220 -148745
rect 110 -148850 120 -148750
rect 210 -148850 220 -148750
rect 110 -148855 220 -148850
rect 1610 -148750 1720 -148745
rect 1610 -148850 1620 -148750
rect 1710 -148850 1720 -148750
rect 1610 -148855 1720 -148850
rect 3110 -148750 3220 -148745
rect 3110 -148850 3120 -148750
rect 3210 -148850 3220 -148750
rect 3110 -148855 3220 -148850
rect 4610 -148750 4720 -148745
rect 4610 -148850 4620 -148750
rect 4710 -148850 4720 -148750
rect 4610 -148855 4720 -148850
rect 6110 -148750 6220 -148745
rect 6110 -148850 6120 -148750
rect 6210 -148850 6220 -148750
rect 6110 -148855 6220 -148850
rect 7610 -148750 7720 -148745
rect 7610 -148850 7620 -148750
rect 7710 -148850 7720 -148750
rect 7610 -148855 7720 -148850
rect 9110 -148750 9220 -148745
rect 9110 -148850 9120 -148750
rect 9210 -148850 9220 -148750
rect 9110 -148855 9220 -148850
rect 10610 -148750 10720 -148745
rect 10610 -148850 10620 -148750
rect 10710 -148850 10720 -148750
rect 10610 -148855 10720 -148850
rect 12110 -148750 12220 -148745
rect 12110 -148850 12120 -148750
rect 12210 -148850 12220 -148750
rect 12110 -148855 12220 -148850
rect 13610 -148750 13720 -148745
rect 13610 -148850 13620 -148750
rect 13710 -148850 13720 -148750
rect 13610 -148855 13720 -148850
rect 15110 -148750 15220 -148745
rect 15110 -148850 15120 -148750
rect 15210 -148850 15220 -148750
rect 15110 -148855 15220 -148850
rect 16610 -148750 16720 -148745
rect 16610 -148850 16620 -148750
rect 16710 -148850 16720 -148750
rect 16610 -148855 16720 -148850
rect 18110 -148750 18220 -148745
rect 18110 -148850 18120 -148750
rect 18210 -148850 18220 -148750
rect 18110 -148855 18220 -148850
rect 19610 -148750 19720 -148745
rect 19610 -148850 19620 -148750
rect 19710 -148850 19720 -148750
rect 19610 -148855 19720 -148850
rect 21110 -148750 21220 -148745
rect 21110 -148850 21120 -148750
rect 21210 -148850 21220 -148750
rect 21110 -148855 21220 -148850
rect 22610 -148750 22720 -148745
rect 22610 -148850 22620 -148750
rect 22710 -148850 22720 -148750
rect 22610 -148855 22720 -148850
rect 24110 -148750 24220 -148745
rect 24110 -148850 24120 -148750
rect 24210 -148850 24220 -148750
rect 24110 -148855 24220 -148850
rect 25610 -148750 25720 -148745
rect 25610 -148850 25620 -148750
rect 25710 -148850 25720 -148750
rect 25610 -148855 25720 -148850
rect 27110 -148750 27220 -148745
rect 27110 -148850 27120 -148750
rect 27210 -148850 27220 -148750
rect 27110 -148855 27220 -148850
rect 28610 -148750 28720 -148745
rect 28610 -148850 28620 -148750
rect 28710 -148850 28720 -148750
rect 28610 -148855 28720 -148850
rect 30110 -148750 30220 -148745
rect 30110 -148850 30120 -148750
rect 30210 -148850 30220 -148750
rect 30110 -148855 30220 -148850
rect 31610 -148750 31720 -148745
rect 31610 -148850 31620 -148750
rect 31710 -148850 31720 -148750
rect 31610 -148855 31720 -148850
rect 33110 -148750 33220 -148745
rect 33110 -148850 33120 -148750
rect 33210 -148850 33220 -148750
rect 33110 -148855 33220 -148850
rect 34610 -148750 34720 -148745
rect 34610 -148850 34620 -148750
rect 34710 -148850 34720 -148750
rect 34610 -148855 34720 -148850
rect 36110 -148750 36220 -148745
rect 36110 -148850 36120 -148750
rect 36210 -148850 36220 -148750
rect 36110 -148855 36220 -148850
rect 37610 -148750 37720 -148745
rect 37610 -148850 37620 -148750
rect 37710 -148850 37720 -148750
rect 37610 -148855 37720 -148850
rect 39110 -148750 39220 -148745
rect 39110 -148850 39120 -148750
rect 39210 -148850 39220 -148750
rect 39110 -148855 39220 -148850
rect 40610 -148750 40720 -148745
rect 40610 -148850 40620 -148750
rect 40710 -148850 40720 -148750
rect 40610 -148855 40720 -148850
rect 42110 -148750 42220 -148745
rect 42110 -148850 42120 -148750
rect 42210 -148850 42220 -148750
rect 42110 -148855 42220 -148850
rect 43610 -148750 43720 -148745
rect 43610 -148850 43620 -148750
rect 43710 -148850 43720 -148750
rect 43610 -148855 43720 -148850
rect 45110 -148750 45220 -148745
rect 45110 -148850 45120 -148750
rect 45210 -148850 45220 -148750
rect 45110 -148855 45220 -148850
rect 46610 -148750 46720 -148745
rect 46610 -148850 46620 -148750
rect 46710 -148850 46720 -148750
rect 46610 -148855 46720 -148850
rect 48110 -148750 48220 -148745
rect 48110 -148850 48120 -148750
rect 48210 -148850 48220 -148750
rect 48110 -148855 48220 -148850
rect 49610 -148750 49720 -148745
rect 49610 -148850 49620 -148750
rect 49710 -148850 49720 -148750
rect 49610 -148855 49720 -148850
rect 51110 -148750 51220 -148745
rect 51110 -148850 51120 -148750
rect 51210 -148850 51220 -148750
rect 51110 -148855 51220 -148850
rect 52610 -148750 52720 -148745
rect 52610 -148850 52620 -148750
rect 52710 -148850 52720 -148750
rect 52610 -148855 52720 -148850
rect 54110 -148750 54220 -148745
rect 54110 -148850 54120 -148750
rect 54210 -148850 54220 -148750
rect 54110 -148855 54220 -148850
rect 55610 -148750 55720 -148745
rect 55610 -148850 55620 -148750
rect 55710 -148850 55720 -148750
rect 55610 -148855 55720 -148850
rect 57110 -148750 57220 -148745
rect 57110 -148850 57120 -148750
rect 57210 -148850 57220 -148750
rect 57110 -148855 57220 -148850
rect 58610 -148750 58720 -148745
rect 58610 -148850 58620 -148750
rect 58710 -148850 58720 -148750
rect 58610 -148855 58720 -148850
rect 60110 -148750 60220 -148745
rect 60110 -148850 60120 -148750
rect 60210 -148850 60220 -148750
rect 60110 -148855 60220 -148850
rect 61610 -148750 61720 -148745
rect 61610 -148850 61620 -148750
rect 61710 -148850 61720 -148750
rect 61610 -148855 61720 -148850
rect 63110 -148750 63220 -148745
rect 63110 -148850 63120 -148750
rect 63210 -148850 63220 -148750
rect 63110 -148855 63220 -148850
rect 64610 -148750 64720 -148745
rect 64610 -148850 64620 -148750
rect 64710 -148850 64720 -148750
rect 64610 -148855 64720 -148850
rect 66110 -148750 66220 -148745
rect 66110 -148850 66120 -148750
rect 66210 -148850 66220 -148750
rect 66110 -148855 66220 -148850
rect 67610 -148750 67720 -148745
rect 67610 -148850 67620 -148750
rect 67710 -148850 67720 -148750
rect 67610 -148855 67720 -148850
rect 69110 -148750 69220 -148745
rect 69110 -148850 69120 -148750
rect 69210 -148850 69220 -148750
rect 69110 -148855 69220 -148850
rect 70610 -148750 70720 -148745
rect 70610 -148850 70620 -148750
rect 70710 -148850 70720 -148750
rect 70610 -148855 70720 -148850
rect 72110 -148750 72220 -148745
rect 72110 -148850 72120 -148750
rect 72210 -148850 72220 -148750
rect 72110 -148855 72220 -148850
rect 73610 -148750 73720 -148745
rect 73610 -148850 73620 -148750
rect 73710 -148850 73720 -148750
rect 73610 -148855 73720 -148850
rect 75110 -148750 75220 -148745
rect 75110 -148850 75120 -148750
rect 75210 -148850 75220 -148750
rect 75110 -148855 75220 -148850
rect 76610 -148750 76720 -148745
rect 76610 -148850 76620 -148750
rect 76710 -148850 76720 -148750
rect 76610 -148855 76720 -148850
rect 78110 -148750 78220 -148745
rect 78110 -148850 78120 -148750
rect 78210 -148850 78220 -148750
rect 78110 -148855 78220 -148850
rect 79610 -148750 79720 -148745
rect 79610 -148850 79620 -148750
rect 79710 -148850 79720 -148750
rect 79610 -148855 79720 -148850
rect 81110 -148750 81220 -148745
rect 81110 -148850 81120 -148750
rect 81210 -148850 81220 -148750
rect 81110 -148855 81220 -148850
rect 82610 -148750 82720 -148745
rect 82610 -148850 82620 -148750
rect 82710 -148850 82720 -148750
rect 82610 -148855 82720 -148850
rect 84110 -148750 84220 -148745
rect 84110 -148850 84120 -148750
rect 84210 -148850 84220 -148750
rect 84110 -148855 84220 -148850
rect 85610 -148750 85720 -148745
rect 85610 -148850 85620 -148750
rect 85710 -148850 85720 -148750
rect 85610 -148855 85720 -148850
rect 87110 -148750 87220 -148745
rect 87110 -148850 87120 -148750
rect 87210 -148850 87220 -148750
rect 87110 -148855 87220 -148850
rect 88610 -148750 88720 -148745
rect 88610 -148850 88620 -148750
rect 88710 -148850 88720 -148750
rect 88610 -148855 88720 -148850
rect 90110 -148750 90220 -148745
rect 90110 -148850 90120 -148750
rect 90210 -148850 90220 -148750
rect 90110 -148855 90220 -148850
rect 91610 -148750 91720 -148745
rect 91610 -148850 91620 -148750
rect 91710 -148850 91720 -148750
rect 91610 -148855 91720 -148850
rect 93110 -148750 93220 -148745
rect 93110 -148850 93120 -148750
rect 93210 -148850 93220 -148750
rect 93110 -148855 93220 -148850
rect 94610 -148750 94720 -148745
rect 94610 -148850 94620 -148750
rect 94710 -148850 94720 -148750
rect 94610 -148855 94720 -148850
rect 96110 -148750 96220 -148745
rect 96110 -148850 96120 -148750
rect 96210 -148850 96220 -148750
rect 96110 -148855 96220 -148850
rect 97610 -148750 97720 -148745
rect 97610 -148850 97620 -148750
rect 97710 -148850 97720 -148750
rect 97610 -148855 97720 -148850
rect 99110 -148750 99220 -148745
rect 99110 -148850 99120 -148750
rect 99210 -148850 99220 -148750
rect 99110 -148855 99220 -148850
rect 100610 -148750 100720 -148745
rect 100610 -148850 100620 -148750
rect 100710 -148850 100720 -148750
rect 100610 -148855 100720 -148850
rect 102110 -148750 102220 -148745
rect 102110 -148850 102120 -148750
rect 102210 -148850 102220 -148750
rect 102110 -148855 102220 -148850
rect 103610 -148750 103720 -148745
rect 103610 -148850 103620 -148750
rect 103710 -148850 103720 -148750
rect 103610 -148855 103720 -148850
rect 105110 -148750 105220 -148745
rect 105110 -148850 105120 -148750
rect 105210 -148850 105220 -148750
rect 105110 -148855 105220 -148850
rect 106610 -148750 106720 -148745
rect 106610 -148850 106620 -148750
rect 106710 -148850 106720 -148750
rect 106610 -148855 106720 -148850
rect 108110 -148750 108220 -148745
rect 108110 -148850 108120 -148750
rect 108210 -148850 108220 -148750
rect 108110 -148855 108220 -148850
rect 109610 -148750 109720 -148745
rect 109610 -148850 109620 -148750
rect 109710 -148850 109720 -148750
rect 109610 -148855 109720 -148850
rect 111110 -148750 111220 -148745
rect 111110 -148850 111120 -148750
rect 111210 -148850 111220 -148750
rect 111110 -148855 111220 -148850
rect 112610 -148750 112720 -148745
rect 112610 -148850 112620 -148750
rect 112710 -148850 112720 -148750
rect 112610 -148855 112720 -148850
rect 114110 -148750 114220 -148745
rect 114110 -148850 114120 -148750
rect 114210 -148850 114220 -148750
rect 114110 -148855 114220 -148850
rect 115610 -148750 115720 -148745
rect 115610 -148850 115620 -148750
rect 115710 -148850 115720 -148750
rect 115610 -148855 115720 -148850
rect 117110 -148750 117220 -148745
rect 117110 -148850 117120 -148750
rect 117210 -148850 117220 -148750
rect 117110 -148855 117220 -148850
rect 118610 -148750 118720 -148745
rect 118610 -148850 118620 -148750
rect 118710 -148850 118720 -148750
rect 118610 -148855 118720 -148850
rect 120110 -148750 120220 -148745
rect 120110 -148850 120120 -148750
rect 120210 -148850 120220 -148750
rect 120110 -148855 120220 -148850
rect 121610 -148750 121720 -148745
rect 121610 -148850 121620 -148750
rect 121710 -148850 121720 -148750
rect 121610 -148855 121720 -148850
rect 123110 -148750 123220 -148745
rect 123110 -148850 123120 -148750
rect 123210 -148850 123220 -148750
rect 123110 -148855 123220 -148850
rect 124610 -148750 124720 -148745
rect 124610 -148850 124620 -148750
rect 124710 -148850 124720 -148750
rect 124610 -148855 124720 -148850
rect 126110 -148750 126220 -148745
rect 126110 -148850 126120 -148750
rect 126210 -148850 126220 -148750
rect 126110 -148855 126220 -148850
rect 127610 -148750 127720 -148745
rect 127610 -148850 127620 -148750
rect 127710 -148850 127720 -148750
rect 127610 -148855 127720 -148850
rect 129110 -148750 129220 -148745
rect 129110 -148850 129120 -148750
rect 129210 -148850 129220 -148750
rect 129110 -148855 129220 -148850
rect 130610 -148750 130720 -148745
rect 130610 -148850 130620 -148750
rect 130710 -148850 130720 -148750
rect 130610 -148855 130720 -148850
rect 132110 -148750 132220 -148745
rect 132110 -148850 132120 -148750
rect 132210 -148850 132220 -148750
rect 132110 -148855 132220 -148850
rect 133610 -148750 133720 -148745
rect 133610 -148850 133620 -148750
rect 133710 -148850 133720 -148750
rect 133610 -148855 133720 -148850
rect 135110 -148750 135220 -148745
rect 135110 -148850 135120 -148750
rect 135210 -148850 135220 -148750
rect 135110 -148855 135220 -148850
rect 136610 -148750 136720 -148745
rect 136610 -148850 136620 -148750
rect 136710 -148850 136720 -148750
rect 136610 -148855 136720 -148850
rect 138110 -148750 138220 -148745
rect 138110 -148850 138120 -148750
rect 138210 -148850 138220 -148750
rect 138110 -148855 138220 -148850
rect 139610 -148750 139720 -148745
rect 139610 -148850 139620 -148750
rect 139710 -148850 139720 -148750
rect 139610 -148855 139720 -148850
rect 141110 -148750 141220 -148745
rect 141110 -148850 141120 -148750
rect 141210 -148850 141220 -148750
rect 141110 -148855 141220 -148850
rect 142610 -148750 142720 -148745
rect 142610 -148850 142620 -148750
rect 142710 -148850 142720 -148750
rect 142610 -148855 142720 -148850
rect 144110 -148750 144220 -148745
rect 144110 -148850 144120 -148750
rect 144210 -148850 144220 -148750
rect 144110 -148855 144220 -148850
rect 145610 -148750 145720 -148745
rect 145610 -148850 145620 -148750
rect 145710 -148850 145720 -148750
rect 145610 -148855 145720 -148850
rect 147110 -148750 147220 -148745
rect 147110 -148850 147120 -148750
rect 147210 -148850 147220 -148750
rect 147110 -148855 147220 -148850
rect 148610 -148750 148720 -148745
rect 148610 -148850 148620 -148750
rect 148710 -148850 148720 -148750
rect 148610 -148855 148720 -148850
rect 270 -148960 150370 -148950
rect 270 -149040 280 -148960
rect 270 -149050 150370 -149040
<< via2 >>
rect 245 1780 290 1825
rect 1745 1780 1790 1825
rect 3245 1780 3290 1825
rect 4745 1780 4790 1825
rect 6245 1780 6290 1825
rect 7745 1780 7790 1825
rect 9245 1780 9290 1825
rect 10745 1780 10790 1825
rect 12245 1780 12290 1825
rect 13745 1780 13790 1825
rect 15245 1780 15290 1825
rect 16745 1780 16790 1825
rect 18245 1780 18290 1825
rect 19745 1780 19790 1825
rect 21245 1780 21290 1825
rect 22745 1780 22790 1825
rect 24245 1780 24290 1825
rect 25745 1780 25790 1825
rect 27245 1780 27290 1825
rect 28745 1780 28790 1825
rect 30245 1780 30290 1825
rect 31745 1780 31790 1825
rect 33245 1780 33290 1825
rect 34745 1780 34790 1825
rect 36245 1780 36290 1825
rect 37745 1780 37790 1825
rect 39245 1780 39290 1825
rect 40745 1780 40790 1825
rect 42245 1780 42290 1825
rect 43745 1780 43790 1825
rect 45245 1780 45290 1825
rect 46745 1780 46790 1825
rect 48245 1780 48290 1825
rect 49745 1780 49790 1825
rect 51245 1780 51290 1825
rect 52745 1780 52790 1825
rect 54245 1780 54290 1825
rect 55745 1780 55790 1825
rect 57245 1780 57290 1825
rect 58745 1780 58790 1825
rect 60245 1780 60290 1825
rect 61745 1780 61790 1825
rect 63245 1780 63290 1825
rect 64745 1780 64790 1825
rect 66245 1780 66290 1825
rect 67745 1780 67790 1825
rect 69245 1780 69290 1825
rect 70745 1780 70790 1825
rect 72245 1780 72290 1825
rect 73745 1780 73790 1825
rect 75245 1780 75290 1825
rect 76745 1780 76790 1825
rect 78245 1780 78290 1825
rect 79745 1780 79790 1825
rect 81245 1780 81290 1825
rect 82745 1780 82790 1825
rect 84245 1780 84290 1825
rect 85745 1780 85790 1825
rect 87245 1780 87290 1825
rect 88745 1780 88790 1825
rect 90245 1780 90290 1825
rect 91745 1780 91790 1825
rect 93245 1780 93290 1825
rect 94745 1780 94790 1825
rect 96245 1780 96290 1825
rect 97745 1780 97790 1825
rect 99245 1780 99290 1825
rect 100745 1780 100790 1825
rect 102245 1780 102290 1825
rect 103745 1780 103790 1825
rect 105245 1780 105290 1825
rect 106745 1780 106790 1825
rect 108245 1780 108290 1825
rect 109745 1780 109790 1825
rect 111245 1780 111290 1825
rect 112745 1780 112790 1825
rect 114245 1780 114290 1825
rect 115745 1780 115790 1825
rect 117245 1780 117290 1825
rect 118745 1780 118790 1825
rect 120245 1780 120290 1825
rect 121745 1780 121790 1825
rect 123245 1780 123290 1825
rect 124745 1780 124790 1825
rect 126245 1780 126290 1825
rect 127745 1780 127790 1825
rect 129245 1780 129290 1825
rect 130745 1780 130790 1825
rect 132245 1780 132290 1825
rect 133745 1780 133790 1825
rect 135245 1780 135290 1825
rect 136745 1780 136790 1825
rect 138245 1780 138290 1825
rect 139745 1780 139790 1825
rect 141245 1780 141290 1825
rect 142745 1780 142790 1825
rect 144245 1780 144290 1825
rect 145745 1780 145790 1825
rect 147245 1780 147290 1825
rect 148745 1780 148790 1825
rect -270 745 -130 780
rect -370 80 -325 115
rect -270 -755 -130 -720
rect -370 -1420 -325 -1385
rect -270 -2255 -130 -2220
rect -370 -2920 -325 -2885
rect -270 -3755 -130 -3720
rect -370 -4420 -325 -4385
rect -270 -5255 -130 -5220
rect -370 -5920 -325 -5885
rect -270 -6755 -130 -6720
rect -370 -7420 -325 -7385
rect -270 -8255 -130 -8220
rect -370 -8920 -325 -8885
rect -270 -9755 -130 -9720
rect -370 -10420 -325 -10385
rect -270 -11255 -130 -11220
rect -370 -11920 -325 -11885
rect -270 -12755 -130 -12720
rect -370 -13420 -325 -13385
rect -270 -14255 -130 -14220
rect -370 -14920 -325 -14885
rect -270 -15755 -130 -15720
rect -370 -16420 -325 -16385
rect -270 -17255 -130 -17220
rect -370 -17920 -325 -17885
rect -270 -18755 -130 -18720
rect -370 -19420 -325 -19385
rect -270 -20255 -130 -20220
rect -370 -20920 -325 -20885
rect -270 -21755 -130 -21720
rect -370 -22420 -325 -22385
rect -270 -23255 -130 -23220
rect -370 -23920 -325 -23885
rect -270 -24755 -130 -24720
rect -370 -25420 -325 -25385
rect -270 -26255 -130 -26220
rect -370 -26920 -325 -26885
rect -270 -27755 -130 -27720
rect -370 -28420 -325 -28385
rect -270 -29255 -130 -29220
rect -370 -29920 -325 -29885
rect -270 -30755 -130 -30720
rect -370 -31420 -325 -31385
rect -270 -32255 -130 -32220
rect -370 -32920 -325 -32885
rect -270 -33755 -130 -33720
rect -370 -34420 -325 -34385
rect -270 -35255 -130 -35220
rect -370 -35920 -325 -35885
rect -270 -36755 -130 -36720
rect -370 -37420 -325 -37385
rect -270 -38255 -130 -38220
rect -370 -38920 -325 -38885
rect -270 -39755 -130 -39720
rect -370 -40420 -325 -40385
rect -270 -41255 -130 -41220
rect -370 -41920 -325 -41885
rect -270 -42755 -130 -42720
rect -370 -43420 -325 -43385
rect -270 -44255 -130 -44220
rect -370 -44920 -325 -44885
rect -270 -45755 -130 -45720
rect -370 -46420 -325 -46385
rect -270 -47255 -130 -47220
rect -370 -47920 -325 -47885
rect -270 -48755 -130 -48720
rect -370 -49420 -325 -49385
rect -270 -50255 -130 -50220
rect -370 -50920 -325 -50885
rect -270 -51755 -130 -51720
rect -370 -52420 -325 -52385
rect -270 -53255 -130 -53220
rect -370 -53920 -325 -53885
rect -270 -54755 -130 -54720
rect -370 -55420 -325 -55385
rect -270 -56255 -130 -56220
rect -370 -56920 -325 -56885
rect -270 -57755 -130 -57720
rect -370 -58420 -325 -58385
rect -270 -59255 -130 -59220
rect -370 -59920 -325 -59885
rect -270 -60755 -130 -60720
rect -370 -61420 -325 -61385
rect -270 -62255 -130 -62220
rect -370 -62920 -325 -62885
rect -270 -63755 -130 -63720
rect -370 -64420 -325 -64385
rect -270 -65255 -130 -65220
rect -370 -65920 -325 -65885
rect -270 -66755 -130 -66720
rect -370 -67420 -325 -67385
rect -270 -68255 -130 -68220
rect -370 -68920 -325 -68885
rect -270 -69755 -130 -69720
rect -370 -70420 -325 -70385
rect -270 -71255 -130 -71220
rect -370 -71920 -325 -71885
rect -270 -72755 -130 -72720
rect -370 -73420 -325 -73385
rect -270 -74255 -130 -74220
rect -370 -74920 -325 -74885
rect -270 -75755 -130 -75720
rect -370 -76420 -325 -76385
rect -270 -77255 -130 -77220
rect -370 -77920 -325 -77885
rect -270 -78755 -130 -78720
rect -370 -79420 -325 -79385
rect -270 -80255 -130 -80220
rect -370 -80920 -325 -80885
rect -270 -81755 -130 -81720
rect -370 -82420 -325 -82385
rect -270 -83255 -130 -83220
rect -370 -83920 -325 -83885
rect -270 -84755 -130 -84720
rect -370 -85420 -325 -85385
rect -270 -86255 -130 -86220
rect -370 -86920 -325 -86885
rect -270 -87755 -130 -87720
rect -370 -88420 -325 -88385
rect -270 -89255 -130 -89220
rect -370 -89920 -325 -89885
rect -270 -90755 -130 -90720
rect -370 -91420 -325 -91385
rect -270 -92255 -130 -92220
rect -370 -92920 -325 -92885
rect -270 -93755 -130 -93720
rect -370 -94420 -325 -94385
rect -270 -95255 -130 -95220
rect -370 -95920 -325 -95885
rect -270 -96755 -130 -96720
rect -370 -97420 -325 -97385
rect -270 -98255 -130 -98220
rect -370 -98920 -325 -98885
rect -270 -99755 -130 -99720
rect -370 -100420 -325 -100385
rect -270 -101255 -130 -101220
rect -370 -101920 -325 -101885
rect -270 -102755 -130 -102720
rect -370 -103420 -325 -103385
rect -270 -104255 -130 -104220
rect -370 -104920 -325 -104885
rect -270 -105755 -130 -105720
rect -370 -106420 -325 -106385
rect -270 -107255 -130 -107220
rect -370 -107920 -325 -107885
rect -270 -108755 -130 -108720
rect -370 -109420 -325 -109385
rect -270 -110255 -130 -110220
rect -370 -110920 -325 -110885
rect -270 -111755 -130 -111720
rect -370 -112420 -325 -112385
rect -270 -113255 -130 -113220
rect -370 -113920 -325 -113885
rect -270 -114755 -130 -114720
rect -370 -115420 -325 -115385
rect -270 -116255 -130 -116220
rect -370 -116920 -325 -116885
rect -270 -117755 -130 -117720
rect -370 -118420 -325 -118385
rect -270 -119255 -130 -119220
rect -370 -119920 -325 -119885
rect -270 -120755 -130 -120720
rect -370 -121420 -325 -121385
rect -270 -122255 -130 -122220
rect -370 -122920 -325 -122885
rect -270 -123755 -130 -123720
rect -370 -124420 -325 -124385
rect -270 -125255 -130 -125220
rect -370 -125920 -325 -125885
rect -270 -126755 -130 -126720
rect -370 -127420 -325 -127385
rect -270 -128255 -130 -128220
rect -370 -128920 -325 -128885
rect -270 -129755 -130 -129720
rect -370 -130420 -325 -130385
rect -270 -131255 -130 -131220
rect -370 -131920 -325 -131885
rect -270 -132755 -130 -132720
rect -370 -133420 -325 -133385
rect -270 -134255 -130 -134220
rect -370 -134920 -325 -134885
rect -270 -135755 -130 -135720
rect -370 -136420 -325 -136385
rect -270 -137255 -130 -137220
rect -370 -137920 -325 -137885
rect -270 -138755 -130 -138720
rect -370 -139420 -325 -139385
rect -270 -140255 -130 -140220
rect -370 -140920 -325 -140885
rect -270 -141755 -130 -141720
rect -370 -142420 -325 -142385
rect -270 -143255 -130 -143220
rect -370 -143920 -325 -143885
rect -270 -144755 -130 -144720
rect -370 -145420 -325 -145385
rect -270 -146255 -130 -146220
rect -370 -146920 -325 -146885
rect -270 -147755 -130 -147720
rect -370 -148420 -325 -148385
rect 280 -148565 1380 -148540
rect 280 -148590 1060 -148565
rect 1060 -148590 1380 -148565
rect 1780 -148565 2880 -148540
rect 1780 -148590 2560 -148565
rect 2560 -148590 2880 -148565
rect 3280 -148565 4380 -148540
rect 3280 -148590 4060 -148565
rect 4060 -148590 4380 -148565
rect 4780 -148565 5880 -148540
rect 4780 -148590 5560 -148565
rect 5560 -148590 5880 -148565
rect 6280 -148565 7380 -148540
rect 6280 -148590 7060 -148565
rect 7060 -148590 7380 -148565
rect 7780 -148565 8880 -148540
rect 7780 -148590 8560 -148565
rect 8560 -148590 8880 -148565
rect 9280 -148565 10380 -148540
rect 9280 -148590 10060 -148565
rect 10060 -148590 10380 -148565
rect 10780 -148565 11880 -148540
rect 10780 -148590 11560 -148565
rect 11560 -148590 11880 -148565
rect 12280 -148565 13380 -148540
rect 12280 -148590 13060 -148565
rect 13060 -148590 13380 -148565
rect 13780 -148565 14880 -148540
rect 13780 -148590 14560 -148565
rect 14560 -148590 14880 -148565
rect 15280 -148565 16380 -148540
rect 15280 -148590 16060 -148565
rect 16060 -148590 16380 -148565
rect 16780 -148565 17880 -148540
rect 16780 -148590 17560 -148565
rect 17560 -148590 17880 -148565
rect 18280 -148565 19380 -148540
rect 18280 -148590 19060 -148565
rect 19060 -148590 19380 -148565
rect 19780 -148565 20880 -148540
rect 19780 -148590 20560 -148565
rect 20560 -148590 20880 -148565
rect 21280 -148565 22380 -148540
rect 21280 -148590 22060 -148565
rect 22060 -148590 22380 -148565
rect 22780 -148565 23880 -148540
rect 22780 -148590 23560 -148565
rect 23560 -148590 23880 -148565
rect 24280 -148565 25380 -148540
rect 24280 -148590 25060 -148565
rect 25060 -148590 25380 -148565
rect 25780 -148565 26880 -148540
rect 25780 -148590 26560 -148565
rect 26560 -148590 26880 -148565
rect 27280 -148565 28380 -148540
rect 27280 -148590 28060 -148565
rect 28060 -148590 28380 -148565
rect 28780 -148565 29880 -148540
rect 28780 -148590 29560 -148565
rect 29560 -148590 29880 -148565
rect 30280 -148565 31380 -148540
rect 30280 -148590 31060 -148565
rect 31060 -148590 31380 -148565
rect 31780 -148565 32880 -148540
rect 31780 -148590 32560 -148565
rect 32560 -148590 32880 -148565
rect 33280 -148565 34380 -148540
rect 33280 -148590 34060 -148565
rect 34060 -148590 34380 -148565
rect 34780 -148565 35880 -148540
rect 34780 -148590 35560 -148565
rect 35560 -148590 35880 -148565
rect 36280 -148565 37380 -148540
rect 36280 -148590 37060 -148565
rect 37060 -148590 37380 -148565
rect 37780 -148565 38880 -148540
rect 37780 -148590 38560 -148565
rect 38560 -148590 38880 -148565
rect 39280 -148565 40380 -148540
rect 39280 -148590 40060 -148565
rect 40060 -148590 40380 -148565
rect 40780 -148565 41880 -148540
rect 40780 -148590 41560 -148565
rect 41560 -148590 41880 -148565
rect 42280 -148565 43380 -148540
rect 42280 -148590 43060 -148565
rect 43060 -148590 43380 -148565
rect 43780 -148565 44880 -148540
rect 43780 -148590 44560 -148565
rect 44560 -148590 44880 -148565
rect 45280 -148565 46380 -148540
rect 45280 -148590 46060 -148565
rect 46060 -148590 46380 -148565
rect 46780 -148565 47880 -148540
rect 46780 -148590 47560 -148565
rect 47560 -148590 47880 -148565
rect 48280 -148565 49380 -148540
rect 48280 -148590 49060 -148565
rect 49060 -148590 49380 -148565
rect 49780 -148565 50880 -148540
rect 49780 -148590 50560 -148565
rect 50560 -148590 50880 -148565
rect 51280 -148565 52380 -148540
rect 51280 -148590 52060 -148565
rect 52060 -148590 52380 -148565
rect 52780 -148565 53880 -148540
rect 52780 -148590 53560 -148565
rect 53560 -148590 53880 -148565
rect 54280 -148565 55380 -148540
rect 54280 -148590 55060 -148565
rect 55060 -148590 55380 -148565
rect 55780 -148565 56880 -148540
rect 55780 -148590 56560 -148565
rect 56560 -148590 56880 -148565
rect 57280 -148565 58380 -148540
rect 57280 -148590 58060 -148565
rect 58060 -148590 58380 -148565
rect 58780 -148565 59880 -148540
rect 58780 -148590 59560 -148565
rect 59560 -148590 59880 -148565
rect 60280 -148565 61380 -148540
rect 60280 -148590 61060 -148565
rect 61060 -148590 61380 -148565
rect 61780 -148565 62880 -148540
rect 61780 -148590 62560 -148565
rect 62560 -148590 62880 -148565
rect 63280 -148565 64380 -148540
rect 63280 -148590 64060 -148565
rect 64060 -148590 64380 -148565
rect 64780 -148565 65880 -148540
rect 64780 -148590 65560 -148565
rect 65560 -148590 65880 -148565
rect 66280 -148565 67380 -148540
rect 66280 -148590 67060 -148565
rect 67060 -148590 67380 -148565
rect 67780 -148565 68880 -148540
rect 67780 -148590 68560 -148565
rect 68560 -148590 68880 -148565
rect 69280 -148565 70380 -148540
rect 69280 -148590 70060 -148565
rect 70060 -148590 70380 -148565
rect 70780 -148565 71880 -148540
rect 70780 -148590 71560 -148565
rect 71560 -148590 71880 -148565
rect 72280 -148565 73380 -148540
rect 72280 -148590 73060 -148565
rect 73060 -148590 73380 -148565
rect 73780 -148565 74880 -148540
rect 73780 -148590 74560 -148565
rect 74560 -148590 74880 -148565
rect 75280 -148565 76380 -148540
rect 75280 -148590 76060 -148565
rect 76060 -148590 76380 -148565
rect 76780 -148565 77880 -148540
rect 76780 -148590 77560 -148565
rect 77560 -148590 77880 -148565
rect 78280 -148565 79380 -148540
rect 78280 -148590 79060 -148565
rect 79060 -148590 79380 -148565
rect 79780 -148565 80880 -148540
rect 79780 -148590 80560 -148565
rect 80560 -148590 80880 -148565
rect 81280 -148565 82380 -148540
rect 81280 -148590 82060 -148565
rect 82060 -148590 82380 -148565
rect 82780 -148565 83880 -148540
rect 82780 -148590 83560 -148565
rect 83560 -148590 83880 -148565
rect 84280 -148565 85380 -148540
rect 84280 -148590 85060 -148565
rect 85060 -148590 85380 -148565
rect 85780 -148565 86880 -148540
rect 85780 -148590 86560 -148565
rect 86560 -148590 86880 -148565
rect 87280 -148565 88380 -148540
rect 87280 -148590 88060 -148565
rect 88060 -148590 88380 -148565
rect 88780 -148565 89880 -148540
rect 88780 -148590 89560 -148565
rect 89560 -148590 89880 -148565
rect 90280 -148565 91380 -148540
rect 90280 -148590 91060 -148565
rect 91060 -148590 91380 -148565
rect 91780 -148565 92880 -148540
rect 91780 -148590 92560 -148565
rect 92560 -148590 92880 -148565
rect 93280 -148565 94380 -148540
rect 93280 -148590 94060 -148565
rect 94060 -148590 94380 -148565
rect 94780 -148565 95880 -148540
rect 94780 -148590 95560 -148565
rect 95560 -148590 95880 -148565
rect 96280 -148565 97380 -148540
rect 96280 -148590 97060 -148565
rect 97060 -148590 97380 -148565
rect 97780 -148565 98880 -148540
rect 97780 -148590 98560 -148565
rect 98560 -148590 98880 -148565
rect 99280 -148565 100380 -148540
rect 99280 -148590 100060 -148565
rect 100060 -148590 100380 -148565
rect 100780 -148565 101880 -148540
rect 100780 -148590 101560 -148565
rect 101560 -148590 101880 -148565
rect 102280 -148565 103380 -148540
rect 102280 -148590 103060 -148565
rect 103060 -148590 103380 -148565
rect 103780 -148565 104880 -148540
rect 103780 -148590 104560 -148565
rect 104560 -148590 104880 -148565
rect 105280 -148565 106380 -148540
rect 105280 -148590 106060 -148565
rect 106060 -148590 106380 -148565
rect 106780 -148565 107880 -148540
rect 106780 -148590 107560 -148565
rect 107560 -148590 107880 -148565
rect 108280 -148565 109380 -148540
rect 108280 -148590 109060 -148565
rect 109060 -148590 109380 -148565
rect 109780 -148565 110880 -148540
rect 109780 -148590 110560 -148565
rect 110560 -148590 110880 -148565
rect 111280 -148565 112380 -148540
rect 111280 -148590 112060 -148565
rect 112060 -148590 112380 -148565
rect 112780 -148565 113880 -148540
rect 112780 -148590 113560 -148565
rect 113560 -148590 113880 -148565
rect 114280 -148565 115380 -148540
rect 114280 -148590 115060 -148565
rect 115060 -148590 115380 -148565
rect 115780 -148565 116880 -148540
rect 115780 -148590 116560 -148565
rect 116560 -148590 116880 -148565
rect 117280 -148565 118380 -148540
rect 117280 -148590 118060 -148565
rect 118060 -148590 118380 -148565
rect 118780 -148565 119880 -148540
rect 118780 -148590 119560 -148565
rect 119560 -148590 119880 -148565
rect 120280 -148565 121380 -148540
rect 120280 -148590 121060 -148565
rect 121060 -148590 121380 -148565
rect 121780 -148565 122880 -148540
rect 121780 -148590 122560 -148565
rect 122560 -148590 122880 -148565
rect 123280 -148565 124380 -148540
rect 123280 -148590 124060 -148565
rect 124060 -148590 124380 -148565
rect 124780 -148565 125880 -148540
rect 124780 -148590 125560 -148565
rect 125560 -148590 125880 -148565
rect 126280 -148565 127380 -148540
rect 126280 -148590 127060 -148565
rect 127060 -148590 127380 -148565
rect 127780 -148565 128880 -148540
rect 127780 -148590 128560 -148565
rect 128560 -148590 128880 -148565
rect 129280 -148565 130380 -148540
rect 129280 -148590 130060 -148565
rect 130060 -148590 130380 -148565
rect 130780 -148565 131880 -148540
rect 130780 -148590 131560 -148565
rect 131560 -148590 131880 -148565
rect 132280 -148565 133380 -148540
rect 132280 -148590 133060 -148565
rect 133060 -148590 133380 -148565
rect 133780 -148565 134880 -148540
rect 133780 -148590 134560 -148565
rect 134560 -148590 134880 -148565
rect 135280 -148565 136380 -148540
rect 135280 -148590 136060 -148565
rect 136060 -148590 136380 -148565
rect 136780 -148565 137880 -148540
rect 136780 -148590 137560 -148565
rect 137560 -148590 137880 -148565
rect 138280 -148565 139380 -148540
rect 138280 -148590 139060 -148565
rect 139060 -148590 139380 -148565
rect 139780 -148565 140880 -148540
rect 139780 -148590 140560 -148565
rect 140560 -148590 140880 -148565
rect 141280 -148565 142380 -148540
rect 141280 -148590 142060 -148565
rect 142060 -148590 142380 -148565
rect 142780 -148565 143880 -148540
rect 142780 -148590 143560 -148565
rect 143560 -148590 143880 -148565
rect 144280 -148565 145380 -148540
rect 144280 -148590 145060 -148565
rect 145060 -148590 145380 -148565
rect 145780 -148565 146880 -148540
rect 145780 -148590 146560 -148565
rect 146560 -148590 146880 -148565
rect 147280 -148565 148380 -148540
rect 147280 -148590 148060 -148565
rect 148060 -148590 148380 -148565
rect 148780 -148565 149880 -148540
rect 148780 -148590 149560 -148565
rect 149560 -148590 149880 -148565
rect 120 -148850 210 -148750
rect 1620 -148850 1710 -148750
rect 3120 -148850 3210 -148750
rect 4620 -148850 4710 -148750
rect 6120 -148850 6210 -148750
rect 7620 -148850 7710 -148750
rect 9120 -148850 9210 -148750
rect 10620 -148850 10710 -148750
rect 12120 -148850 12210 -148750
rect 13620 -148850 13710 -148750
rect 15120 -148850 15210 -148750
rect 16620 -148850 16710 -148750
rect 18120 -148850 18210 -148750
rect 19620 -148850 19710 -148750
rect 21120 -148850 21210 -148750
rect 22620 -148850 22710 -148750
rect 24120 -148850 24210 -148750
rect 25620 -148850 25710 -148750
rect 27120 -148850 27210 -148750
rect 28620 -148850 28710 -148750
rect 30120 -148850 30210 -148750
rect 31620 -148850 31710 -148750
rect 33120 -148850 33210 -148750
rect 34620 -148850 34710 -148750
rect 36120 -148850 36210 -148750
rect 37620 -148850 37710 -148750
rect 39120 -148850 39210 -148750
rect 40620 -148850 40710 -148750
rect 42120 -148850 42210 -148750
rect 43620 -148850 43710 -148750
rect 45120 -148850 45210 -148750
rect 46620 -148850 46710 -148750
rect 48120 -148850 48210 -148750
rect 49620 -148850 49710 -148750
rect 51120 -148850 51210 -148750
rect 52620 -148850 52710 -148750
rect 54120 -148850 54210 -148750
rect 55620 -148850 55710 -148750
rect 57120 -148850 57210 -148750
rect 58620 -148850 58710 -148750
rect 60120 -148850 60210 -148750
rect 61620 -148850 61710 -148750
rect 63120 -148850 63210 -148750
rect 64620 -148850 64710 -148750
rect 66120 -148850 66210 -148750
rect 67620 -148850 67710 -148750
rect 69120 -148850 69210 -148750
rect 70620 -148850 70710 -148750
rect 72120 -148850 72210 -148750
rect 73620 -148850 73710 -148750
rect 75120 -148850 75210 -148750
rect 76620 -148850 76710 -148750
rect 78120 -148850 78210 -148750
rect 79620 -148850 79710 -148750
rect 81120 -148850 81210 -148750
rect 82620 -148850 82710 -148750
rect 84120 -148850 84210 -148750
rect 85620 -148850 85710 -148750
rect 87120 -148850 87210 -148750
rect 88620 -148850 88710 -148750
rect 90120 -148850 90210 -148750
rect 91620 -148850 91710 -148750
rect 93120 -148850 93210 -148750
rect 94620 -148850 94710 -148750
rect 96120 -148850 96210 -148750
rect 97620 -148850 97710 -148750
rect 99120 -148850 99210 -148750
rect 100620 -148850 100710 -148750
rect 102120 -148850 102210 -148750
rect 103620 -148850 103710 -148750
rect 105120 -148850 105210 -148750
rect 106620 -148850 106710 -148750
rect 108120 -148850 108210 -148750
rect 109620 -148850 109710 -148750
rect 111120 -148850 111210 -148750
rect 112620 -148850 112710 -148750
rect 114120 -148850 114210 -148750
rect 115620 -148850 115710 -148750
rect 117120 -148850 117210 -148750
rect 118620 -148850 118710 -148750
rect 120120 -148850 120210 -148750
rect 121620 -148850 121710 -148750
rect 123120 -148850 123210 -148750
rect 124620 -148850 124710 -148750
rect 126120 -148850 126210 -148750
rect 127620 -148850 127710 -148750
rect 129120 -148850 129210 -148750
rect 130620 -148850 130710 -148750
rect 132120 -148850 132210 -148750
rect 133620 -148850 133710 -148750
rect 135120 -148850 135210 -148750
rect 136620 -148850 136710 -148750
rect 138120 -148850 138210 -148750
rect 139620 -148850 139710 -148750
rect 141120 -148850 141210 -148750
rect 142620 -148850 142710 -148750
rect 144120 -148850 144210 -148750
rect 145620 -148850 145710 -148750
rect 147120 -148850 147210 -148750
rect 148620 -148850 148710 -148750
<< metal3 >>
rect -600 1420 -555 2500
rect 240 1825 295 1830
rect 240 1780 245 1825
rect 290 1780 295 1825
rect 240 1775 295 1780
rect 1740 1825 1795 1830
rect 1740 1780 1745 1825
rect 1790 1780 1795 1825
rect 1740 1775 1795 1780
rect 3240 1825 3295 1830
rect 3240 1780 3245 1825
rect 3290 1780 3295 1825
rect 3240 1775 3295 1780
rect 4740 1825 4795 1830
rect 4740 1780 4745 1825
rect 4790 1780 4795 1825
rect 4740 1775 4795 1780
rect 6240 1825 6295 1830
rect 6240 1780 6245 1825
rect 6290 1780 6295 1825
rect 6240 1775 6295 1780
rect 7740 1825 7795 1830
rect 7740 1780 7745 1825
rect 7790 1780 7795 1825
rect 7740 1775 7795 1780
rect 9240 1825 9295 1830
rect 9240 1780 9245 1825
rect 9290 1780 9295 1825
rect 9240 1775 9295 1780
rect 10740 1825 10795 1830
rect 10740 1780 10745 1825
rect 10790 1780 10795 1825
rect 10740 1775 10795 1780
rect 12240 1825 12295 1830
rect 12240 1780 12245 1825
rect 12290 1780 12295 1825
rect 12240 1775 12295 1780
rect 13740 1825 13795 1830
rect 13740 1780 13745 1825
rect 13790 1780 13795 1825
rect 13740 1775 13795 1780
rect 15240 1825 15295 1830
rect 15240 1780 15245 1825
rect 15290 1780 15295 1825
rect 15240 1775 15295 1780
rect 16740 1825 16795 1830
rect 16740 1780 16745 1825
rect 16790 1780 16795 1825
rect 16740 1775 16795 1780
rect 18240 1825 18295 1830
rect 18240 1780 18245 1825
rect 18290 1780 18295 1825
rect 18240 1775 18295 1780
rect 19740 1825 19795 1830
rect 19740 1780 19745 1825
rect 19790 1780 19795 1825
rect 19740 1775 19795 1780
rect 21240 1825 21295 1830
rect 21240 1780 21245 1825
rect 21290 1780 21295 1825
rect 21240 1775 21295 1780
rect 22740 1825 22795 1830
rect 22740 1780 22745 1825
rect 22790 1780 22795 1825
rect 22740 1775 22795 1780
rect 24240 1825 24295 1830
rect 24240 1780 24245 1825
rect 24290 1780 24295 1825
rect 24240 1775 24295 1780
rect 25740 1825 25795 1830
rect 25740 1780 25745 1825
rect 25790 1780 25795 1825
rect 25740 1775 25795 1780
rect 27240 1825 27295 1830
rect 27240 1780 27245 1825
rect 27290 1780 27295 1825
rect 27240 1775 27295 1780
rect 28740 1825 28795 1830
rect 28740 1780 28745 1825
rect 28790 1780 28795 1825
rect 28740 1775 28795 1780
rect 30240 1825 30295 1830
rect 30240 1780 30245 1825
rect 30290 1780 30295 1825
rect 30240 1775 30295 1780
rect 31740 1825 31795 1830
rect 31740 1780 31745 1825
rect 31790 1780 31795 1825
rect 31740 1775 31795 1780
rect 33240 1825 33295 1830
rect 33240 1780 33245 1825
rect 33290 1780 33295 1825
rect 33240 1775 33295 1780
rect 34740 1825 34795 1830
rect 34740 1780 34745 1825
rect 34790 1780 34795 1825
rect 34740 1775 34795 1780
rect 36240 1825 36295 1830
rect 36240 1780 36245 1825
rect 36290 1780 36295 1825
rect 36240 1775 36295 1780
rect 37740 1825 37795 1830
rect 37740 1780 37745 1825
rect 37790 1780 37795 1825
rect 37740 1775 37795 1780
rect 39240 1825 39295 1830
rect 39240 1780 39245 1825
rect 39290 1780 39295 1825
rect 39240 1775 39295 1780
rect 40740 1825 40795 1830
rect 40740 1780 40745 1825
rect 40790 1780 40795 1825
rect 40740 1775 40795 1780
rect 42240 1825 42295 1830
rect 42240 1780 42245 1825
rect 42290 1780 42295 1825
rect 42240 1775 42295 1780
rect 43740 1825 43795 1830
rect 43740 1780 43745 1825
rect 43790 1780 43795 1825
rect 43740 1775 43795 1780
rect 45240 1825 45295 1830
rect 45240 1780 45245 1825
rect 45290 1780 45295 1825
rect 45240 1775 45295 1780
rect 46740 1825 46795 1830
rect 46740 1780 46745 1825
rect 46790 1780 46795 1825
rect 46740 1775 46795 1780
rect 48240 1825 48295 1830
rect 48240 1780 48245 1825
rect 48290 1780 48295 1825
rect 48240 1775 48295 1780
rect 49740 1825 49795 1830
rect 49740 1780 49745 1825
rect 49790 1780 49795 1825
rect 49740 1775 49795 1780
rect 51240 1825 51295 1830
rect 51240 1780 51245 1825
rect 51290 1780 51295 1825
rect 51240 1775 51295 1780
rect 52740 1825 52795 1830
rect 52740 1780 52745 1825
rect 52790 1780 52795 1825
rect 52740 1775 52795 1780
rect 54240 1825 54295 1830
rect 54240 1780 54245 1825
rect 54290 1780 54295 1825
rect 54240 1775 54295 1780
rect 55740 1825 55795 1830
rect 55740 1780 55745 1825
rect 55790 1780 55795 1825
rect 55740 1775 55795 1780
rect 57240 1825 57295 1830
rect 57240 1780 57245 1825
rect 57290 1780 57295 1825
rect 57240 1775 57295 1780
rect 58740 1825 58795 1830
rect 58740 1780 58745 1825
rect 58790 1780 58795 1825
rect 58740 1775 58795 1780
rect 60240 1825 60295 1830
rect 60240 1780 60245 1825
rect 60290 1780 60295 1825
rect 60240 1775 60295 1780
rect 61740 1825 61795 1830
rect 61740 1780 61745 1825
rect 61790 1780 61795 1825
rect 61740 1775 61795 1780
rect 63240 1825 63295 1830
rect 63240 1780 63245 1825
rect 63290 1780 63295 1825
rect 63240 1775 63295 1780
rect 64740 1825 64795 1830
rect 64740 1780 64745 1825
rect 64790 1780 64795 1825
rect 64740 1775 64795 1780
rect 66240 1825 66295 1830
rect 66240 1780 66245 1825
rect 66290 1780 66295 1825
rect 66240 1775 66295 1780
rect 67740 1825 67795 1830
rect 67740 1780 67745 1825
rect 67790 1780 67795 1825
rect 67740 1775 67795 1780
rect 69240 1825 69295 1830
rect 69240 1780 69245 1825
rect 69290 1780 69295 1825
rect 69240 1775 69295 1780
rect 70740 1825 70795 1830
rect 70740 1780 70745 1825
rect 70790 1780 70795 1825
rect 70740 1775 70795 1780
rect 72240 1825 72295 1830
rect 72240 1780 72245 1825
rect 72290 1780 72295 1825
rect 72240 1775 72295 1780
rect 73740 1825 73795 1830
rect 73740 1780 73745 1825
rect 73790 1780 73795 1825
rect 73740 1775 73795 1780
rect 75240 1825 75295 1830
rect 75240 1780 75245 1825
rect 75290 1780 75295 1825
rect 75240 1775 75295 1780
rect 76740 1825 76795 1830
rect 76740 1780 76745 1825
rect 76790 1780 76795 1825
rect 76740 1775 76795 1780
rect 78240 1825 78295 1830
rect 78240 1780 78245 1825
rect 78290 1780 78295 1825
rect 78240 1775 78295 1780
rect 79740 1825 79795 1830
rect 79740 1780 79745 1825
rect 79790 1780 79795 1825
rect 79740 1775 79795 1780
rect 81240 1825 81295 1830
rect 81240 1780 81245 1825
rect 81290 1780 81295 1825
rect 81240 1775 81295 1780
rect 82740 1825 82795 1830
rect 82740 1780 82745 1825
rect 82790 1780 82795 1825
rect 82740 1775 82795 1780
rect 84240 1825 84295 1830
rect 84240 1780 84245 1825
rect 84290 1780 84295 1825
rect 84240 1775 84295 1780
rect 85740 1825 85795 1830
rect 85740 1780 85745 1825
rect 85790 1780 85795 1825
rect 85740 1775 85795 1780
rect 87240 1825 87295 1830
rect 87240 1780 87245 1825
rect 87290 1780 87295 1825
rect 87240 1775 87295 1780
rect 88740 1825 88795 1830
rect 88740 1780 88745 1825
rect 88790 1780 88795 1825
rect 88740 1775 88795 1780
rect 90240 1825 90295 1830
rect 90240 1780 90245 1825
rect 90290 1780 90295 1825
rect 90240 1775 90295 1780
rect 91740 1825 91795 1830
rect 91740 1780 91745 1825
rect 91790 1780 91795 1825
rect 91740 1775 91795 1780
rect 93240 1825 93295 1830
rect 93240 1780 93245 1825
rect 93290 1780 93295 1825
rect 93240 1775 93295 1780
rect 94740 1825 94795 1830
rect 94740 1780 94745 1825
rect 94790 1780 94795 1825
rect 94740 1775 94795 1780
rect 96240 1825 96295 1830
rect 96240 1780 96245 1825
rect 96290 1780 96295 1825
rect 96240 1775 96295 1780
rect 97740 1825 97795 1830
rect 97740 1780 97745 1825
rect 97790 1780 97795 1825
rect 97740 1775 97795 1780
rect 99240 1825 99295 1830
rect 99240 1780 99245 1825
rect 99290 1780 99295 1825
rect 99240 1775 99295 1780
rect 100740 1825 100795 1830
rect 100740 1780 100745 1825
rect 100790 1780 100795 1825
rect 100740 1775 100795 1780
rect 102240 1825 102295 1830
rect 102240 1780 102245 1825
rect 102290 1780 102295 1825
rect 102240 1775 102295 1780
rect 103740 1825 103795 1830
rect 103740 1780 103745 1825
rect 103790 1780 103795 1825
rect 103740 1775 103795 1780
rect 105240 1825 105295 1830
rect 105240 1780 105245 1825
rect 105290 1780 105295 1825
rect 105240 1775 105295 1780
rect 106740 1825 106795 1830
rect 106740 1780 106745 1825
rect 106790 1780 106795 1825
rect 106740 1775 106795 1780
rect 108240 1825 108295 1830
rect 108240 1780 108245 1825
rect 108290 1780 108295 1825
rect 108240 1775 108295 1780
rect 109740 1825 109795 1830
rect 109740 1780 109745 1825
rect 109790 1780 109795 1825
rect 109740 1775 109795 1780
rect 111240 1825 111295 1830
rect 111240 1780 111245 1825
rect 111290 1780 111295 1825
rect 111240 1775 111295 1780
rect 112740 1825 112795 1830
rect 112740 1780 112745 1825
rect 112790 1780 112795 1825
rect 112740 1775 112795 1780
rect 114240 1825 114295 1830
rect 114240 1780 114245 1825
rect 114290 1780 114295 1825
rect 114240 1775 114295 1780
rect 115740 1825 115795 1830
rect 115740 1780 115745 1825
rect 115790 1780 115795 1825
rect 115740 1775 115795 1780
rect 117240 1825 117295 1830
rect 117240 1780 117245 1825
rect 117290 1780 117295 1825
rect 117240 1775 117295 1780
rect 118740 1825 118795 1830
rect 118740 1780 118745 1825
rect 118790 1780 118795 1825
rect 118740 1775 118795 1780
rect 120240 1825 120295 1830
rect 120240 1780 120245 1825
rect 120290 1780 120295 1825
rect 120240 1775 120295 1780
rect 121740 1825 121795 1830
rect 121740 1780 121745 1825
rect 121790 1780 121795 1825
rect 121740 1775 121795 1780
rect 123240 1825 123295 1830
rect 123240 1780 123245 1825
rect 123290 1780 123295 1825
rect 123240 1775 123295 1780
rect 124740 1825 124795 1830
rect 124740 1780 124745 1825
rect 124790 1780 124795 1825
rect 124740 1775 124795 1780
rect 126240 1825 126295 1830
rect 126240 1780 126245 1825
rect 126290 1780 126295 1825
rect 126240 1775 126295 1780
rect 127740 1825 127795 1830
rect 127740 1780 127745 1825
rect 127790 1780 127795 1825
rect 127740 1775 127795 1780
rect 129240 1825 129295 1830
rect 129240 1780 129245 1825
rect 129290 1780 129295 1825
rect 129240 1775 129295 1780
rect 130740 1825 130795 1830
rect 130740 1780 130745 1825
rect 130790 1780 130795 1825
rect 130740 1775 130795 1780
rect 132240 1825 132295 1830
rect 132240 1780 132245 1825
rect 132290 1780 132295 1825
rect 132240 1775 132295 1780
rect 133740 1825 133795 1830
rect 133740 1780 133745 1825
rect 133790 1780 133795 1825
rect 133740 1775 133795 1780
rect 135240 1825 135295 1830
rect 135240 1780 135245 1825
rect 135290 1780 135295 1825
rect 135240 1775 135295 1780
rect 136740 1825 136795 1830
rect 136740 1780 136745 1825
rect 136790 1780 136795 1825
rect 136740 1775 136795 1780
rect 138240 1825 138295 1830
rect 138240 1780 138245 1825
rect 138290 1780 138295 1825
rect 138240 1775 138295 1780
rect 139740 1825 139795 1830
rect 139740 1780 139745 1825
rect 139790 1780 139795 1825
rect 139740 1775 139795 1780
rect 141240 1825 141295 1830
rect 141240 1780 141245 1825
rect 141290 1780 141295 1825
rect 141240 1775 141295 1780
rect 142740 1825 142795 1830
rect 142740 1780 142745 1825
rect 142790 1780 142795 1825
rect 142740 1775 142795 1780
rect 144240 1825 144295 1830
rect 144240 1780 144245 1825
rect 144290 1780 144295 1825
rect 144240 1775 144295 1780
rect 145740 1825 145795 1830
rect 145740 1780 145745 1825
rect 145790 1780 145795 1825
rect 145740 1775 145795 1780
rect 147240 1825 147295 1830
rect 147240 1780 147245 1825
rect 147290 1780 147295 1825
rect 147240 1775 147295 1780
rect 148740 1825 148795 1830
rect 148740 1780 148745 1825
rect 148790 1780 148795 1825
rect 148740 1775 148795 1780
rect -600 1375 100 1420
rect -600 -80 -555 1375
rect -240 1275 -185 1280
rect -240 1270 260 1275
rect -240 1235 -235 1270
rect -190 1235 260 1270
rect -240 1230 260 1235
rect -240 1225 -185 1230
rect -280 780 220 785
rect -280 745 -270 780
rect -130 745 220 780
rect -280 740 220 745
rect -380 115 20 125
rect -380 80 -370 115
rect -325 80 20 115
rect -375 70 -320 80
rect -600 -125 100 -80
rect -600 -1580 -555 -125
rect -240 -225 -185 -220
rect -240 -230 260 -225
rect -240 -265 -235 -230
rect -190 -265 260 -230
rect -240 -270 260 -265
rect -240 -275 -185 -270
rect -280 -720 220 -715
rect -280 -755 -270 -720
rect -130 -755 220 -720
rect -280 -760 220 -755
rect -380 -1385 20 -1375
rect -380 -1420 -370 -1385
rect -325 -1420 20 -1385
rect -375 -1430 -320 -1420
rect -600 -1625 100 -1580
rect -600 -3080 -555 -1625
rect -240 -1725 -185 -1720
rect -240 -1730 260 -1725
rect -240 -1765 -235 -1730
rect -190 -1765 260 -1730
rect -240 -1770 260 -1765
rect -240 -1775 -185 -1770
rect -280 -2220 220 -2215
rect -280 -2255 -270 -2220
rect -130 -2255 220 -2220
rect -280 -2260 220 -2255
rect -380 -2885 20 -2875
rect -380 -2920 -370 -2885
rect -325 -2920 20 -2885
rect -375 -2930 -320 -2920
rect -600 -3125 100 -3080
rect -600 -4580 -555 -3125
rect -240 -3225 -185 -3220
rect -240 -3230 260 -3225
rect -240 -3265 -235 -3230
rect -190 -3265 260 -3230
rect -240 -3270 260 -3265
rect -240 -3275 -185 -3270
rect -280 -3720 220 -3715
rect -280 -3755 -270 -3720
rect -130 -3755 220 -3720
rect -280 -3760 220 -3755
rect -380 -4385 20 -4375
rect -380 -4420 -370 -4385
rect -325 -4420 20 -4385
rect -375 -4430 -320 -4420
rect -600 -4625 100 -4580
rect -600 -6080 -555 -4625
rect -240 -4725 -185 -4720
rect -240 -4730 260 -4725
rect -240 -4765 -235 -4730
rect -190 -4765 260 -4730
rect -240 -4770 260 -4765
rect -240 -4775 -185 -4770
rect -280 -5220 220 -5215
rect -280 -5255 -270 -5220
rect -130 -5255 220 -5220
rect -280 -5260 220 -5255
rect -380 -5885 20 -5875
rect -380 -5920 -370 -5885
rect -325 -5920 20 -5885
rect -375 -5930 -320 -5920
rect -600 -6125 100 -6080
rect -600 -7580 -555 -6125
rect -240 -6225 -185 -6220
rect -240 -6230 260 -6225
rect -240 -6265 -235 -6230
rect -190 -6265 260 -6230
rect -240 -6270 260 -6265
rect -240 -6275 -185 -6270
rect -280 -6720 220 -6715
rect -280 -6755 -270 -6720
rect -130 -6755 220 -6720
rect -280 -6760 220 -6755
rect -380 -7385 20 -7375
rect -380 -7420 -370 -7385
rect -325 -7420 20 -7385
rect -375 -7430 -320 -7420
rect -600 -7625 100 -7580
rect -600 -9080 -555 -7625
rect -240 -7725 -185 -7720
rect -240 -7730 260 -7725
rect -240 -7765 -235 -7730
rect -190 -7765 260 -7730
rect -240 -7770 260 -7765
rect -240 -7775 -185 -7770
rect -280 -8220 220 -8215
rect -280 -8255 -270 -8220
rect -130 -8255 220 -8220
rect -280 -8260 220 -8255
rect -380 -8885 20 -8875
rect -380 -8920 -370 -8885
rect -325 -8920 20 -8885
rect -375 -8930 -320 -8920
rect -600 -9125 100 -9080
rect -600 -10580 -555 -9125
rect -240 -9225 -185 -9220
rect -240 -9230 260 -9225
rect -240 -9265 -235 -9230
rect -190 -9265 260 -9230
rect -240 -9270 260 -9265
rect -240 -9275 -185 -9270
rect -280 -9720 220 -9715
rect -280 -9755 -270 -9720
rect -130 -9755 220 -9720
rect -280 -9760 220 -9755
rect -380 -10385 20 -10375
rect -380 -10420 -370 -10385
rect -325 -10420 20 -10385
rect -375 -10430 -320 -10420
rect -600 -10625 100 -10580
rect -600 -12080 -555 -10625
rect -240 -10725 -185 -10720
rect -240 -10730 260 -10725
rect -240 -10765 -235 -10730
rect -190 -10765 260 -10730
rect -240 -10770 260 -10765
rect -240 -10775 -185 -10770
rect -280 -11220 220 -11215
rect -280 -11255 -270 -11220
rect -130 -11255 220 -11220
rect -280 -11260 220 -11255
rect -380 -11885 20 -11875
rect -380 -11920 -370 -11885
rect -325 -11920 20 -11885
rect -375 -11930 -320 -11920
rect -600 -12125 100 -12080
rect -600 -13580 -555 -12125
rect -240 -12225 -185 -12220
rect -240 -12230 260 -12225
rect -240 -12265 -235 -12230
rect -190 -12265 260 -12230
rect -240 -12270 260 -12265
rect -240 -12275 -185 -12270
rect -280 -12720 220 -12715
rect -280 -12755 -270 -12720
rect -130 -12755 220 -12720
rect -280 -12760 220 -12755
rect -380 -13385 20 -13375
rect -380 -13420 -370 -13385
rect -325 -13420 20 -13385
rect -375 -13430 -320 -13420
rect -600 -13625 100 -13580
rect -600 -15080 -555 -13625
rect -240 -13725 -185 -13720
rect -240 -13730 260 -13725
rect -240 -13765 -235 -13730
rect -190 -13765 260 -13730
rect -240 -13770 260 -13765
rect -240 -13775 -185 -13770
rect -280 -14220 220 -14215
rect -280 -14255 -270 -14220
rect -130 -14255 220 -14220
rect -280 -14260 220 -14255
rect -380 -14885 20 -14875
rect -380 -14920 -370 -14885
rect -325 -14920 20 -14885
rect -375 -14930 -320 -14920
rect -600 -15125 100 -15080
rect -600 -16580 -555 -15125
rect -240 -15225 -185 -15220
rect -240 -15230 260 -15225
rect -240 -15265 -235 -15230
rect -190 -15265 260 -15230
rect -240 -15270 260 -15265
rect -240 -15275 -185 -15270
rect -280 -15720 220 -15715
rect -280 -15755 -270 -15720
rect -130 -15755 220 -15720
rect -280 -15760 220 -15755
rect -380 -16385 20 -16375
rect -380 -16420 -370 -16385
rect -325 -16420 20 -16385
rect -375 -16430 -320 -16420
rect -600 -16625 100 -16580
rect -600 -18080 -555 -16625
rect -240 -16725 -185 -16720
rect -240 -16730 260 -16725
rect -240 -16765 -235 -16730
rect -190 -16765 260 -16730
rect -240 -16770 260 -16765
rect -240 -16775 -185 -16770
rect -280 -17220 220 -17215
rect -280 -17255 -270 -17220
rect -130 -17255 220 -17220
rect -280 -17260 220 -17255
rect -380 -17885 20 -17875
rect -380 -17920 -370 -17885
rect -325 -17920 20 -17885
rect -375 -17930 -320 -17920
rect -600 -18125 100 -18080
rect -600 -19580 -555 -18125
rect -240 -18225 -185 -18220
rect -240 -18230 260 -18225
rect -240 -18265 -235 -18230
rect -190 -18265 260 -18230
rect -240 -18270 260 -18265
rect -240 -18275 -185 -18270
rect -280 -18720 220 -18715
rect -280 -18755 -270 -18720
rect -130 -18755 220 -18720
rect -280 -18760 220 -18755
rect -380 -19385 20 -19375
rect -380 -19420 -370 -19385
rect -325 -19420 20 -19385
rect -375 -19430 -320 -19420
rect -600 -19625 100 -19580
rect -600 -21080 -555 -19625
rect -240 -19725 -185 -19720
rect -240 -19730 260 -19725
rect -240 -19765 -235 -19730
rect -190 -19765 260 -19730
rect -240 -19770 260 -19765
rect -240 -19775 -185 -19770
rect -280 -20220 220 -20215
rect -280 -20255 -270 -20220
rect -130 -20255 220 -20220
rect -280 -20260 220 -20255
rect -380 -20885 20 -20875
rect -380 -20920 -370 -20885
rect -325 -20920 20 -20885
rect -375 -20930 -320 -20920
rect -600 -21125 100 -21080
rect -600 -22580 -555 -21125
rect -240 -21225 -185 -21220
rect -240 -21230 260 -21225
rect -240 -21265 -235 -21230
rect -190 -21265 260 -21230
rect -240 -21270 260 -21265
rect -240 -21275 -185 -21270
rect -280 -21720 220 -21715
rect -280 -21755 -270 -21720
rect -130 -21755 220 -21720
rect -280 -21760 220 -21755
rect -380 -22385 20 -22375
rect -380 -22420 -370 -22385
rect -325 -22420 20 -22385
rect -375 -22430 -320 -22420
rect -600 -22625 100 -22580
rect -600 -24080 -555 -22625
rect -240 -22725 -185 -22720
rect -240 -22730 260 -22725
rect -240 -22765 -235 -22730
rect -190 -22765 260 -22730
rect -240 -22770 260 -22765
rect -240 -22775 -185 -22770
rect -280 -23220 220 -23215
rect -280 -23255 -270 -23220
rect -130 -23255 220 -23220
rect -280 -23260 220 -23255
rect -380 -23885 20 -23875
rect -380 -23920 -370 -23885
rect -325 -23920 20 -23885
rect -375 -23930 -320 -23920
rect -600 -24125 100 -24080
rect -600 -25580 -555 -24125
rect -240 -24225 -185 -24220
rect -240 -24230 260 -24225
rect -240 -24265 -235 -24230
rect -190 -24265 260 -24230
rect -240 -24270 260 -24265
rect -240 -24275 -185 -24270
rect -280 -24720 220 -24715
rect -280 -24755 -270 -24720
rect -130 -24755 220 -24720
rect -280 -24760 220 -24755
rect -380 -25385 20 -25375
rect -380 -25420 -370 -25385
rect -325 -25420 20 -25385
rect -375 -25430 -320 -25420
rect -600 -25625 100 -25580
rect -600 -27080 -555 -25625
rect -240 -25725 -185 -25720
rect -240 -25730 260 -25725
rect -240 -25765 -235 -25730
rect -190 -25765 260 -25730
rect -240 -25770 260 -25765
rect -240 -25775 -185 -25770
rect -280 -26220 220 -26215
rect -280 -26255 -270 -26220
rect -130 -26255 220 -26220
rect -280 -26260 220 -26255
rect -380 -26885 20 -26875
rect -380 -26920 -370 -26885
rect -325 -26920 20 -26885
rect -375 -26930 -320 -26920
rect -600 -27125 100 -27080
rect -600 -28580 -555 -27125
rect -240 -27225 -185 -27220
rect -240 -27230 260 -27225
rect -240 -27265 -235 -27230
rect -190 -27265 260 -27230
rect -240 -27270 260 -27265
rect -240 -27275 -185 -27270
rect -280 -27720 220 -27715
rect -280 -27755 -270 -27720
rect -130 -27755 220 -27720
rect -280 -27760 220 -27755
rect -380 -28385 20 -28375
rect -380 -28420 -370 -28385
rect -325 -28420 20 -28385
rect -375 -28430 -320 -28420
rect -600 -28625 100 -28580
rect -600 -30080 -555 -28625
rect -240 -28725 -185 -28720
rect -240 -28730 260 -28725
rect -240 -28765 -235 -28730
rect -190 -28765 260 -28730
rect -240 -28770 260 -28765
rect -240 -28775 -185 -28770
rect -280 -29220 220 -29215
rect -280 -29255 -270 -29220
rect -130 -29255 220 -29220
rect -280 -29260 220 -29255
rect -380 -29885 20 -29875
rect -380 -29920 -370 -29885
rect -325 -29920 20 -29885
rect -375 -29930 -320 -29920
rect -600 -30125 100 -30080
rect -600 -31580 -555 -30125
rect -240 -30225 -185 -30220
rect -240 -30230 260 -30225
rect -240 -30265 -235 -30230
rect -190 -30265 260 -30230
rect -240 -30270 260 -30265
rect -240 -30275 -185 -30270
rect -280 -30720 220 -30715
rect -280 -30755 -270 -30720
rect -130 -30755 220 -30720
rect -280 -30760 220 -30755
rect -380 -31385 20 -31375
rect -380 -31420 -370 -31385
rect -325 -31420 20 -31385
rect -375 -31430 -320 -31420
rect -600 -31625 100 -31580
rect -600 -33080 -555 -31625
rect -240 -31725 -185 -31720
rect -240 -31730 260 -31725
rect -240 -31765 -235 -31730
rect -190 -31765 260 -31730
rect -240 -31770 260 -31765
rect -240 -31775 -185 -31770
rect -280 -32220 220 -32215
rect -280 -32255 -270 -32220
rect -130 -32255 220 -32220
rect -280 -32260 220 -32255
rect -380 -32885 20 -32875
rect -380 -32920 -370 -32885
rect -325 -32920 20 -32885
rect -375 -32930 -320 -32920
rect -600 -33125 100 -33080
rect -600 -34580 -555 -33125
rect -240 -33225 -185 -33220
rect -240 -33230 260 -33225
rect -240 -33265 -235 -33230
rect -190 -33265 260 -33230
rect -240 -33270 260 -33265
rect -240 -33275 -185 -33270
rect -280 -33720 220 -33715
rect -280 -33755 -270 -33720
rect -130 -33755 220 -33720
rect -280 -33760 220 -33755
rect -380 -34385 20 -34375
rect -380 -34420 -370 -34385
rect -325 -34420 20 -34385
rect -375 -34430 -320 -34420
rect -600 -34625 100 -34580
rect -600 -36080 -555 -34625
rect -240 -34725 -185 -34720
rect -240 -34730 260 -34725
rect -240 -34765 -235 -34730
rect -190 -34765 260 -34730
rect -240 -34770 260 -34765
rect -240 -34775 -185 -34770
rect -280 -35220 220 -35215
rect -280 -35255 -270 -35220
rect -130 -35255 220 -35220
rect -280 -35260 220 -35255
rect -380 -35885 20 -35875
rect -380 -35920 -370 -35885
rect -325 -35920 20 -35885
rect -375 -35930 -320 -35920
rect -600 -36125 100 -36080
rect -600 -37580 -555 -36125
rect -240 -36225 -185 -36220
rect -240 -36230 260 -36225
rect -240 -36265 -235 -36230
rect -190 -36265 260 -36230
rect -240 -36270 260 -36265
rect -240 -36275 -185 -36270
rect -280 -36720 220 -36715
rect -280 -36755 -270 -36720
rect -130 -36755 220 -36720
rect -280 -36760 220 -36755
rect -380 -37385 20 -37375
rect -380 -37420 -370 -37385
rect -325 -37420 20 -37385
rect -375 -37430 -320 -37420
rect -600 -37625 100 -37580
rect -600 -39080 -555 -37625
rect -240 -37725 -185 -37720
rect -240 -37730 260 -37725
rect -240 -37765 -235 -37730
rect -190 -37765 260 -37730
rect -240 -37770 260 -37765
rect -240 -37775 -185 -37770
rect -280 -38220 220 -38215
rect -280 -38255 -270 -38220
rect -130 -38255 220 -38220
rect -280 -38260 220 -38255
rect -380 -38885 20 -38875
rect -380 -38920 -370 -38885
rect -325 -38920 20 -38885
rect -375 -38930 -320 -38920
rect -600 -39125 100 -39080
rect -600 -40580 -555 -39125
rect -240 -39225 -185 -39220
rect -240 -39230 260 -39225
rect -240 -39265 -235 -39230
rect -190 -39265 260 -39230
rect -240 -39270 260 -39265
rect -240 -39275 -185 -39270
rect -280 -39720 220 -39715
rect -280 -39755 -270 -39720
rect -130 -39755 220 -39720
rect -280 -39760 220 -39755
rect -380 -40385 20 -40375
rect -380 -40420 -370 -40385
rect -325 -40420 20 -40385
rect -375 -40430 -320 -40420
rect -600 -40625 100 -40580
rect -600 -42080 -555 -40625
rect -240 -40725 -185 -40720
rect -240 -40730 260 -40725
rect -240 -40765 -235 -40730
rect -190 -40765 260 -40730
rect -240 -40770 260 -40765
rect -240 -40775 -185 -40770
rect -280 -41220 220 -41215
rect -280 -41255 -270 -41220
rect -130 -41255 220 -41220
rect -280 -41260 220 -41255
rect -380 -41885 20 -41875
rect -380 -41920 -370 -41885
rect -325 -41920 20 -41885
rect -375 -41930 -320 -41920
rect -600 -42125 100 -42080
rect -600 -43580 -555 -42125
rect -240 -42225 -185 -42220
rect -240 -42230 260 -42225
rect -240 -42265 -235 -42230
rect -190 -42265 260 -42230
rect -240 -42270 260 -42265
rect -240 -42275 -185 -42270
rect -280 -42720 220 -42715
rect -280 -42755 -270 -42720
rect -130 -42755 220 -42720
rect -280 -42760 220 -42755
rect -380 -43385 20 -43375
rect -380 -43420 -370 -43385
rect -325 -43420 20 -43385
rect -375 -43430 -320 -43420
rect -600 -43625 100 -43580
rect -600 -45080 -555 -43625
rect -240 -43725 -185 -43720
rect -240 -43730 260 -43725
rect -240 -43765 -235 -43730
rect -190 -43765 260 -43730
rect -240 -43770 260 -43765
rect -240 -43775 -185 -43770
rect -280 -44220 220 -44215
rect -280 -44255 -270 -44220
rect -130 -44255 220 -44220
rect -280 -44260 220 -44255
rect -380 -44885 20 -44875
rect -380 -44920 -370 -44885
rect -325 -44920 20 -44885
rect -375 -44930 -320 -44920
rect -600 -45125 100 -45080
rect -600 -46580 -555 -45125
rect -240 -45225 -185 -45220
rect -240 -45230 260 -45225
rect -240 -45265 -235 -45230
rect -190 -45265 260 -45230
rect -240 -45270 260 -45265
rect -240 -45275 -185 -45270
rect -280 -45720 220 -45715
rect -280 -45755 -270 -45720
rect -130 -45755 220 -45720
rect -280 -45760 220 -45755
rect -380 -46385 20 -46375
rect -380 -46420 -370 -46385
rect -325 -46420 20 -46385
rect -375 -46430 -320 -46420
rect -600 -46625 100 -46580
rect -600 -48080 -555 -46625
rect -240 -46725 -185 -46720
rect -240 -46730 260 -46725
rect -240 -46765 -235 -46730
rect -190 -46765 260 -46730
rect -240 -46770 260 -46765
rect -240 -46775 -185 -46770
rect -280 -47220 220 -47215
rect -280 -47255 -270 -47220
rect -130 -47255 220 -47220
rect -280 -47260 220 -47255
rect -380 -47885 20 -47875
rect -380 -47920 -370 -47885
rect -325 -47920 20 -47885
rect -375 -47930 -320 -47920
rect -600 -48125 100 -48080
rect -600 -49580 -555 -48125
rect -240 -48225 -185 -48220
rect -240 -48230 260 -48225
rect -240 -48265 -235 -48230
rect -190 -48265 260 -48230
rect -240 -48270 260 -48265
rect -240 -48275 -185 -48270
rect -280 -48720 220 -48715
rect -280 -48755 -270 -48720
rect -130 -48755 220 -48720
rect -280 -48760 220 -48755
rect -380 -49385 20 -49375
rect -380 -49420 -370 -49385
rect -325 -49420 20 -49385
rect -375 -49430 -320 -49420
rect -600 -49625 100 -49580
rect -600 -51080 -555 -49625
rect -240 -49725 -185 -49720
rect -240 -49730 260 -49725
rect -240 -49765 -235 -49730
rect -190 -49765 260 -49730
rect -240 -49770 260 -49765
rect -240 -49775 -185 -49770
rect -280 -50220 220 -50215
rect -280 -50255 -270 -50220
rect -130 -50255 220 -50220
rect -280 -50260 220 -50255
rect -380 -50885 20 -50875
rect -380 -50920 -370 -50885
rect -325 -50920 20 -50885
rect -375 -50930 -320 -50920
rect -600 -51125 100 -51080
rect -600 -52580 -555 -51125
rect -240 -51225 -185 -51220
rect -240 -51230 260 -51225
rect -240 -51265 -235 -51230
rect -190 -51265 260 -51230
rect -240 -51270 260 -51265
rect -240 -51275 -185 -51270
rect -280 -51720 220 -51715
rect -280 -51755 -270 -51720
rect -130 -51755 220 -51720
rect -280 -51760 220 -51755
rect -380 -52385 20 -52375
rect -380 -52420 -370 -52385
rect -325 -52420 20 -52385
rect -375 -52430 -320 -52420
rect -600 -52625 100 -52580
rect -600 -54080 -555 -52625
rect -240 -52725 -185 -52720
rect -240 -52730 260 -52725
rect -240 -52765 -235 -52730
rect -190 -52765 260 -52730
rect -240 -52770 260 -52765
rect -240 -52775 -185 -52770
rect -280 -53220 220 -53215
rect -280 -53255 -270 -53220
rect -130 -53255 220 -53220
rect -280 -53260 220 -53255
rect -380 -53885 20 -53875
rect -380 -53920 -370 -53885
rect -325 -53920 20 -53885
rect -375 -53930 -320 -53920
rect -600 -54125 100 -54080
rect -600 -55580 -555 -54125
rect -240 -54225 -185 -54220
rect -240 -54230 260 -54225
rect -240 -54265 -235 -54230
rect -190 -54265 260 -54230
rect -240 -54270 260 -54265
rect -240 -54275 -185 -54270
rect -280 -54720 220 -54715
rect -280 -54755 -270 -54720
rect -130 -54755 220 -54720
rect -280 -54760 220 -54755
rect -380 -55385 20 -55375
rect -380 -55420 -370 -55385
rect -325 -55420 20 -55385
rect -375 -55430 -320 -55420
rect -600 -55625 100 -55580
rect -600 -57080 -555 -55625
rect -240 -55725 -185 -55720
rect -240 -55730 260 -55725
rect -240 -55765 -235 -55730
rect -190 -55765 260 -55730
rect -240 -55770 260 -55765
rect -240 -55775 -185 -55770
rect -280 -56220 220 -56215
rect -280 -56255 -270 -56220
rect -130 -56255 220 -56220
rect -280 -56260 220 -56255
rect -380 -56885 20 -56875
rect -380 -56920 -370 -56885
rect -325 -56920 20 -56885
rect -375 -56930 -320 -56920
rect -600 -57125 100 -57080
rect -600 -58580 -555 -57125
rect -240 -57225 -185 -57220
rect -240 -57230 260 -57225
rect -240 -57265 -235 -57230
rect -190 -57265 260 -57230
rect -240 -57270 260 -57265
rect -240 -57275 -185 -57270
rect -280 -57720 220 -57715
rect -280 -57755 -270 -57720
rect -130 -57755 220 -57720
rect -280 -57760 220 -57755
rect -380 -58385 20 -58375
rect -380 -58420 -370 -58385
rect -325 -58420 20 -58385
rect -375 -58430 -320 -58420
rect -600 -58625 100 -58580
rect -600 -60080 -555 -58625
rect -240 -58725 -185 -58720
rect -240 -58730 260 -58725
rect -240 -58765 -235 -58730
rect -190 -58765 260 -58730
rect -240 -58770 260 -58765
rect -240 -58775 -185 -58770
rect -280 -59220 220 -59215
rect -280 -59255 -270 -59220
rect -130 -59255 220 -59220
rect -280 -59260 220 -59255
rect -380 -59885 20 -59875
rect -380 -59920 -370 -59885
rect -325 -59920 20 -59885
rect -375 -59930 -320 -59920
rect -600 -60125 100 -60080
rect -600 -61580 -555 -60125
rect -240 -60225 -185 -60220
rect -240 -60230 260 -60225
rect -240 -60265 -235 -60230
rect -190 -60265 260 -60230
rect -240 -60270 260 -60265
rect -240 -60275 -185 -60270
rect -280 -60720 220 -60715
rect -280 -60755 -270 -60720
rect -130 -60755 220 -60720
rect -280 -60760 220 -60755
rect -380 -61385 20 -61375
rect -380 -61420 -370 -61385
rect -325 -61420 20 -61385
rect -375 -61430 -320 -61420
rect -600 -61625 100 -61580
rect -600 -63080 -555 -61625
rect -240 -61725 -185 -61720
rect -240 -61730 260 -61725
rect -240 -61765 -235 -61730
rect -190 -61765 260 -61730
rect -240 -61770 260 -61765
rect -240 -61775 -185 -61770
rect -280 -62220 220 -62215
rect -280 -62255 -270 -62220
rect -130 -62255 220 -62220
rect -280 -62260 220 -62255
rect -380 -62885 20 -62875
rect -380 -62920 -370 -62885
rect -325 -62920 20 -62885
rect -375 -62930 -320 -62920
rect -600 -63125 100 -63080
rect -600 -64580 -555 -63125
rect -240 -63225 -185 -63220
rect -240 -63230 260 -63225
rect -240 -63265 -235 -63230
rect -190 -63265 260 -63230
rect -240 -63270 260 -63265
rect -240 -63275 -185 -63270
rect -280 -63720 220 -63715
rect -280 -63755 -270 -63720
rect -130 -63755 220 -63720
rect -280 -63760 220 -63755
rect -380 -64385 20 -64375
rect -380 -64420 -370 -64385
rect -325 -64420 20 -64385
rect -375 -64430 -320 -64420
rect -600 -64625 100 -64580
rect -600 -66080 -555 -64625
rect -240 -64725 -185 -64720
rect -240 -64730 260 -64725
rect -240 -64765 -235 -64730
rect -190 -64765 260 -64730
rect -240 -64770 260 -64765
rect -240 -64775 -185 -64770
rect -280 -65220 220 -65215
rect -280 -65255 -270 -65220
rect -130 -65255 220 -65220
rect -280 -65260 220 -65255
rect -380 -65885 20 -65875
rect -380 -65920 -370 -65885
rect -325 -65920 20 -65885
rect -375 -65930 -320 -65920
rect -600 -66125 100 -66080
rect -600 -67580 -555 -66125
rect -240 -66225 -185 -66220
rect -240 -66230 260 -66225
rect -240 -66265 -235 -66230
rect -190 -66265 260 -66230
rect -240 -66270 260 -66265
rect -240 -66275 -185 -66270
rect -280 -66720 220 -66715
rect -280 -66755 -270 -66720
rect -130 -66755 220 -66720
rect -280 -66760 220 -66755
rect -380 -67385 20 -67375
rect -380 -67420 -370 -67385
rect -325 -67420 20 -67385
rect -375 -67430 -320 -67420
rect -600 -67625 100 -67580
rect -600 -69080 -555 -67625
rect -240 -67725 -185 -67720
rect -240 -67730 260 -67725
rect -240 -67765 -235 -67730
rect -190 -67765 260 -67730
rect -240 -67770 260 -67765
rect -240 -67775 -185 -67770
rect -280 -68220 220 -68215
rect -280 -68255 -270 -68220
rect -130 -68255 220 -68220
rect -280 -68260 220 -68255
rect -380 -68885 20 -68875
rect -380 -68920 -370 -68885
rect -325 -68920 20 -68885
rect -375 -68930 -320 -68920
rect -600 -69125 100 -69080
rect -600 -70580 -555 -69125
rect -240 -69225 -185 -69220
rect -240 -69230 260 -69225
rect -240 -69265 -235 -69230
rect -190 -69265 260 -69230
rect -240 -69270 260 -69265
rect -240 -69275 -185 -69270
rect -280 -69720 220 -69715
rect -280 -69755 -270 -69720
rect -130 -69755 220 -69720
rect -280 -69760 220 -69755
rect -380 -70385 20 -70375
rect -380 -70420 -370 -70385
rect -325 -70420 20 -70385
rect -375 -70430 -320 -70420
rect -600 -70625 100 -70580
rect -600 -72080 -555 -70625
rect -240 -70725 -185 -70720
rect -240 -70730 260 -70725
rect -240 -70765 -235 -70730
rect -190 -70765 260 -70730
rect -240 -70770 260 -70765
rect -240 -70775 -185 -70770
rect -280 -71220 220 -71215
rect -280 -71255 -270 -71220
rect -130 -71255 220 -71220
rect -280 -71260 220 -71255
rect -380 -71885 20 -71875
rect -380 -71920 -370 -71885
rect -325 -71920 20 -71885
rect -375 -71930 -320 -71920
rect -600 -72125 100 -72080
rect -600 -73580 -555 -72125
rect -240 -72225 -185 -72220
rect -240 -72230 260 -72225
rect -240 -72265 -235 -72230
rect -190 -72265 260 -72230
rect -240 -72270 260 -72265
rect -240 -72275 -185 -72270
rect -280 -72720 220 -72715
rect -280 -72755 -270 -72720
rect -130 -72755 220 -72720
rect -280 -72760 220 -72755
rect -380 -73385 20 -73375
rect -380 -73420 -370 -73385
rect -325 -73420 20 -73385
rect -375 -73430 -320 -73420
rect -600 -73625 100 -73580
rect -600 -75080 -555 -73625
rect -240 -73725 -185 -73720
rect -240 -73730 260 -73725
rect -240 -73765 -235 -73730
rect -190 -73765 260 -73730
rect -240 -73770 260 -73765
rect -240 -73775 -185 -73770
rect -280 -74220 220 -74215
rect -280 -74255 -270 -74220
rect -130 -74255 220 -74220
rect -280 -74260 220 -74255
rect -380 -74885 20 -74875
rect -380 -74920 -370 -74885
rect -325 -74920 20 -74885
rect -375 -74930 -320 -74920
rect -600 -75125 100 -75080
rect -600 -76580 -555 -75125
rect -240 -75225 -185 -75220
rect -240 -75230 260 -75225
rect -240 -75265 -235 -75230
rect -190 -75265 260 -75230
rect -240 -75270 260 -75265
rect -240 -75275 -185 -75270
rect -280 -75720 220 -75715
rect -280 -75755 -270 -75720
rect -130 -75755 220 -75720
rect -280 -75760 220 -75755
rect -380 -76385 20 -76375
rect -380 -76420 -370 -76385
rect -325 -76420 20 -76385
rect -375 -76430 -320 -76420
rect -600 -76625 100 -76580
rect -600 -78080 -555 -76625
rect -240 -76725 -185 -76720
rect -240 -76730 260 -76725
rect -240 -76765 -235 -76730
rect -190 -76765 260 -76730
rect -240 -76770 260 -76765
rect -240 -76775 -185 -76770
rect -280 -77220 220 -77215
rect -280 -77255 -270 -77220
rect -130 -77255 220 -77220
rect -280 -77260 220 -77255
rect -380 -77885 20 -77875
rect -380 -77920 -370 -77885
rect -325 -77920 20 -77885
rect -375 -77930 -320 -77920
rect -600 -78125 100 -78080
rect -600 -79580 -555 -78125
rect -240 -78225 -185 -78220
rect -240 -78230 260 -78225
rect -240 -78265 -235 -78230
rect -190 -78265 260 -78230
rect -240 -78270 260 -78265
rect -240 -78275 -185 -78270
rect -280 -78720 220 -78715
rect -280 -78755 -270 -78720
rect -130 -78755 220 -78720
rect -280 -78760 220 -78755
rect -380 -79385 20 -79375
rect -380 -79420 -370 -79385
rect -325 -79420 20 -79385
rect -375 -79430 -320 -79420
rect -600 -79625 100 -79580
rect -600 -81080 -555 -79625
rect -240 -79725 -185 -79720
rect -240 -79730 260 -79725
rect -240 -79765 -235 -79730
rect -190 -79765 260 -79730
rect -240 -79770 260 -79765
rect -240 -79775 -185 -79770
rect -280 -80220 220 -80215
rect -280 -80255 -270 -80220
rect -130 -80255 220 -80220
rect -280 -80260 220 -80255
rect -380 -80885 20 -80875
rect -380 -80920 -370 -80885
rect -325 -80920 20 -80885
rect -375 -80930 -320 -80920
rect -600 -81125 100 -81080
rect -600 -82580 -555 -81125
rect -240 -81225 -185 -81220
rect -240 -81230 260 -81225
rect -240 -81265 -235 -81230
rect -190 -81265 260 -81230
rect -240 -81270 260 -81265
rect -240 -81275 -185 -81270
rect -280 -81720 220 -81715
rect -280 -81755 -270 -81720
rect -130 -81755 220 -81720
rect -280 -81760 220 -81755
rect -380 -82385 20 -82375
rect -380 -82420 -370 -82385
rect -325 -82420 20 -82385
rect -375 -82430 -320 -82420
rect -600 -82625 100 -82580
rect -600 -84080 -555 -82625
rect -240 -82725 -185 -82720
rect -240 -82730 260 -82725
rect -240 -82765 -235 -82730
rect -190 -82765 260 -82730
rect -240 -82770 260 -82765
rect -240 -82775 -185 -82770
rect -280 -83220 220 -83215
rect -280 -83255 -270 -83220
rect -130 -83255 220 -83220
rect -280 -83260 220 -83255
rect -380 -83885 20 -83875
rect -380 -83920 -370 -83885
rect -325 -83920 20 -83885
rect -375 -83930 -320 -83920
rect -600 -84125 100 -84080
rect -600 -85580 -555 -84125
rect -240 -84225 -185 -84220
rect -240 -84230 260 -84225
rect -240 -84265 -235 -84230
rect -190 -84265 260 -84230
rect -240 -84270 260 -84265
rect -240 -84275 -185 -84270
rect -280 -84720 220 -84715
rect -280 -84755 -270 -84720
rect -130 -84755 220 -84720
rect -280 -84760 220 -84755
rect -380 -85385 20 -85375
rect -380 -85420 -370 -85385
rect -325 -85420 20 -85385
rect -375 -85430 -320 -85420
rect -600 -85625 100 -85580
rect -600 -87080 -555 -85625
rect -240 -85725 -185 -85720
rect -240 -85730 260 -85725
rect -240 -85765 -235 -85730
rect -190 -85765 260 -85730
rect -240 -85770 260 -85765
rect -240 -85775 -185 -85770
rect -280 -86220 220 -86215
rect -280 -86255 -270 -86220
rect -130 -86255 220 -86220
rect -280 -86260 220 -86255
rect -380 -86885 20 -86875
rect -380 -86920 -370 -86885
rect -325 -86920 20 -86885
rect -375 -86930 -320 -86920
rect -600 -87125 100 -87080
rect -600 -88580 -555 -87125
rect -240 -87225 -185 -87220
rect -240 -87230 260 -87225
rect -240 -87265 -235 -87230
rect -190 -87265 260 -87230
rect -240 -87270 260 -87265
rect -240 -87275 -185 -87270
rect -280 -87720 220 -87715
rect -280 -87755 -270 -87720
rect -130 -87755 220 -87720
rect -280 -87760 220 -87755
rect -380 -88385 20 -88375
rect -380 -88420 -370 -88385
rect -325 -88420 20 -88385
rect -375 -88430 -320 -88420
rect -600 -88625 100 -88580
rect -600 -90080 -555 -88625
rect -240 -88725 -185 -88720
rect -240 -88730 260 -88725
rect -240 -88765 -235 -88730
rect -190 -88765 260 -88730
rect -240 -88770 260 -88765
rect -240 -88775 -185 -88770
rect -280 -89220 220 -89215
rect -280 -89255 -270 -89220
rect -130 -89255 220 -89220
rect -280 -89260 220 -89255
rect -380 -89885 20 -89875
rect -380 -89920 -370 -89885
rect -325 -89920 20 -89885
rect -375 -89930 -320 -89920
rect -600 -90125 100 -90080
rect -600 -91580 -555 -90125
rect -240 -90225 -185 -90220
rect -240 -90230 260 -90225
rect -240 -90265 -235 -90230
rect -190 -90265 260 -90230
rect -240 -90270 260 -90265
rect -240 -90275 -185 -90270
rect -280 -90720 220 -90715
rect -280 -90755 -270 -90720
rect -130 -90755 220 -90720
rect -280 -90760 220 -90755
rect -380 -91385 20 -91375
rect -380 -91420 -370 -91385
rect -325 -91420 20 -91385
rect -375 -91430 -320 -91420
rect -600 -91625 100 -91580
rect -600 -93080 -555 -91625
rect -240 -91725 -185 -91720
rect -240 -91730 260 -91725
rect -240 -91765 -235 -91730
rect -190 -91765 260 -91730
rect -240 -91770 260 -91765
rect -240 -91775 -185 -91770
rect -280 -92220 220 -92215
rect -280 -92255 -270 -92220
rect -130 -92255 220 -92220
rect -280 -92260 220 -92255
rect -380 -92885 20 -92875
rect -380 -92920 -370 -92885
rect -325 -92920 20 -92885
rect -375 -92930 -320 -92920
rect -600 -93125 100 -93080
rect -600 -94580 -555 -93125
rect -240 -93225 -185 -93220
rect -240 -93230 260 -93225
rect -240 -93265 -235 -93230
rect -190 -93265 260 -93230
rect -240 -93270 260 -93265
rect -240 -93275 -185 -93270
rect -280 -93720 220 -93715
rect -280 -93755 -270 -93720
rect -130 -93755 220 -93720
rect -280 -93760 220 -93755
rect -380 -94385 20 -94375
rect -380 -94420 -370 -94385
rect -325 -94420 20 -94385
rect -375 -94430 -320 -94420
rect -600 -94625 100 -94580
rect -600 -96080 -555 -94625
rect -240 -94725 -185 -94720
rect -240 -94730 260 -94725
rect -240 -94765 -235 -94730
rect -190 -94765 260 -94730
rect -240 -94770 260 -94765
rect -240 -94775 -185 -94770
rect -280 -95220 220 -95215
rect -280 -95255 -270 -95220
rect -130 -95255 220 -95220
rect -280 -95260 220 -95255
rect -380 -95885 20 -95875
rect -380 -95920 -370 -95885
rect -325 -95920 20 -95885
rect -375 -95930 -320 -95920
rect -600 -96125 100 -96080
rect -600 -97580 -555 -96125
rect -240 -96225 -185 -96220
rect -240 -96230 260 -96225
rect -240 -96265 -235 -96230
rect -190 -96265 260 -96230
rect -240 -96270 260 -96265
rect -240 -96275 -185 -96270
rect -280 -96720 220 -96715
rect -280 -96755 -270 -96720
rect -130 -96755 220 -96720
rect -280 -96760 220 -96755
rect -380 -97385 20 -97375
rect -380 -97420 -370 -97385
rect -325 -97420 20 -97385
rect -375 -97430 -320 -97420
rect -600 -97625 100 -97580
rect -600 -99080 -555 -97625
rect -240 -97725 -185 -97720
rect -240 -97730 260 -97725
rect -240 -97765 -235 -97730
rect -190 -97765 260 -97730
rect -240 -97770 260 -97765
rect -240 -97775 -185 -97770
rect -280 -98220 220 -98215
rect -280 -98255 -270 -98220
rect -130 -98255 220 -98220
rect -280 -98260 220 -98255
rect -380 -98885 20 -98875
rect -380 -98920 -370 -98885
rect -325 -98920 20 -98885
rect -375 -98930 -320 -98920
rect -600 -99125 100 -99080
rect -600 -100580 -555 -99125
rect -240 -99225 -185 -99220
rect -240 -99230 260 -99225
rect -240 -99265 -235 -99230
rect -190 -99265 260 -99230
rect -240 -99270 260 -99265
rect -240 -99275 -185 -99270
rect -280 -99720 220 -99715
rect -280 -99755 -270 -99720
rect -130 -99755 220 -99720
rect -280 -99760 220 -99755
rect -380 -100385 20 -100375
rect -380 -100420 -370 -100385
rect -325 -100420 20 -100385
rect -375 -100430 -320 -100420
rect -600 -100625 100 -100580
rect -600 -102080 -555 -100625
rect -240 -100725 -185 -100720
rect -240 -100730 260 -100725
rect -240 -100765 -235 -100730
rect -190 -100765 260 -100730
rect -240 -100770 260 -100765
rect -240 -100775 -185 -100770
rect -280 -101220 220 -101215
rect -280 -101255 -270 -101220
rect -130 -101255 220 -101220
rect -280 -101260 220 -101255
rect -380 -101885 20 -101875
rect -380 -101920 -370 -101885
rect -325 -101920 20 -101885
rect -375 -101930 -320 -101920
rect -600 -102125 100 -102080
rect -600 -103580 -555 -102125
rect -240 -102225 -185 -102220
rect -240 -102230 260 -102225
rect -240 -102265 -235 -102230
rect -190 -102265 260 -102230
rect -240 -102270 260 -102265
rect -240 -102275 -185 -102270
rect -280 -102720 220 -102715
rect -280 -102755 -270 -102720
rect -130 -102755 220 -102720
rect -280 -102760 220 -102755
rect -380 -103385 20 -103375
rect -380 -103420 -370 -103385
rect -325 -103420 20 -103385
rect -375 -103430 -320 -103420
rect -600 -103625 100 -103580
rect -600 -105080 -555 -103625
rect -240 -103725 -185 -103720
rect -240 -103730 260 -103725
rect -240 -103765 -235 -103730
rect -190 -103765 260 -103730
rect -240 -103770 260 -103765
rect -240 -103775 -185 -103770
rect -280 -104220 220 -104215
rect -280 -104255 -270 -104220
rect -130 -104255 220 -104220
rect -280 -104260 220 -104255
rect -380 -104885 20 -104875
rect -380 -104920 -370 -104885
rect -325 -104920 20 -104885
rect -375 -104930 -320 -104920
rect -600 -105125 100 -105080
rect -600 -106580 -555 -105125
rect -240 -105225 -185 -105220
rect -240 -105230 260 -105225
rect -240 -105265 -235 -105230
rect -190 -105265 260 -105230
rect -240 -105270 260 -105265
rect -240 -105275 -185 -105270
rect -280 -105720 220 -105715
rect -280 -105755 -270 -105720
rect -130 -105755 220 -105720
rect -280 -105760 220 -105755
rect -380 -106385 20 -106375
rect -380 -106420 -370 -106385
rect -325 -106420 20 -106385
rect -375 -106430 -320 -106420
rect -600 -106625 100 -106580
rect -600 -108080 -555 -106625
rect -240 -106725 -185 -106720
rect -240 -106730 260 -106725
rect -240 -106765 -235 -106730
rect -190 -106765 260 -106730
rect -240 -106770 260 -106765
rect -240 -106775 -185 -106770
rect -280 -107220 220 -107215
rect -280 -107255 -270 -107220
rect -130 -107255 220 -107220
rect -280 -107260 220 -107255
rect -380 -107885 20 -107875
rect -380 -107920 -370 -107885
rect -325 -107920 20 -107885
rect -375 -107930 -320 -107920
rect -600 -108125 100 -108080
rect -600 -109580 -555 -108125
rect -240 -108225 -185 -108220
rect -240 -108230 260 -108225
rect -240 -108265 -235 -108230
rect -190 -108265 260 -108230
rect -240 -108270 260 -108265
rect -240 -108275 -185 -108270
rect -280 -108720 220 -108715
rect -280 -108755 -270 -108720
rect -130 -108755 220 -108720
rect -280 -108760 220 -108755
rect -380 -109385 20 -109375
rect -380 -109420 -370 -109385
rect -325 -109420 20 -109385
rect -375 -109430 -320 -109420
rect -600 -109625 100 -109580
rect -600 -111080 -555 -109625
rect -240 -109725 -185 -109720
rect -240 -109730 260 -109725
rect -240 -109765 -235 -109730
rect -190 -109765 260 -109730
rect -240 -109770 260 -109765
rect -240 -109775 -185 -109770
rect -280 -110220 220 -110215
rect -280 -110255 -270 -110220
rect -130 -110255 220 -110220
rect -280 -110260 220 -110255
rect -380 -110885 20 -110875
rect -380 -110920 -370 -110885
rect -325 -110920 20 -110885
rect -375 -110930 -320 -110920
rect -600 -111125 100 -111080
rect -600 -112580 -555 -111125
rect -240 -111225 -185 -111220
rect -240 -111230 260 -111225
rect -240 -111265 -235 -111230
rect -190 -111265 260 -111230
rect -240 -111270 260 -111265
rect -240 -111275 -185 -111270
rect -280 -111720 220 -111715
rect -280 -111755 -270 -111720
rect -130 -111755 220 -111720
rect -280 -111760 220 -111755
rect -380 -112385 20 -112375
rect -380 -112420 -370 -112385
rect -325 -112420 20 -112385
rect -375 -112430 -320 -112420
rect -600 -112625 100 -112580
rect -600 -114080 -555 -112625
rect -240 -112725 -185 -112720
rect -240 -112730 260 -112725
rect -240 -112765 -235 -112730
rect -190 -112765 260 -112730
rect -240 -112770 260 -112765
rect -240 -112775 -185 -112770
rect -280 -113220 220 -113215
rect -280 -113255 -270 -113220
rect -130 -113255 220 -113220
rect -280 -113260 220 -113255
rect -380 -113885 20 -113875
rect -380 -113920 -370 -113885
rect -325 -113920 20 -113885
rect -375 -113930 -320 -113920
rect -600 -114125 100 -114080
rect -600 -115580 -555 -114125
rect -240 -114225 -185 -114220
rect -240 -114230 260 -114225
rect -240 -114265 -235 -114230
rect -190 -114265 260 -114230
rect -240 -114270 260 -114265
rect -240 -114275 -185 -114270
rect -280 -114720 220 -114715
rect -280 -114755 -270 -114720
rect -130 -114755 220 -114720
rect -280 -114760 220 -114755
rect -380 -115385 20 -115375
rect -380 -115420 -370 -115385
rect -325 -115420 20 -115385
rect -375 -115430 -320 -115420
rect -600 -115625 100 -115580
rect -600 -117080 -555 -115625
rect -240 -115725 -185 -115720
rect -240 -115730 260 -115725
rect -240 -115765 -235 -115730
rect -190 -115765 260 -115730
rect -240 -115770 260 -115765
rect -240 -115775 -185 -115770
rect -280 -116220 220 -116215
rect -280 -116255 -270 -116220
rect -130 -116255 220 -116220
rect -280 -116260 220 -116255
rect -380 -116885 20 -116875
rect -380 -116920 -370 -116885
rect -325 -116920 20 -116885
rect -375 -116930 -320 -116920
rect -600 -117125 100 -117080
rect -600 -118580 -555 -117125
rect -240 -117225 -185 -117220
rect -240 -117230 260 -117225
rect -240 -117265 -235 -117230
rect -190 -117265 260 -117230
rect -240 -117270 260 -117265
rect -240 -117275 -185 -117270
rect -280 -117720 220 -117715
rect -280 -117755 -270 -117720
rect -130 -117755 220 -117720
rect -280 -117760 220 -117755
rect -380 -118385 20 -118375
rect -380 -118420 -370 -118385
rect -325 -118420 20 -118385
rect -375 -118430 -320 -118420
rect -600 -118625 100 -118580
rect -600 -120080 -555 -118625
rect -240 -118725 -185 -118720
rect -240 -118730 260 -118725
rect -240 -118765 -235 -118730
rect -190 -118765 260 -118730
rect -240 -118770 260 -118765
rect -240 -118775 -185 -118770
rect -280 -119220 220 -119215
rect -280 -119255 -270 -119220
rect -130 -119255 220 -119220
rect -280 -119260 220 -119255
rect -380 -119885 20 -119875
rect -380 -119920 -370 -119885
rect -325 -119920 20 -119885
rect -375 -119930 -320 -119920
rect -600 -120125 100 -120080
rect -600 -121580 -555 -120125
rect -240 -120225 -185 -120220
rect -240 -120230 260 -120225
rect -240 -120265 -235 -120230
rect -190 -120265 260 -120230
rect -240 -120270 260 -120265
rect -240 -120275 -185 -120270
rect -280 -120720 220 -120715
rect -280 -120755 -270 -120720
rect -130 -120755 220 -120720
rect -280 -120760 220 -120755
rect -380 -121385 20 -121375
rect -380 -121420 -370 -121385
rect -325 -121420 20 -121385
rect -375 -121430 -320 -121420
rect -600 -121625 100 -121580
rect -600 -123080 -555 -121625
rect -240 -121725 -185 -121720
rect -240 -121730 260 -121725
rect -240 -121765 -235 -121730
rect -190 -121765 260 -121730
rect -240 -121770 260 -121765
rect -240 -121775 -185 -121770
rect -280 -122220 220 -122215
rect -280 -122255 -270 -122220
rect -130 -122255 220 -122220
rect -280 -122260 220 -122255
rect -380 -122885 20 -122875
rect -380 -122920 -370 -122885
rect -325 -122920 20 -122885
rect -375 -122930 -320 -122920
rect -600 -123125 100 -123080
rect -600 -124580 -555 -123125
rect -240 -123225 -185 -123220
rect -240 -123230 260 -123225
rect -240 -123265 -235 -123230
rect -190 -123265 260 -123230
rect -240 -123270 260 -123265
rect -240 -123275 -185 -123270
rect -280 -123720 220 -123715
rect -280 -123755 -270 -123720
rect -130 -123755 220 -123720
rect -280 -123760 220 -123755
rect -380 -124385 20 -124375
rect -380 -124420 -370 -124385
rect -325 -124420 20 -124385
rect -375 -124430 -320 -124420
rect -600 -124625 100 -124580
rect -600 -126080 -555 -124625
rect -240 -124725 -185 -124720
rect -240 -124730 260 -124725
rect -240 -124765 -235 -124730
rect -190 -124765 260 -124730
rect -240 -124770 260 -124765
rect -240 -124775 -185 -124770
rect -280 -125220 220 -125215
rect -280 -125255 -270 -125220
rect -130 -125255 220 -125220
rect -280 -125260 220 -125255
rect -380 -125885 20 -125875
rect -380 -125920 -370 -125885
rect -325 -125920 20 -125885
rect -375 -125930 -320 -125920
rect -600 -126125 100 -126080
rect -600 -127580 -555 -126125
rect -240 -126225 -185 -126220
rect -240 -126230 260 -126225
rect -240 -126265 -235 -126230
rect -190 -126265 260 -126230
rect -240 -126270 260 -126265
rect -240 -126275 -185 -126270
rect -280 -126720 220 -126715
rect -280 -126755 -270 -126720
rect -130 -126755 220 -126720
rect -280 -126760 220 -126755
rect -380 -127385 20 -127375
rect -380 -127420 -370 -127385
rect -325 -127420 20 -127385
rect -375 -127430 -320 -127420
rect -600 -127625 100 -127580
rect -600 -129080 -555 -127625
rect -240 -127725 -185 -127720
rect -240 -127730 260 -127725
rect -240 -127765 -235 -127730
rect -190 -127765 260 -127730
rect -240 -127770 260 -127765
rect -240 -127775 -185 -127770
rect -280 -128220 220 -128215
rect -280 -128255 -270 -128220
rect -130 -128255 220 -128220
rect -280 -128260 220 -128255
rect -380 -128885 20 -128875
rect -380 -128920 -370 -128885
rect -325 -128920 20 -128885
rect -375 -128930 -320 -128920
rect -600 -129125 100 -129080
rect -600 -130580 -555 -129125
rect -240 -129225 -185 -129220
rect -240 -129230 260 -129225
rect -240 -129265 -235 -129230
rect -190 -129265 260 -129230
rect -240 -129270 260 -129265
rect -240 -129275 -185 -129270
rect -280 -129720 220 -129715
rect -280 -129755 -270 -129720
rect -130 -129755 220 -129720
rect -280 -129760 220 -129755
rect -380 -130385 20 -130375
rect -380 -130420 -370 -130385
rect -325 -130420 20 -130385
rect -375 -130430 -320 -130420
rect -600 -130625 100 -130580
rect -600 -132080 -555 -130625
rect -240 -130725 -185 -130720
rect -240 -130730 260 -130725
rect -240 -130765 -235 -130730
rect -190 -130765 260 -130730
rect -240 -130770 260 -130765
rect -240 -130775 -185 -130770
rect -280 -131220 220 -131215
rect -280 -131255 -270 -131220
rect -130 -131255 220 -131220
rect -280 -131260 220 -131255
rect -380 -131885 20 -131875
rect -380 -131920 -370 -131885
rect -325 -131920 20 -131885
rect -375 -131930 -320 -131920
rect -600 -132125 100 -132080
rect -600 -133580 -555 -132125
rect -240 -132225 -185 -132220
rect -240 -132230 260 -132225
rect -240 -132265 -235 -132230
rect -190 -132265 260 -132230
rect -240 -132270 260 -132265
rect -240 -132275 -185 -132270
rect -280 -132720 220 -132715
rect -280 -132755 -270 -132720
rect -130 -132755 220 -132720
rect -280 -132760 220 -132755
rect -380 -133385 20 -133375
rect -380 -133420 -370 -133385
rect -325 -133420 20 -133385
rect -375 -133430 -320 -133420
rect -600 -133625 100 -133580
rect -600 -135080 -555 -133625
rect -240 -133725 -185 -133720
rect -240 -133730 260 -133725
rect -240 -133765 -235 -133730
rect -190 -133765 260 -133730
rect -240 -133770 260 -133765
rect -240 -133775 -185 -133770
rect -280 -134220 220 -134215
rect -280 -134255 -270 -134220
rect -130 -134255 220 -134220
rect -280 -134260 220 -134255
rect -380 -134885 20 -134875
rect -380 -134920 -370 -134885
rect -325 -134920 20 -134885
rect -375 -134930 -320 -134920
rect -600 -135125 100 -135080
rect -600 -136580 -555 -135125
rect -240 -135225 -185 -135220
rect -240 -135230 260 -135225
rect -240 -135265 -235 -135230
rect -190 -135265 260 -135230
rect -240 -135270 260 -135265
rect -240 -135275 -185 -135270
rect -280 -135720 220 -135715
rect -280 -135755 -270 -135720
rect -130 -135755 220 -135720
rect -280 -135760 220 -135755
rect -380 -136385 20 -136375
rect -380 -136420 -370 -136385
rect -325 -136420 20 -136385
rect -375 -136430 -320 -136420
rect -600 -136625 100 -136580
rect -600 -138080 -555 -136625
rect -240 -136725 -185 -136720
rect -240 -136730 260 -136725
rect -240 -136765 -235 -136730
rect -190 -136765 260 -136730
rect -240 -136770 260 -136765
rect -240 -136775 -185 -136770
rect -280 -137220 220 -137215
rect -280 -137255 -270 -137220
rect -130 -137255 220 -137220
rect -280 -137260 220 -137255
rect -380 -137885 20 -137875
rect -380 -137920 -370 -137885
rect -325 -137920 20 -137885
rect -375 -137930 -320 -137920
rect -600 -138125 100 -138080
rect -600 -139580 -555 -138125
rect -240 -138225 -185 -138220
rect -240 -138230 260 -138225
rect -240 -138265 -235 -138230
rect -190 -138265 260 -138230
rect -240 -138270 260 -138265
rect -240 -138275 -185 -138270
rect -280 -138720 220 -138715
rect -280 -138755 -270 -138720
rect -130 -138755 220 -138720
rect -280 -138760 220 -138755
rect -380 -139385 20 -139375
rect -380 -139420 -370 -139385
rect -325 -139420 20 -139385
rect -375 -139430 -320 -139420
rect -600 -139625 100 -139580
rect -600 -141080 -555 -139625
rect -240 -139725 -185 -139720
rect -240 -139730 260 -139725
rect -240 -139765 -235 -139730
rect -190 -139765 260 -139730
rect -240 -139770 260 -139765
rect -240 -139775 -185 -139770
rect -280 -140220 220 -140215
rect -280 -140255 -270 -140220
rect -130 -140255 220 -140220
rect -280 -140260 220 -140255
rect -380 -140885 20 -140875
rect -380 -140920 -370 -140885
rect -325 -140920 20 -140885
rect -375 -140930 -320 -140920
rect -600 -141125 100 -141080
rect -600 -142580 -555 -141125
rect -240 -141225 -185 -141220
rect -240 -141230 260 -141225
rect -240 -141265 -235 -141230
rect -190 -141265 260 -141230
rect -240 -141270 260 -141265
rect -240 -141275 -185 -141270
rect -280 -141720 220 -141715
rect -280 -141755 -270 -141720
rect -130 -141755 220 -141720
rect -280 -141760 220 -141755
rect -380 -142385 20 -142375
rect -380 -142420 -370 -142385
rect -325 -142420 20 -142385
rect -375 -142430 -320 -142420
rect -600 -142625 100 -142580
rect -600 -144080 -555 -142625
rect -240 -142725 -185 -142720
rect -240 -142730 260 -142725
rect -240 -142765 -235 -142730
rect -190 -142765 260 -142730
rect -240 -142770 260 -142765
rect -240 -142775 -185 -142770
rect -280 -143220 220 -143215
rect -280 -143255 -270 -143220
rect -130 -143255 220 -143220
rect -280 -143260 220 -143255
rect -380 -143885 20 -143875
rect -380 -143920 -370 -143885
rect -325 -143920 20 -143885
rect -375 -143930 -320 -143920
rect -600 -144125 100 -144080
rect -600 -145580 -555 -144125
rect -240 -144225 -185 -144220
rect -240 -144230 260 -144225
rect -240 -144265 -235 -144230
rect -190 -144265 260 -144230
rect -240 -144270 260 -144265
rect -240 -144275 -185 -144270
rect -280 -144720 220 -144715
rect -280 -144755 -270 -144720
rect -130 -144755 220 -144720
rect -280 -144760 220 -144755
rect -380 -145385 20 -145375
rect -380 -145420 -370 -145385
rect -325 -145420 20 -145385
rect -375 -145430 -320 -145420
rect -600 -145625 100 -145580
rect -600 -147080 -555 -145625
rect -240 -145725 -185 -145720
rect -240 -145730 260 -145725
rect -240 -145765 -235 -145730
rect -190 -145765 260 -145730
rect -240 -145770 260 -145765
rect -240 -145775 -185 -145770
rect -280 -146220 220 -146215
rect -280 -146255 -270 -146220
rect -130 -146255 220 -146220
rect -280 -146260 220 -146255
rect -380 -146885 20 -146875
rect -380 -146920 -370 -146885
rect -325 -146920 20 -146885
rect -375 -146930 -320 -146920
rect -600 -147125 100 -147080
rect -600 -147500 -555 -147125
rect -240 -147225 -185 -147220
rect -240 -147230 260 -147225
rect -240 -147265 -235 -147230
rect -190 -147265 260 -147230
rect -240 -147270 260 -147265
rect -240 -147275 -185 -147270
rect -280 -147720 220 -147715
rect -280 -147755 -270 -147720
rect -130 -147755 220 -147720
rect -280 -147760 220 -147755
rect -380 -148385 20 -148375
rect -380 -148420 -370 -148385
rect -325 -148420 20 -148385
rect -375 -148430 -320 -148420
rect 270 -148540 1390 -148530
rect 270 -148590 280 -148540
rect 1380 -148590 1390 -148540
rect 270 -148600 1390 -148590
rect 1770 -148540 2890 -148530
rect 1770 -148590 1780 -148540
rect 2880 -148590 2890 -148540
rect 1770 -148600 2890 -148590
rect 3270 -148540 4390 -148530
rect 3270 -148590 3280 -148540
rect 4380 -148590 4390 -148540
rect 3270 -148600 4390 -148590
rect 4770 -148540 5890 -148530
rect 4770 -148590 4780 -148540
rect 5880 -148590 5890 -148540
rect 4770 -148600 5890 -148590
rect 6270 -148540 7390 -148530
rect 6270 -148590 6280 -148540
rect 7380 -148590 7390 -148540
rect 6270 -148600 7390 -148590
rect 7770 -148540 8890 -148530
rect 7770 -148590 7780 -148540
rect 8880 -148590 8890 -148540
rect 7770 -148600 8890 -148590
rect 9270 -148540 10390 -148530
rect 9270 -148590 9280 -148540
rect 10380 -148590 10390 -148540
rect 9270 -148600 10390 -148590
rect 10770 -148540 11890 -148530
rect 10770 -148590 10780 -148540
rect 11880 -148590 11890 -148540
rect 10770 -148600 11890 -148590
rect 12270 -148540 13390 -148530
rect 12270 -148590 12280 -148540
rect 13380 -148590 13390 -148540
rect 12270 -148600 13390 -148590
rect 13770 -148540 14890 -148530
rect 13770 -148590 13780 -148540
rect 14880 -148590 14890 -148540
rect 13770 -148600 14890 -148590
rect 15270 -148540 16390 -148530
rect 15270 -148590 15280 -148540
rect 16380 -148590 16390 -148540
rect 15270 -148600 16390 -148590
rect 16770 -148540 17890 -148530
rect 16770 -148590 16780 -148540
rect 17880 -148590 17890 -148540
rect 16770 -148600 17890 -148590
rect 18270 -148540 19390 -148530
rect 18270 -148590 18280 -148540
rect 19380 -148590 19390 -148540
rect 18270 -148600 19390 -148590
rect 19770 -148540 20890 -148530
rect 19770 -148590 19780 -148540
rect 20880 -148590 20890 -148540
rect 19770 -148600 20890 -148590
rect 21270 -148540 22390 -148530
rect 21270 -148590 21280 -148540
rect 22380 -148590 22390 -148540
rect 21270 -148600 22390 -148590
rect 22770 -148540 23890 -148530
rect 22770 -148590 22780 -148540
rect 23880 -148590 23890 -148540
rect 22770 -148600 23890 -148590
rect 24270 -148540 25390 -148530
rect 24270 -148590 24280 -148540
rect 25380 -148590 25390 -148540
rect 24270 -148600 25390 -148590
rect 25770 -148540 26890 -148530
rect 25770 -148590 25780 -148540
rect 26880 -148590 26890 -148540
rect 25770 -148600 26890 -148590
rect 27270 -148540 28390 -148530
rect 27270 -148590 27280 -148540
rect 28380 -148590 28390 -148540
rect 27270 -148600 28390 -148590
rect 28770 -148540 29890 -148530
rect 28770 -148590 28780 -148540
rect 29880 -148590 29890 -148540
rect 28770 -148600 29890 -148590
rect 30270 -148540 31390 -148530
rect 30270 -148590 30280 -148540
rect 31380 -148590 31390 -148540
rect 30270 -148600 31390 -148590
rect 31770 -148540 32890 -148530
rect 31770 -148590 31780 -148540
rect 32880 -148590 32890 -148540
rect 31770 -148600 32890 -148590
rect 33270 -148540 34390 -148530
rect 33270 -148590 33280 -148540
rect 34380 -148590 34390 -148540
rect 33270 -148600 34390 -148590
rect 34770 -148540 35890 -148530
rect 34770 -148590 34780 -148540
rect 35880 -148590 35890 -148540
rect 34770 -148600 35890 -148590
rect 36270 -148540 37390 -148530
rect 36270 -148590 36280 -148540
rect 37380 -148590 37390 -148540
rect 36270 -148600 37390 -148590
rect 37770 -148540 38890 -148530
rect 37770 -148590 37780 -148540
rect 38880 -148590 38890 -148540
rect 37770 -148600 38890 -148590
rect 39270 -148540 40390 -148530
rect 39270 -148590 39280 -148540
rect 40380 -148590 40390 -148540
rect 39270 -148600 40390 -148590
rect 40770 -148540 41890 -148530
rect 40770 -148590 40780 -148540
rect 41880 -148590 41890 -148540
rect 40770 -148600 41890 -148590
rect 42270 -148540 43390 -148530
rect 42270 -148590 42280 -148540
rect 43380 -148590 43390 -148540
rect 42270 -148600 43390 -148590
rect 43770 -148540 44890 -148530
rect 43770 -148590 43780 -148540
rect 44880 -148590 44890 -148540
rect 43770 -148600 44890 -148590
rect 45270 -148540 46390 -148530
rect 45270 -148590 45280 -148540
rect 46380 -148590 46390 -148540
rect 45270 -148600 46390 -148590
rect 46770 -148540 47890 -148530
rect 46770 -148590 46780 -148540
rect 47880 -148590 47890 -148540
rect 46770 -148600 47890 -148590
rect 48270 -148540 49390 -148530
rect 48270 -148590 48280 -148540
rect 49380 -148590 49390 -148540
rect 48270 -148600 49390 -148590
rect 49770 -148540 50890 -148530
rect 49770 -148590 49780 -148540
rect 50880 -148590 50890 -148540
rect 49770 -148600 50890 -148590
rect 51270 -148540 52390 -148530
rect 51270 -148590 51280 -148540
rect 52380 -148590 52390 -148540
rect 51270 -148600 52390 -148590
rect 52770 -148540 53890 -148530
rect 52770 -148590 52780 -148540
rect 53880 -148590 53890 -148540
rect 52770 -148600 53890 -148590
rect 54270 -148540 55390 -148530
rect 54270 -148590 54280 -148540
rect 55380 -148590 55390 -148540
rect 54270 -148600 55390 -148590
rect 55770 -148540 56890 -148530
rect 55770 -148590 55780 -148540
rect 56880 -148590 56890 -148540
rect 55770 -148600 56890 -148590
rect 57270 -148540 58390 -148530
rect 57270 -148590 57280 -148540
rect 58380 -148590 58390 -148540
rect 57270 -148600 58390 -148590
rect 58770 -148540 59890 -148530
rect 58770 -148590 58780 -148540
rect 59880 -148590 59890 -148540
rect 58770 -148600 59890 -148590
rect 60270 -148540 61390 -148530
rect 60270 -148590 60280 -148540
rect 61380 -148590 61390 -148540
rect 60270 -148600 61390 -148590
rect 61770 -148540 62890 -148530
rect 61770 -148590 61780 -148540
rect 62880 -148590 62890 -148540
rect 61770 -148600 62890 -148590
rect 63270 -148540 64390 -148530
rect 63270 -148590 63280 -148540
rect 64380 -148590 64390 -148540
rect 63270 -148600 64390 -148590
rect 64770 -148540 65890 -148530
rect 64770 -148590 64780 -148540
rect 65880 -148590 65890 -148540
rect 64770 -148600 65890 -148590
rect 66270 -148540 67390 -148530
rect 66270 -148590 66280 -148540
rect 67380 -148590 67390 -148540
rect 66270 -148600 67390 -148590
rect 67770 -148540 68890 -148530
rect 67770 -148590 67780 -148540
rect 68880 -148590 68890 -148540
rect 67770 -148600 68890 -148590
rect 69270 -148540 70390 -148530
rect 69270 -148590 69280 -148540
rect 70380 -148590 70390 -148540
rect 69270 -148600 70390 -148590
rect 70770 -148540 71890 -148530
rect 70770 -148590 70780 -148540
rect 71880 -148590 71890 -148540
rect 70770 -148600 71890 -148590
rect 72270 -148540 73390 -148530
rect 72270 -148590 72280 -148540
rect 73380 -148590 73390 -148540
rect 72270 -148600 73390 -148590
rect 73770 -148540 74890 -148530
rect 73770 -148590 73780 -148540
rect 74880 -148590 74890 -148540
rect 73770 -148600 74890 -148590
rect 75270 -148540 76390 -148530
rect 75270 -148590 75280 -148540
rect 76380 -148590 76390 -148540
rect 75270 -148600 76390 -148590
rect 76770 -148540 77890 -148530
rect 76770 -148590 76780 -148540
rect 77880 -148590 77890 -148540
rect 76770 -148600 77890 -148590
rect 78270 -148540 79390 -148530
rect 78270 -148590 78280 -148540
rect 79380 -148590 79390 -148540
rect 78270 -148600 79390 -148590
rect 79770 -148540 80890 -148530
rect 79770 -148590 79780 -148540
rect 80880 -148590 80890 -148540
rect 79770 -148600 80890 -148590
rect 81270 -148540 82390 -148530
rect 81270 -148590 81280 -148540
rect 82380 -148590 82390 -148540
rect 81270 -148600 82390 -148590
rect 82770 -148540 83890 -148530
rect 82770 -148590 82780 -148540
rect 83880 -148590 83890 -148540
rect 82770 -148600 83890 -148590
rect 84270 -148540 85390 -148530
rect 84270 -148590 84280 -148540
rect 85380 -148590 85390 -148540
rect 84270 -148600 85390 -148590
rect 85770 -148540 86890 -148530
rect 85770 -148590 85780 -148540
rect 86880 -148590 86890 -148540
rect 85770 -148600 86890 -148590
rect 87270 -148540 88390 -148530
rect 87270 -148590 87280 -148540
rect 88380 -148590 88390 -148540
rect 87270 -148600 88390 -148590
rect 88770 -148540 89890 -148530
rect 88770 -148590 88780 -148540
rect 89880 -148590 89890 -148540
rect 88770 -148600 89890 -148590
rect 90270 -148540 91390 -148530
rect 90270 -148590 90280 -148540
rect 91380 -148590 91390 -148540
rect 90270 -148600 91390 -148590
rect 91770 -148540 92890 -148530
rect 91770 -148590 91780 -148540
rect 92880 -148590 92890 -148540
rect 91770 -148600 92890 -148590
rect 93270 -148540 94390 -148530
rect 93270 -148590 93280 -148540
rect 94380 -148590 94390 -148540
rect 93270 -148600 94390 -148590
rect 94770 -148540 95890 -148530
rect 94770 -148590 94780 -148540
rect 95880 -148590 95890 -148540
rect 94770 -148600 95890 -148590
rect 96270 -148540 97390 -148530
rect 96270 -148590 96280 -148540
rect 97380 -148590 97390 -148540
rect 96270 -148600 97390 -148590
rect 97770 -148540 98890 -148530
rect 97770 -148590 97780 -148540
rect 98880 -148590 98890 -148540
rect 97770 -148600 98890 -148590
rect 99270 -148540 100390 -148530
rect 99270 -148590 99280 -148540
rect 100380 -148590 100390 -148540
rect 99270 -148600 100390 -148590
rect 100770 -148540 101890 -148530
rect 100770 -148590 100780 -148540
rect 101880 -148590 101890 -148540
rect 100770 -148600 101890 -148590
rect 102270 -148540 103390 -148530
rect 102270 -148590 102280 -148540
rect 103380 -148590 103390 -148540
rect 102270 -148600 103390 -148590
rect 103770 -148540 104890 -148530
rect 103770 -148590 103780 -148540
rect 104880 -148590 104890 -148540
rect 103770 -148600 104890 -148590
rect 105270 -148540 106390 -148530
rect 105270 -148590 105280 -148540
rect 106380 -148590 106390 -148540
rect 105270 -148600 106390 -148590
rect 106770 -148540 107890 -148530
rect 106770 -148590 106780 -148540
rect 107880 -148590 107890 -148540
rect 106770 -148600 107890 -148590
rect 108270 -148540 109390 -148530
rect 108270 -148590 108280 -148540
rect 109380 -148590 109390 -148540
rect 108270 -148600 109390 -148590
rect 109770 -148540 110890 -148530
rect 109770 -148590 109780 -148540
rect 110880 -148590 110890 -148540
rect 109770 -148600 110890 -148590
rect 111270 -148540 112390 -148530
rect 111270 -148590 111280 -148540
rect 112380 -148590 112390 -148540
rect 111270 -148600 112390 -148590
rect 112770 -148540 113890 -148530
rect 112770 -148590 112780 -148540
rect 113880 -148590 113890 -148540
rect 112770 -148600 113890 -148590
rect 114270 -148540 115390 -148530
rect 114270 -148590 114280 -148540
rect 115380 -148590 115390 -148540
rect 114270 -148600 115390 -148590
rect 115770 -148540 116890 -148530
rect 115770 -148590 115780 -148540
rect 116880 -148590 116890 -148540
rect 115770 -148600 116890 -148590
rect 117270 -148540 118390 -148530
rect 117270 -148590 117280 -148540
rect 118380 -148590 118390 -148540
rect 117270 -148600 118390 -148590
rect 118770 -148540 119890 -148530
rect 118770 -148590 118780 -148540
rect 119880 -148590 119890 -148540
rect 118770 -148600 119890 -148590
rect 120270 -148540 121390 -148530
rect 120270 -148590 120280 -148540
rect 121380 -148590 121390 -148540
rect 120270 -148600 121390 -148590
rect 121770 -148540 122890 -148530
rect 121770 -148590 121780 -148540
rect 122880 -148590 122890 -148540
rect 121770 -148600 122890 -148590
rect 123270 -148540 124390 -148530
rect 123270 -148590 123280 -148540
rect 124380 -148590 124390 -148540
rect 123270 -148600 124390 -148590
rect 124770 -148540 125890 -148530
rect 124770 -148590 124780 -148540
rect 125880 -148590 125890 -148540
rect 124770 -148600 125890 -148590
rect 126270 -148540 127390 -148530
rect 126270 -148590 126280 -148540
rect 127380 -148590 127390 -148540
rect 126270 -148600 127390 -148590
rect 127770 -148540 128890 -148530
rect 127770 -148590 127780 -148540
rect 128880 -148590 128890 -148540
rect 127770 -148600 128890 -148590
rect 129270 -148540 130390 -148530
rect 129270 -148590 129280 -148540
rect 130380 -148590 130390 -148540
rect 129270 -148600 130390 -148590
rect 130770 -148540 131890 -148530
rect 130770 -148590 130780 -148540
rect 131880 -148590 131890 -148540
rect 130770 -148600 131890 -148590
rect 132270 -148540 133390 -148530
rect 132270 -148590 132280 -148540
rect 133380 -148590 133390 -148540
rect 132270 -148600 133390 -148590
rect 133770 -148540 134890 -148530
rect 133770 -148590 133780 -148540
rect 134880 -148590 134890 -148540
rect 133770 -148600 134890 -148590
rect 135270 -148540 136390 -148530
rect 135270 -148590 135280 -148540
rect 136380 -148590 136390 -148540
rect 135270 -148600 136390 -148590
rect 136770 -148540 137890 -148530
rect 136770 -148590 136780 -148540
rect 137880 -148590 137890 -148540
rect 136770 -148600 137890 -148590
rect 138270 -148540 139390 -148530
rect 138270 -148590 138280 -148540
rect 139380 -148590 139390 -148540
rect 138270 -148600 139390 -148590
rect 139770 -148540 140890 -148530
rect 139770 -148590 139780 -148540
rect 140880 -148590 140890 -148540
rect 139770 -148600 140890 -148590
rect 141270 -148540 142390 -148530
rect 141270 -148590 141280 -148540
rect 142380 -148590 142390 -148540
rect 141270 -148600 142390 -148590
rect 142770 -148540 143890 -148530
rect 142770 -148590 142780 -148540
rect 143880 -148590 143890 -148540
rect 142770 -148600 143890 -148590
rect 144270 -148540 145390 -148530
rect 144270 -148590 144280 -148540
rect 145380 -148590 145390 -148540
rect 144270 -148600 145390 -148590
rect 145770 -148540 146890 -148530
rect 145770 -148590 145780 -148540
rect 146880 -148590 146890 -148540
rect 145770 -148600 146890 -148590
rect 147270 -148540 148390 -148530
rect 147270 -148590 147280 -148540
rect 148380 -148590 148390 -148540
rect 147270 -148600 148390 -148590
rect 148770 -148540 149890 -148530
rect 148770 -148590 148780 -148540
rect 149880 -148590 149890 -148540
rect 148770 -148600 149890 -148590
rect 110 -148750 220 -148745
rect 110 -148850 120 -148750
rect 210 -148850 220 -148750
rect 110 -148855 220 -148850
rect 1610 -148750 1720 -148745
rect 1610 -148850 1620 -148750
rect 1710 -148850 1720 -148750
rect 1610 -148855 1720 -148850
rect 3110 -148750 3220 -148745
rect 3110 -148850 3120 -148750
rect 3210 -148850 3220 -148750
rect 3110 -148855 3220 -148850
rect 4610 -148750 4720 -148745
rect 4610 -148850 4620 -148750
rect 4710 -148850 4720 -148750
rect 4610 -148855 4720 -148850
rect 6110 -148750 6220 -148745
rect 6110 -148850 6120 -148750
rect 6210 -148850 6220 -148750
rect 6110 -148855 6220 -148850
rect 7610 -148750 7720 -148745
rect 7610 -148850 7620 -148750
rect 7710 -148850 7720 -148750
rect 7610 -148855 7720 -148850
rect 9110 -148750 9220 -148745
rect 9110 -148850 9120 -148750
rect 9210 -148850 9220 -148750
rect 9110 -148855 9220 -148850
rect 10610 -148750 10720 -148745
rect 10610 -148850 10620 -148750
rect 10710 -148850 10720 -148750
rect 10610 -148855 10720 -148850
rect 12110 -148750 12220 -148745
rect 12110 -148850 12120 -148750
rect 12210 -148850 12220 -148750
rect 12110 -148855 12220 -148850
rect 13610 -148750 13720 -148745
rect 13610 -148850 13620 -148750
rect 13710 -148850 13720 -148750
rect 13610 -148855 13720 -148850
rect 15110 -148750 15220 -148745
rect 15110 -148850 15120 -148750
rect 15210 -148850 15220 -148750
rect 15110 -148855 15220 -148850
rect 16610 -148750 16720 -148745
rect 16610 -148850 16620 -148750
rect 16710 -148850 16720 -148750
rect 16610 -148855 16720 -148850
rect 18110 -148750 18220 -148745
rect 18110 -148850 18120 -148750
rect 18210 -148850 18220 -148750
rect 18110 -148855 18220 -148850
rect 19610 -148750 19720 -148745
rect 19610 -148850 19620 -148750
rect 19710 -148850 19720 -148750
rect 19610 -148855 19720 -148850
rect 21110 -148750 21220 -148745
rect 21110 -148850 21120 -148750
rect 21210 -148850 21220 -148750
rect 21110 -148855 21220 -148850
rect 22610 -148750 22720 -148745
rect 22610 -148850 22620 -148750
rect 22710 -148850 22720 -148750
rect 22610 -148855 22720 -148850
rect 24110 -148750 24220 -148745
rect 24110 -148850 24120 -148750
rect 24210 -148850 24220 -148750
rect 24110 -148855 24220 -148850
rect 25610 -148750 25720 -148745
rect 25610 -148850 25620 -148750
rect 25710 -148850 25720 -148750
rect 25610 -148855 25720 -148850
rect 27110 -148750 27220 -148745
rect 27110 -148850 27120 -148750
rect 27210 -148850 27220 -148750
rect 27110 -148855 27220 -148850
rect 28610 -148750 28720 -148745
rect 28610 -148850 28620 -148750
rect 28710 -148850 28720 -148750
rect 28610 -148855 28720 -148850
rect 30110 -148750 30220 -148745
rect 30110 -148850 30120 -148750
rect 30210 -148850 30220 -148750
rect 30110 -148855 30220 -148850
rect 31610 -148750 31720 -148745
rect 31610 -148850 31620 -148750
rect 31710 -148850 31720 -148750
rect 31610 -148855 31720 -148850
rect 33110 -148750 33220 -148745
rect 33110 -148850 33120 -148750
rect 33210 -148850 33220 -148750
rect 33110 -148855 33220 -148850
rect 34610 -148750 34720 -148745
rect 34610 -148850 34620 -148750
rect 34710 -148850 34720 -148750
rect 34610 -148855 34720 -148850
rect 36110 -148750 36220 -148745
rect 36110 -148850 36120 -148750
rect 36210 -148850 36220 -148750
rect 36110 -148855 36220 -148850
rect 37610 -148750 37720 -148745
rect 37610 -148850 37620 -148750
rect 37710 -148850 37720 -148750
rect 37610 -148855 37720 -148850
rect 39110 -148750 39220 -148745
rect 39110 -148850 39120 -148750
rect 39210 -148850 39220 -148750
rect 39110 -148855 39220 -148850
rect 40610 -148750 40720 -148745
rect 40610 -148850 40620 -148750
rect 40710 -148850 40720 -148750
rect 40610 -148855 40720 -148850
rect 42110 -148750 42220 -148745
rect 42110 -148850 42120 -148750
rect 42210 -148850 42220 -148750
rect 42110 -148855 42220 -148850
rect 43610 -148750 43720 -148745
rect 43610 -148850 43620 -148750
rect 43710 -148850 43720 -148750
rect 43610 -148855 43720 -148850
rect 45110 -148750 45220 -148745
rect 45110 -148850 45120 -148750
rect 45210 -148850 45220 -148750
rect 45110 -148855 45220 -148850
rect 46610 -148750 46720 -148745
rect 46610 -148850 46620 -148750
rect 46710 -148850 46720 -148750
rect 46610 -148855 46720 -148850
rect 48110 -148750 48220 -148745
rect 48110 -148850 48120 -148750
rect 48210 -148850 48220 -148750
rect 48110 -148855 48220 -148850
rect 49610 -148750 49720 -148745
rect 49610 -148850 49620 -148750
rect 49710 -148850 49720 -148750
rect 49610 -148855 49720 -148850
rect 51110 -148750 51220 -148745
rect 51110 -148850 51120 -148750
rect 51210 -148850 51220 -148750
rect 51110 -148855 51220 -148850
rect 52610 -148750 52720 -148745
rect 52610 -148850 52620 -148750
rect 52710 -148850 52720 -148750
rect 52610 -148855 52720 -148850
rect 54110 -148750 54220 -148745
rect 54110 -148850 54120 -148750
rect 54210 -148850 54220 -148750
rect 54110 -148855 54220 -148850
rect 55610 -148750 55720 -148745
rect 55610 -148850 55620 -148750
rect 55710 -148850 55720 -148750
rect 55610 -148855 55720 -148850
rect 57110 -148750 57220 -148745
rect 57110 -148850 57120 -148750
rect 57210 -148850 57220 -148750
rect 57110 -148855 57220 -148850
rect 58610 -148750 58720 -148745
rect 58610 -148850 58620 -148750
rect 58710 -148850 58720 -148750
rect 58610 -148855 58720 -148850
rect 60110 -148750 60220 -148745
rect 60110 -148850 60120 -148750
rect 60210 -148850 60220 -148750
rect 60110 -148855 60220 -148850
rect 61610 -148750 61720 -148745
rect 61610 -148850 61620 -148750
rect 61710 -148850 61720 -148750
rect 61610 -148855 61720 -148850
rect 63110 -148750 63220 -148745
rect 63110 -148850 63120 -148750
rect 63210 -148850 63220 -148750
rect 63110 -148855 63220 -148850
rect 64610 -148750 64720 -148745
rect 64610 -148850 64620 -148750
rect 64710 -148850 64720 -148750
rect 64610 -148855 64720 -148850
rect 66110 -148750 66220 -148745
rect 66110 -148850 66120 -148750
rect 66210 -148850 66220 -148750
rect 66110 -148855 66220 -148850
rect 67610 -148750 67720 -148745
rect 67610 -148850 67620 -148750
rect 67710 -148850 67720 -148750
rect 67610 -148855 67720 -148850
rect 69110 -148750 69220 -148745
rect 69110 -148850 69120 -148750
rect 69210 -148850 69220 -148750
rect 69110 -148855 69220 -148850
rect 70610 -148750 70720 -148745
rect 70610 -148850 70620 -148750
rect 70710 -148850 70720 -148750
rect 70610 -148855 70720 -148850
rect 72110 -148750 72220 -148745
rect 72110 -148850 72120 -148750
rect 72210 -148850 72220 -148750
rect 72110 -148855 72220 -148850
rect 73610 -148750 73720 -148745
rect 73610 -148850 73620 -148750
rect 73710 -148850 73720 -148750
rect 73610 -148855 73720 -148850
rect 75110 -148750 75220 -148745
rect 75110 -148850 75120 -148750
rect 75210 -148850 75220 -148750
rect 75110 -148855 75220 -148850
rect 76610 -148750 76720 -148745
rect 76610 -148850 76620 -148750
rect 76710 -148850 76720 -148750
rect 76610 -148855 76720 -148850
rect 78110 -148750 78220 -148745
rect 78110 -148850 78120 -148750
rect 78210 -148850 78220 -148750
rect 78110 -148855 78220 -148850
rect 79610 -148750 79720 -148745
rect 79610 -148850 79620 -148750
rect 79710 -148850 79720 -148750
rect 79610 -148855 79720 -148850
rect 81110 -148750 81220 -148745
rect 81110 -148850 81120 -148750
rect 81210 -148850 81220 -148750
rect 81110 -148855 81220 -148850
rect 82610 -148750 82720 -148745
rect 82610 -148850 82620 -148750
rect 82710 -148850 82720 -148750
rect 82610 -148855 82720 -148850
rect 84110 -148750 84220 -148745
rect 84110 -148850 84120 -148750
rect 84210 -148850 84220 -148750
rect 84110 -148855 84220 -148850
rect 85610 -148750 85720 -148745
rect 85610 -148850 85620 -148750
rect 85710 -148850 85720 -148750
rect 85610 -148855 85720 -148850
rect 87110 -148750 87220 -148745
rect 87110 -148850 87120 -148750
rect 87210 -148850 87220 -148750
rect 87110 -148855 87220 -148850
rect 88610 -148750 88720 -148745
rect 88610 -148850 88620 -148750
rect 88710 -148850 88720 -148750
rect 88610 -148855 88720 -148850
rect 90110 -148750 90220 -148745
rect 90110 -148850 90120 -148750
rect 90210 -148850 90220 -148750
rect 90110 -148855 90220 -148850
rect 91610 -148750 91720 -148745
rect 91610 -148850 91620 -148750
rect 91710 -148850 91720 -148750
rect 91610 -148855 91720 -148850
rect 93110 -148750 93220 -148745
rect 93110 -148850 93120 -148750
rect 93210 -148850 93220 -148750
rect 93110 -148855 93220 -148850
rect 94610 -148750 94720 -148745
rect 94610 -148850 94620 -148750
rect 94710 -148850 94720 -148750
rect 94610 -148855 94720 -148850
rect 96110 -148750 96220 -148745
rect 96110 -148850 96120 -148750
rect 96210 -148850 96220 -148750
rect 96110 -148855 96220 -148850
rect 97610 -148750 97720 -148745
rect 97610 -148850 97620 -148750
rect 97710 -148850 97720 -148750
rect 97610 -148855 97720 -148850
rect 99110 -148750 99220 -148745
rect 99110 -148850 99120 -148750
rect 99210 -148850 99220 -148750
rect 99110 -148855 99220 -148850
rect 100610 -148750 100720 -148745
rect 100610 -148850 100620 -148750
rect 100710 -148850 100720 -148750
rect 100610 -148855 100720 -148850
rect 102110 -148750 102220 -148745
rect 102110 -148850 102120 -148750
rect 102210 -148850 102220 -148750
rect 102110 -148855 102220 -148850
rect 103610 -148750 103720 -148745
rect 103610 -148850 103620 -148750
rect 103710 -148850 103720 -148750
rect 103610 -148855 103720 -148850
rect 105110 -148750 105220 -148745
rect 105110 -148850 105120 -148750
rect 105210 -148850 105220 -148750
rect 105110 -148855 105220 -148850
rect 106610 -148750 106720 -148745
rect 106610 -148850 106620 -148750
rect 106710 -148850 106720 -148750
rect 106610 -148855 106720 -148850
rect 108110 -148750 108220 -148745
rect 108110 -148850 108120 -148750
rect 108210 -148850 108220 -148750
rect 108110 -148855 108220 -148850
rect 109610 -148750 109720 -148745
rect 109610 -148850 109620 -148750
rect 109710 -148850 109720 -148750
rect 109610 -148855 109720 -148850
rect 111110 -148750 111220 -148745
rect 111110 -148850 111120 -148750
rect 111210 -148850 111220 -148750
rect 111110 -148855 111220 -148850
rect 112610 -148750 112720 -148745
rect 112610 -148850 112620 -148750
rect 112710 -148850 112720 -148750
rect 112610 -148855 112720 -148850
rect 114110 -148750 114220 -148745
rect 114110 -148850 114120 -148750
rect 114210 -148850 114220 -148750
rect 114110 -148855 114220 -148850
rect 115610 -148750 115720 -148745
rect 115610 -148850 115620 -148750
rect 115710 -148850 115720 -148750
rect 115610 -148855 115720 -148850
rect 117110 -148750 117220 -148745
rect 117110 -148850 117120 -148750
rect 117210 -148850 117220 -148750
rect 117110 -148855 117220 -148850
rect 118610 -148750 118720 -148745
rect 118610 -148850 118620 -148750
rect 118710 -148850 118720 -148750
rect 118610 -148855 118720 -148850
rect 120110 -148750 120220 -148745
rect 120110 -148850 120120 -148750
rect 120210 -148850 120220 -148750
rect 120110 -148855 120220 -148850
rect 121610 -148750 121720 -148745
rect 121610 -148850 121620 -148750
rect 121710 -148850 121720 -148750
rect 121610 -148855 121720 -148850
rect 123110 -148750 123220 -148745
rect 123110 -148850 123120 -148750
rect 123210 -148850 123220 -148750
rect 123110 -148855 123220 -148850
rect 124610 -148750 124720 -148745
rect 124610 -148850 124620 -148750
rect 124710 -148850 124720 -148750
rect 124610 -148855 124720 -148850
rect 126110 -148750 126220 -148745
rect 126110 -148850 126120 -148750
rect 126210 -148850 126220 -148750
rect 126110 -148855 126220 -148850
rect 127610 -148750 127720 -148745
rect 127610 -148850 127620 -148750
rect 127710 -148850 127720 -148750
rect 127610 -148855 127720 -148850
rect 129110 -148750 129220 -148745
rect 129110 -148850 129120 -148750
rect 129210 -148850 129220 -148750
rect 129110 -148855 129220 -148850
rect 130610 -148750 130720 -148745
rect 130610 -148850 130620 -148750
rect 130710 -148850 130720 -148750
rect 130610 -148855 130720 -148850
rect 132110 -148750 132220 -148745
rect 132110 -148850 132120 -148750
rect 132210 -148850 132220 -148750
rect 132110 -148855 132220 -148850
rect 133610 -148750 133720 -148745
rect 133610 -148850 133620 -148750
rect 133710 -148850 133720 -148750
rect 133610 -148855 133720 -148850
rect 135110 -148750 135220 -148745
rect 135110 -148850 135120 -148750
rect 135210 -148850 135220 -148750
rect 135110 -148855 135220 -148850
rect 136610 -148750 136720 -148745
rect 136610 -148850 136620 -148750
rect 136710 -148850 136720 -148750
rect 136610 -148855 136720 -148850
rect 138110 -148750 138220 -148745
rect 138110 -148850 138120 -148750
rect 138210 -148850 138220 -148750
rect 138110 -148855 138220 -148850
rect 139610 -148750 139720 -148745
rect 139610 -148850 139620 -148750
rect 139710 -148850 139720 -148750
rect 139610 -148855 139720 -148850
rect 141110 -148750 141220 -148745
rect 141110 -148850 141120 -148750
rect 141210 -148850 141220 -148750
rect 141110 -148855 141220 -148850
rect 142610 -148750 142720 -148745
rect 142610 -148850 142620 -148750
rect 142710 -148850 142720 -148750
rect 142610 -148855 142720 -148850
rect 144110 -148750 144220 -148745
rect 144110 -148850 144120 -148750
rect 144210 -148850 144220 -148750
rect 144110 -148855 144220 -148850
rect 145610 -148750 145720 -148745
rect 145610 -148850 145620 -148750
rect 145710 -148850 145720 -148750
rect 145610 -148855 145720 -148850
rect 147110 -148750 147220 -148745
rect 147110 -148850 147120 -148750
rect 147210 -148850 147220 -148750
rect 147110 -148855 147220 -148850
rect 148610 -148750 148720 -148745
rect 148610 -148850 148620 -148750
rect 148710 -148850 148720 -148750
rect 148610 -148855 148720 -148850
<< via3 >>
rect 245 1780 290 1825
rect 1745 1780 1790 1825
rect 3245 1780 3290 1825
rect 4745 1780 4790 1825
rect 6245 1780 6290 1825
rect 7745 1780 7790 1825
rect 9245 1780 9290 1825
rect 10745 1780 10790 1825
rect 12245 1780 12290 1825
rect 13745 1780 13790 1825
rect 15245 1780 15290 1825
rect 16745 1780 16790 1825
rect 18245 1780 18290 1825
rect 19745 1780 19790 1825
rect 21245 1780 21290 1825
rect 22745 1780 22790 1825
rect 24245 1780 24290 1825
rect 25745 1780 25790 1825
rect 27245 1780 27290 1825
rect 28745 1780 28790 1825
rect 30245 1780 30290 1825
rect 31745 1780 31790 1825
rect 33245 1780 33290 1825
rect 34745 1780 34790 1825
rect 36245 1780 36290 1825
rect 37745 1780 37790 1825
rect 39245 1780 39290 1825
rect 40745 1780 40790 1825
rect 42245 1780 42290 1825
rect 43745 1780 43790 1825
rect 45245 1780 45290 1825
rect 46745 1780 46790 1825
rect 48245 1780 48290 1825
rect 49745 1780 49790 1825
rect 51245 1780 51290 1825
rect 52745 1780 52790 1825
rect 54245 1780 54290 1825
rect 55745 1780 55790 1825
rect 57245 1780 57290 1825
rect 58745 1780 58790 1825
rect 60245 1780 60290 1825
rect 61745 1780 61790 1825
rect 63245 1780 63290 1825
rect 64745 1780 64790 1825
rect 66245 1780 66290 1825
rect 67745 1780 67790 1825
rect 69245 1780 69290 1825
rect 70745 1780 70790 1825
rect 72245 1780 72290 1825
rect 73745 1780 73790 1825
rect 75245 1780 75290 1825
rect 76745 1780 76790 1825
rect 78245 1780 78290 1825
rect 79745 1780 79790 1825
rect 81245 1780 81290 1825
rect 82745 1780 82790 1825
rect 84245 1780 84290 1825
rect 85745 1780 85790 1825
rect 87245 1780 87290 1825
rect 88745 1780 88790 1825
rect 90245 1780 90290 1825
rect 91745 1780 91790 1825
rect 93245 1780 93290 1825
rect 94745 1780 94790 1825
rect 96245 1780 96290 1825
rect 97745 1780 97790 1825
rect 99245 1780 99290 1825
rect 100745 1780 100790 1825
rect 102245 1780 102290 1825
rect 103745 1780 103790 1825
rect 105245 1780 105290 1825
rect 106745 1780 106790 1825
rect 108245 1780 108290 1825
rect 109745 1780 109790 1825
rect 111245 1780 111290 1825
rect 112745 1780 112790 1825
rect 114245 1780 114290 1825
rect 115745 1780 115790 1825
rect 117245 1780 117290 1825
rect 118745 1780 118790 1825
rect 120245 1780 120290 1825
rect 121745 1780 121790 1825
rect 123245 1780 123290 1825
rect 124745 1780 124790 1825
rect 126245 1780 126290 1825
rect 127745 1780 127790 1825
rect 129245 1780 129290 1825
rect 130745 1780 130790 1825
rect 132245 1780 132290 1825
rect 133745 1780 133790 1825
rect 135245 1780 135290 1825
rect 136745 1780 136790 1825
rect 138245 1780 138290 1825
rect 139745 1780 139790 1825
rect 141245 1780 141290 1825
rect 142745 1780 142790 1825
rect 144245 1780 144290 1825
rect 145745 1780 145790 1825
rect 147245 1780 147290 1825
rect 148745 1780 148790 1825
rect -235 1235 -190 1270
rect -235 -265 -190 -230
rect -235 -1765 -190 -1730
rect -235 -3265 -190 -3230
rect -235 -4765 -190 -4730
rect -235 -6265 -190 -6230
rect -235 -7765 -190 -7730
rect -235 -9265 -190 -9230
rect -235 -10765 -190 -10730
rect -235 -12265 -190 -12230
rect -235 -13765 -190 -13730
rect -235 -15265 -190 -15230
rect -235 -16765 -190 -16730
rect -235 -18265 -190 -18230
rect -235 -19765 -190 -19730
rect -235 -21265 -190 -21230
rect -235 -22765 -190 -22730
rect -235 -24265 -190 -24230
rect -235 -25765 -190 -25730
rect -235 -27265 -190 -27230
rect -235 -28765 -190 -28730
rect -235 -30265 -190 -30230
rect -235 -31765 -190 -31730
rect -235 -33265 -190 -33230
rect -235 -34765 -190 -34730
rect -235 -36265 -190 -36230
rect -235 -37765 -190 -37730
rect -235 -39265 -190 -39230
rect -235 -40765 -190 -40730
rect -235 -42265 -190 -42230
rect -235 -43765 -190 -43730
rect -235 -45265 -190 -45230
rect -235 -46765 -190 -46730
rect -235 -48265 -190 -48230
rect -235 -49765 -190 -49730
rect -235 -51265 -190 -51230
rect -235 -52765 -190 -52730
rect -235 -54265 -190 -54230
rect -235 -55765 -190 -55730
rect -235 -57265 -190 -57230
rect -235 -58765 -190 -58730
rect -235 -60265 -190 -60230
rect -235 -61765 -190 -61730
rect -235 -63265 -190 -63230
rect -235 -64765 -190 -64730
rect -235 -66265 -190 -66230
rect -235 -67765 -190 -67730
rect -235 -69265 -190 -69230
rect -235 -70765 -190 -70730
rect -235 -72265 -190 -72230
rect -235 -73765 -190 -73730
rect -235 -75265 -190 -75230
rect -235 -76765 -190 -76730
rect -235 -78265 -190 -78230
rect -235 -79765 -190 -79730
rect -235 -81265 -190 -81230
rect -235 -82765 -190 -82730
rect -235 -84265 -190 -84230
rect -235 -85765 -190 -85730
rect -235 -87265 -190 -87230
rect -235 -88765 -190 -88730
rect -235 -90265 -190 -90230
rect -235 -91765 -190 -91730
rect -235 -93265 -190 -93230
rect -235 -94765 -190 -94730
rect -235 -96265 -190 -96230
rect -235 -97765 -190 -97730
rect -235 -99265 -190 -99230
rect -235 -100765 -190 -100730
rect -235 -102265 -190 -102230
rect -235 -103765 -190 -103730
rect -235 -105265 -190 -105230
rect -235 -106765 -190 -106730
rect -235 -108265 -190 -108230
rect -235 -109765 -190 -109730
rect -235 -111265 -190 -111230
rect -235 -112765 -190 -112730
rect -235 -114265 -190 -114230
rect -235 -115765 -190 -115730
rect -235 -117265 -190 -117230
rect -235 -118765 -190 -118730
rect -235 -120265 -190 -120230
rect -235 -121765 -190 -121730
rect -235 -123265 -190 -123230
rect -235 -124765 -190 -124730
rect -235 -126265 -190 -126230
rect -235 -127765 -190 -127730
rect -235 -129265 -190 -129230
rect -235 -130765 -190 -130730
rect -235 -132265 -190 -132230
rect -235 -133765 -190 -133730
rect -235 -135265 -190 -135230
rect -235 -136765 -190 -136730
rect -235 -138265 -190 -138230
rect -235 -139765 -190 -139730
rect -235 -141265 -190 -141230
rect -235 -142765 -190 -142730
rect -235 -144265 -190 -144230
rect -235 -145765 -190 -145730
rect -235 -147265 -190 -147230
rect 280 -148590 1380 -148540
rect 1780 -148590 2880 -148540
rect 3280 -148590 4380 -148540
rect 4780 -148590 5880 -148540
rect 6280 -148590 7380 -148540
rect 7780 -148590 8880 -148540
rect 9280 -148590 10380 -148540
rect 10780 -148590 11880 -148540
rect 12280 -148590 13380 -148540
rect 13780 -148590 14880 -148540
rect 15280 -148590 16380 -148540
rect 16780 -148590 17880 -148540
rect 18280 -148590 19380 -148540
rect 19780 -148590 20880 -148540
rect 21280 -148590 22380 -148540
rect 22780 -148590 23880 -148540
rect 24280 -148590 25380 -148540
rect 25780 -148590 26880 -148540
rect 27280 -148590 28380 -148540
rect 28780 -148590 29880 -148540
rect 30280 -148590 31380 -148540
rect 31780 -148590 32880 -148540
rect 33280 -148590 34380 -148540
rect 34780 -148590 35880 -148540
rect 36280 -148590 37380 -148540
rect 37780 -148590 38880 -148540
rect 39280 -148590 40380 -148540
rect 40780 -148590 41880 -148540
rect 42280 -148590 43380 -148540
rect 43780 -148590 44880 -148540
rect 45280 -148590 46380 -148540
rect 46780 -148590 47880 -148540
rect 48280 -148590 49380 -148540
rect 49780 -148590 50880 -148540
rect 51280 -148590 52380 -148540
rect 52780 -148590 53880 -148540
rect 54280 -148590 55380 -148540
rect 55780 -148590 56880 -148540
rect 57280 -148590 58380 -148540
rect 58780 -148590 59880 -148540
rect 60280 -148590 61380 -148540
rect 61780 -148590 62880 -148540
rect 63280 -148590 64380 -148540
rect 64780 -148590 65880 -148540
rect 66280 -148590 67380 -148540
rect 67780 -148590 68880 -148540
rect 69280 -148590 70380 -148540
rect 70780 -148590 71880 -148540
rect 72280 -148590 73380 -148540
rect 73780 -148590 74880 -148540
rect 75280 -148590 76380 -148540
rect 76780 -148590 77880 -148540
rect 78280 -148590 79380 -148540
rect 79780 -148590 80880 -148540
rect 81280 -148590 82380 -148540
rect 82780 -148590 83880 -148540
rect 84280 -148590 85380 -148540
rect 85780 -148590 86880 -148540
rect 87280 -148590 88380 -148540
rect 88780 -148590 89880 -148540
rect 90280 -148590 91380 -148540
rect 91780 -148590 92880 -148540
rect 93280 -148590 94380 -148540
rect 94780 -148590 95880 -148540
rect 96280 -148590 97380 -148540
rect 97780 -148590 98880 -148540
rect 99280 -148590 100380 -148540
rect 100780 -148590 101880 -148540
rect 102280 -148590 103380 -148540
rect 103780 -148590 104880 -148540
rect 105280 -148590 106380 -148540
rect 106780 -148590 107880 -148540
rect 108280 -148590 109380 -148540
rect 109780 -148590 110880 -148540
rect 111280 -148590 112380 -148540
rect 112780 -148590 113880 -148540
rect 114280 -148590 115380 -148540
rect 115780 -148590 116880 -148540
rect 117280 -148590 118380 -148540
rect 118780 -148590 119880 -148540
rect 120280 -148590 121380 -148540
rect 121780 -148590 122880 -148540
rect 123280 -148590 124380 -148540
rect 124780 -148590 125880 -148540
rect 126280 -148590 127380 -148540
rect 127780 -148590 128880 -148540
rect 129280 -148590 130380 -148540
rect 130780 -148590 131880 -148540
rect 132280 -148590 133380 -148540
rect 133780 -148590 134880 -148540
rect 135280 -148590 136380 -148540
rect 136780 -148590 137880 -148540
rect 138280 -148590 139380 -148540
rect 139780 -148590 140880 -148540
rect 141280 -148590 142380 -148540
rect 142780 -148590 143880 -148540
rect 144280 -148590 145380 -148540
rect 145780 -148590 146880 -148540
rect 147280 -148590 148380 -148540
rect 148780 -148590 149880 -148540
rect 120 -148850 210 -148750
rect 1620 -148850 1710 -148750
rect 3120 -148850 3210 -148750
rect 4620 -148850 4710 -148750
rect 6120 -148850 6210 -148750
rect 7620 -148850 7710 -148750
rect 9120 -148850 9210 -148750
rect 10620 -148850 10710 -148750
rect 12120 -148850 12210 -148750
rect 13620 -148850 13710 -148750
rect 15120 -148850 15210 -148750
rect 16620 -148850 16710 -148750
rect 18120 -148850 18210 -148750
rect 19620 -148850 19710 -148750
rect 21120 -148850 21210 -148750
rect 22620 -148850 22710 -148750
rect 24120 -148850 24210 -148750
rect 25620 -148850 25710 -148750
rect 27120 -148850 27210 -148750
rect 28620 -148850 28710 -148750
rect 30120 -148850 30210 -148750
rect 31620 -148850 31710 -148750
rect 33120 -148850 33210 -148750
rect 34620 -148850 34710 -148750
rect 36120 -148850 36210 -148750
rect 37620 -148850 37710 -148750
rect 39120 -148850 39210 -148750
rect 40620 -148850 40710 -148750
rect 42120 -148850 42210 -148750
rect 43620 -148850 43710 -148750
rect 45120 -148850 45210 -148750
rect 46620 -148850 46710 -148750
rect 48120 -148850 48210 -148750
rect 49620 -148850 49710 -148750
rect 51120 -148850 51210 -148750
rect 52620 -148850 52710 -148750
rect 54120 -148850 54210 -148750
rect 55620 -148850 55710 -148750
rect 57120 -148850 57210 -148750
rect 58620 -148850 58710 -148750
rect 60120 -148850 60210 -148750
rect 61620 -148850 61710 -148750
rect 63120 -148850 63210 -148750
rect 64620 -148850 64710 -148750
rect 66120 -148850 66210 -148750
rect 67620 -148850 67710 -148750
rect 69120 -148850 69210 -148750
rect 70620 -148850 70710 -148750
rect 72120 -148850 72210 -148750
rect 73620 -148850 73710 -148750
rect 75120 -148850 75210 -148750
rect 76620 -148850 76710 -148750
rect 78120 -148850 78210 -148750
rect 79620 -148850 79710 -148750
rect 81120 -148850 81210 -148750
rect 82620 -148850 82710 -148750
rect 84120 -148850 84210 -148750
rect 85620 -148850 85710 -148750
rect 87120 -148850 87210 -148750
rect 88620 -148850 88710 -148750
rect 90120 -148850 90210 -148750
rect 91620 -148850 91710 -148750
rect 93120 -148850 93210 -148750
rect 94620 -148850 94710 -148750
rect 96120 -148850 96210 -148750
rect 97620 -148850 97710 -148750
rect 99120 -148850 99210 -148750
rect 100620 -148850 100710 -148750
rect 102120 -148850 102210 -148750
rect 103620 -148850 103710 -148750
rect 105120 -148850 105210 -148750
rect 106620 -148850 106710 -148750
rect 108120 -148850 108210 -148750
rect 109620 -148850 109710 -148750
rect 111120 -148850 111210 -148750
rect 112620 -148850 112710 -148750
rect 114120 -148850 114210 -148750
rect 115620 -148850 115710 -148750
rect 117120 -148850 117210 -148750
rect 118620 -148850 118710 -148750
rect 120120 -148850 120210 -148750
rect 121620 -148850 121710 -148750
rect 123120 -148850 123210 -148750
rect 124620 -148850 124710 -148750
rect 126120 -148850 126210 -148750
rect 127620 -148850 127710 -148750
rect 129120 -148850 129210 -148750
rect 130620 -148850 130710 -148750
rect 132120 -148850 132210 -148750
rect 133620 -148850 133710 -148750
rect 135120 -148850 135210 -148750
rect 136620 -148850 136710 -148750
rect 138120 -148850 138210 -148750
rect 139620 -148850 139710 -148750
rect 141120 -148850 141210 -148750
rect 142620 -148850 142710 -148750
rect 144120 -148850 144210 -148750
rect 145620 -148850 145710 -148750
rect 147120 -148850 147210 -148750
rect 148620 -148850 148710 -148750
<< metal4 >>
rect -1500 1825 149600 1830
rect -1500 1780 245 1825
rect 290 1780 1745 1825
rect 1790 1780 3245 1825
rect 3290 1780 4745 1825
rect 4790 1780 6245 1825
rect 6290 1780 7745 1825
rect 7790 1780 9245 1825
rect 9290 1780 10745 1825
rect 10790 1780 12245 1825
rect 12290 1780 13745 1825
rect 13790 1780 15245 1825
rect 15290 1780 16745 1825
rect 16790 1780 18245 1825
rect 18290 1780 19745 1825
rect 19790 1780 21245 1825
rect 21290 1780 22745 1825
rect 22790 1780 24245 1825
rect 24290 1780 25745 1825
rect 25790 1780 27245 1825
rect 27290 1780 28745 1825
rect 28790 1780 30245 1825
rect 30290 1780 31745 1825
rect 31790 1780 33245 1825
rect 33290 1780 34745 1825
rect 34790 1780 36245 1825
rect 36290 1780 37745 1825
rect 37790 1780 39245 1825
rect 39290 1780 40745 1825
rect 40790 1780 42245 1825
rect 42290 1780 43745 1825
rect 43790 1780 45245 1825
rect 45290 1780 46745 1825
rect 46790 1780 48245 1825
rect 48290 1780 49745 1825
rect 49790 1780 51245 1825
rect 51290 1780 52745 1825
rect 52790 1780 54245 1825
rect 54290 1780 55745 1825
rect 55790 1780 57245 1825
rect 57290 1780 58745 1825
rect 58790 1780 60245 1825
rect 60290 1780 61745 1825
rect 61790 1780 63245 1825
rect 63290 1780 64745 1825
rect 64790 1780 66245 1825
rect 66290 1780 67745 1825
rect 67790 1780 69245 1825
rect 69290 1780 70745 1825
rect 70790 1780 72245 1825
rect 72290 1780 73745 1825
rect 73790 1780 75245 1825
rect 75290 1780 76745 1825
rect 76790 1780 78245 1825
rect 78290 1780 79745 1825
rect 79790 1780 81245 1825
rect 81290 1780 82745 1825
rect 82790 1780 84245 1825
rect 84290 1780 85745 1825
rect 85790 1780 87245 1825
rect 87290 1780 88745 1825
rect 88790 1780 90245 1825
rect 90290 1780 91745 1825
rect 91790 1780 93245 1825
rect 93290 1780 94745 1825
rect 94790 1780 96245 1825
rect 96290 1780 97745 1825
rect 97790 1780 99245 1825
rect 99290 1780 100745 1825
rect 100790 1780 102245 1825
rect 102290 1780 103745 1825
rect 103790 1780 105245 1825
rect 105290 1780 106745 1825
rect 106790 1780 108245 1825
rect 108290 1780 109745 1825
rect 109790 1780 111245 1825
rect 111290 1780 112745 1825
rect 112790 1780 114245 1825
rect 114290 1780 115745 1825
rect 115790 1780 117245 1825
rect 117290 1780 118745 1825
rect 118790 1780 120245 1825
rect 120290 1780 121745 1825
rect 121790 1780 123245 1825
rect 123290 1780 124745 1825
rect 124790 1780 126245 1825
rect 126290 1780 127745 1825
rect 127790 1780 129245 1825
rect 129290 1780 130745 1825
rect 130790 1780 132245 1825
rect 132290 1780 133745 1825
rect 133790 1780 135245 1825
rect 135290 1780 136745 1825
rect 136790 1780 138245 1825
rect 138290 1780 139745 1825
rect 139790 1780 141245 1825
rect 141290 1780 142745 1825
rect 142790 1780 144245 1825
rect 144290 1780 145745 1825
rect 145790 1780 147245 1825
rect 147290 1780 148745 1825
rect 148790 1780 149600 1825
rect -1500 1775 149600 1780
rect -240 1270 -185 1300
rect -240 1235 -235 1270
rect -190 1235 -185 1270
rect -240 -230 -185 1235
rect -240 -265 -235 -230
rect -190 -265 -185 -230
rect -240 -1730 -185 -265
rect -240 -1765 -235 -1730
rect -190 -1765 -185 -1730
rect -240 -3230 -185 -1765
rect -240 -3265 -235 -3230
rect -190 -3265 -185 -3230
rect -240 -4730 -185 -3265
rect -240 -4765 -235 -4730
rect -190 -4765 -185 -4730
rect -240 -6230 -185 -4765
rect -240 -6265 -235 -6230
rect -190 -6265 -185 -6230
rect -240 -7730 -185 -6265
rect -240 -7765 -235 -7730
rect -190 -7765 -185 -7730
rect -240 -9230 -185 -7765
rect -240 -9265 -235 -9230
rect -190 -9265 -185 -9230
rect -240 -10730 -185 -9265
rect -240 -10765 -235 -10730
rect -190 -10765 -185 -10730
rect -240 -12230 -185 -10765
rect -240 -12265 -235 -12230
rect -190 -12265 -185 -12230
rect -240 -13730 -185 -12265
rect -240 -13765 -235 -13730
rect -190 -13765 -185 -13730
rect -240 -15230 -185 -13765
rect -240 -15265 -235 -15230
rect -190 -15265 -185 -15230
rect -240 -16730 -185 -15265
rect -240 -16765 -235 -16730
rect -190 -16765 -185 -16730
rect -240 -18230 -185 -16765
rect -240 -18265 -235 -18230
rect -190 -18265 -185 -18230
rect -240 -19730 -185 -18265
rect -240 -19765 -235 -19730
rect -190 -19765 -185 -19730
rect -240 -21230 -185 -19765
rect -240 -21265 -235 -21230
rect -190 -21265 -185 -21230
rect -240 -22730 -185 -21265
rect -240 -22765 -235 -22730
rect -190 -22765 -185 -22730
rect -240 -24230 -185 -22765
rect -240 -24265 -235 -24230
rect -190 -24265 -185 -24230
rect -240 -25730 -185 -24265
rect -240 -25765 -235 -25730
rect -190 -25765 -185 -25730
rect -240 -27230 -185 -25765
rect -240 -27265 -235 -27230
rect -190 -27265 -185 -27230
rect -240 -28730 -185 -27265
rect -240 -28765 -235 -28730
rect -190 -28765 -185 -28730
rect -240 -30230 -185 -28765
rect -240 -30265 -235 -30230
rect -190 -30265 -185 -30230
rect -240 -31730 -185 -30265
rect -240 -31765 -235 -31730
rect -190 -31765 -185 -31730
rect -240 -33230 -185 -31765
rect -240 -33265 -235 -33230
rect -190 -33265 -185 -33230
rect -240 -34730 -185 -33265
rect -240 -34765 -235 -34730
rect -190 -34765 -185 -34730
rect -240 -36230 -185 -34765
rect -240 -36265 -235 -36230
rect -190 -36265 -185 -36230
rect -240 -37730 -185 -36265
rect -240 -37765 -235 -37730
rect -190 -37765 -185 -37730
rect -240 -39230 -185 -37765
rect -240 -39265 -235 -39230
rect -190 -39265 -185 -39230
rect -240 -40730 -185 -39265
rect -240 -40765 -235 -40730
rect -190 -40765 -185 -40730
rect -240 -42230 -185 -40765
rect -240 -42265 -235 -42230
rect -190 -42265 -185 -42230
rect -240 -43730 -185 -42265
rect -240 -43765 -235 -43730
rect -190 -43765 -185 -43730
rect -240 -45230 -185 -43765
rect -240 -45265 -235 -45230
rect -190 -45265 -185 -45230
rect -240 -46730 -185 -45265
rect -240 -46765 -235 -46730
rect -190 -46765 -185 -46730
rect -240 -48230 -185 -46765
rect -240 -48265 -235 -48230
rect -190 -48265 -185 -48230
rect -240 -49730 -185 -48265
rect -240 -49765 -235 -49730
rect -190 -49765 -185 -49730
rect -240 -51230 -185 -49765
rect -240 -51265 -235 -51230
rect -190 -51265 -185 -51230
rect -240 -52730 -185 -51265
rect -240 -52765 -235 -52730
rect -190 -52765 -185 -52730
rect -240 -54230 -185 -52765
rect -240 -54265 -235 -54230
rect -190 -54265 -185 -54230
rect -240 -55730 -185 -54265
rect -240 -55765 -235 -55730
rect -190 -55765 -185 -55730
rect -240 -57230 -185 -55765
rect -240 -57265 -235 -57230
rect -190 -57265 -185 -57230
rect -240 -58730 -185 -57265
rect -240 -58765 -235 -58730
rect -190 -58765 -185 -58730
rect -240 -60230 -185 -58765
rect -240 -60265 -235 -60230
rect -190 -60265 -185 -60230
rect -240 -61730 -185 -60265
rect -240 -61765 -235 -61730
rect -190 -61765 -185 -61730
rect -240 -63230 -185 -61765
rect -240 -63265 -235 -63230
rect -190 -63265 -185 -63230
rect -240 -64730 -185 -63265
rect -240 -64765 -235 -64730
rect -190 -64765 -185 -64730
rect -240 -66230 -185 -64765
rect -240 -66265 -235 -66230
rect -190 -66265 -185 -66230
rect -240 -67730 -185 -66265
rect -240 -67765 -235 -67730
rect -190 -67765 -185 -67730
rect -240 -69230 -185 -67765
rect -240 -69265 -235 -69230
rect -190 -69265 -185 -69230
rect -240 -70730 -185 -69265
rect -240 -70765 -235 -70730
rect -190 -70765 -185 -70730
rect -240 -72230 -185 -70765
rect -240 -72265 -235 -72230
rect -190 -72265 -185 -72230
rect -240 -73730 -185 -72265
rect -240 -73765 -235 -73730
rect -190 -73765 -185 -73730
rect -240 -75230 -185 -73765
rect -240 -75265 -235 -75230
rect -190 -75265 -185 -75230
rect -240 -76730 -185 -75265
rect -240 -76765 -235 -76730
rect -190 -76765 -185 -76730
rect -240 -78230 -185 -76765
rect -240 -78265 -235 -78230
rect -190 -78265 -185 -78230
rect -240 -79730 -185 -78265
rect -240 -79765 -235 -79730
rect -190 -79765 -185 -79730
rect -240 -81230 -185 -79765
rect -240 -81265 -235 -81230
rect -190 -81265 -185 -81230
rect -240 -82730 -185 -81265
rect -240 -82765 -235 -82730
rect -190 -82765 -185 -82730
rect -240 -84230 -185 -82765
rect -240 -84265 -235 -84230
rect -190 -84265 -185 -84230
rect -240 -85730 -185 -84265
rect -240 -85765 -235 -85730
rect -190 -85765 -185 -85730
rect -240 -87230 -185 -85765
rect -240 -87265 -235 -87230
rect -190 -87265 -185 -87230
rect -240 -88730 -185 -87265
rect -240 -88765 -235 -88730
rect -190 -88765 -185 -88730
rect -240 -90230 -185 -88765
rect -240 -90265 -235 -90230
rect -190 -90265 -185 -90230
rect -240 -91730 -185 -90265
rect -240 -91765 -235 -91730
rect -190 -91765 -185 -91730
rect -240 -93230 -185 -91765
rect -240 -93265 -235 -93230
rect -190 -93265 -185 -93230
rect -240 -94730 -185 -93265
rect -240 -94765 -235 -94730
rect -190 -94765 -185 -94730
rect -240 -96230 -185 -94765
rect -240 -96265 -235 -96230
rect -190 -96265 -185 -96230
rect -240 -97730 -185 -96265
rect -240 -97765 -235 -97730
rect -190 -97765 -185 -97730
rect -240 -99230 -185 -97765
rect -240 -99265 -235 -99230
rect -190 -99265 -185 -99230
rect -240 -100730 -185 -99265
rect -240 -100765 -235 -100730
rect -190 -100765 -185 -100730
rect -240 -102230 -185 -100765
rect -240 -102265 -235 -102230
rect -190 -102265 -185 -102230
rect -240 -103730 -185 -102265
rect -240 -103765 -235 -103730
rect -190 -103765 -185 -103730
rect -240 -105230 -185 -103765
rect -240 -105265 -235 -105230
rect -190 -105265 -185 -105230
rect -240 -106730 -185 -105265
rect -240 -106765 -235 -106730
rect -190 -106765 -185 -106730
rect -240 -108230 -185 -106765
rect -240 -108265 -235 -108230
rect -190 -108265 -185 -108230
rect -240 -109730 -185 -108265
rect -240 -109765 -235 -109730
rect -190 -109765 -185 -109730
rect -240 -111230 -185 -109765
rect -240 -111265 -235 -111230
rect -190 -111265 -185 -111230
rect -240 -112730 -185 -111265
rect -240 -112765 -235 -112730
rect -190 -112765 -185 -112730
rect -240 -114230 -185 -112765
rect -240 -114265 -235 -114230
rect -190 -114265 -185 -114230
rect -240 -115730 -185 -114265
rect -240 -115765 -235 -115730
rect -190 -115765 -185 -115730
rect -240 -117230 -185 -115765
rect -240 -117265 -235 -117230
rect -190 -117265 -185 -117230
rect -240 -118730 -185 -117265
rect -240 -118765 -235 -118730
rect -190 -118765 -185 -118730
rect -240 -120230 -185 -118765
rect -240 -120265 -235 -120230
rect -190 -120265 -185 -120230
rect -240 -121730 -185 -120265
rect -240 -121765 -235 -121730
rect -190 -121765 -185 -121730
rect -240 -123230 -185 -121765
rect -240 -123265 -235 -123230
rect -190 -123265 -185 -123230
rect -240 -124730 -185 -123265
rect -240 -124765 -235 -124730
rect -190 -124765 -185 -124730
rect -240 -126230 -185 -124765
rect -240 -126265 -235 -126230
rect -190 -126265 -185 -126230
rect -240 -127730 -185 -126265
rect -240 -127765 -235 -127730
rect -190 -127765 -185 -127730
rect -240 -129230 -185 -127765
rect -240 -129265 -235 -129230
rect -190 -129265 -185 -129230
rect -240 -130730 -185 -129265
rect -240 -130765 -235 -130730
rect -190 -130765 -185 -130730
rect -240 -132230 -185 -130765
rect -240 -132265 -235 -132230
rect -190 -132265 -185 -132230
rect -240 -133730 -185 -132265
rect -240 -133765 -235 -133730
rect -190 -133765 -185 -133730
rect -240 -135230 -185 -133765
rect -240 -135265 -235 -135230
rect -190 -135265 -185 -135230
rect -240 -136730 -185 -135265
rect -240 -136765 -235 -136730
rect -190 -136765 -185 -136730
rect -240 -138230 -185 -136765
rect -240 -138265 -235 -138230
rect -190 -138265 -185 -138230
rect -240 -139730 -185 -138265
rect -240 -139765 -235 -139730
rect -190 -139765 -185 -139730
rect -240 -141230 -185 -139765
rect -240 -141265 -235 -141230
rect -190 -141265 -185 -141230
rect -240 -142730 -185 -141265
rect -240 -142765 -235 -142730
rect -190 -142765 -185 -142730
rect -240 -144230 -185 -142765
rect -240 -144265 -235 -144230
rect -190 -144265 -185 -144230
rect -240 -145730 -185 -144265
rect -240 -145765 -235 -145730
rect -190 -145765 -185 -145730
rect -240 -147230 -185 -145765
rect -240 -147265 -235 -147230
rect -190 -147265 -185 -147230
rect -240 -149300 -185 -147265
rect 1315 -148530 1390 -148500
rect 2815 -148530 2890 -148500
rect 4315 -148530 4390 -148500
rect 5815 -148530 5890 -148500
rect 7315 -148530 7390 -148500
rect 8815 -148530 8890 -148500
rect 10315 -148530 10390 -148500
rect 11815 -148530 11890 -148500
rect 13315 -148530 13390 -148500
rect 14815 -148530 14890 -148500
rect 16315 -148530 16390 -148500
rect 17815 -148530 17890 -148500
rect 19315 -148530 19390 -148500
rect 20815 -148530 20890 -148500
rect 22315 -148530 22390 -148500
rect 23815 -148530 23890 -148500
rect 25315 -148530 25390 -148500
rect 26815 -148530 26890 -148500
rect 28315 -148530 28390 -148500
rect 29815 -148530 29890 -148500
rect 31315 -148530 31390 -148500
rect 32815 -148530 32890 -148500
rect 34315 -148530 34390 -148500
rect 35815 -148530 35890 -148500
rect 37315 -148530 37390 -148500
rect 38815 -148530 38890 -148500
rect 40315 -148530 40390 -148500
rect 41815 -148530 41890 -148500
rect 43315 -148530 43390 -148500
rect 44815 -148530 44890 -148500
rect 46315 -148530 46390 -148500
rect 47815 -148530 47890 -148500
rect 49315 -148530 49390 -148500
rect 50815 -148530 50890 -148500
rect 52315 -148530 52390 -148500
rect 53815 -148530 53890 -148500
rect 55315 -148530 55390 -148500
rect 56815 -148530 56890 -148500
rect 58315 -148530 58390 -148500
rect 59815 -148530 59890 -148500
rect 61315 -148530 61390 -148500
rect 62815 -148530 62890 -148500
rect 64315 -148530 64390 -148500
rect 65815 -148530 65890 -148500
rect 67315 -148530 67390 -148500
rect 68815 -148530 68890 -148500
rect 70315 -148530 70390 -148500
rect 71815 -148530 71890 -148500
rect 73315 -148530 73390 -148500
rect 74815 -148530 74890 -148500
rect 76315 -148530 76390 -148500
rect 77815 -148530 77890 -148500
rect 79315 -148530 79390 -148500
rect 80815 -148530 80890 -148500
rect 82315 -148530 82390 -148500
rect 83815 -148530 83890 -148500
rect 85315 -148530 85390 -148500
rect 86815 -148530 86890 -148500
rect 88315 -148530 88390 -148500
rect 89815 -148530 89890 -148500
rect 91315 -148530 91390 -148500
rect 92815 -148530 92890 -148500
rect 94315 -148530 94390 -148500
rect 95815 -148530 95890 -148500
rect 97315 -148530 97390 -148500
rect 98815 -148530 98890 -148500
rect 100315 -148530 100390 -148500
rect 101815 -148530 101890 -148500
rect 103315 -148530 103390 -148500
rect 104815 -148530 104890 -148500
rect 106315 -148530 106390 -148500
rect 107815 -148530 107890 -148500
rect 109315 -148530 109390 -148500
rect 110815 -148530 110890 -148500
rect 112315 -148530 112390 -148500
rect 113815 -148530 113890 -148500
rect 115315 -148530 115390 -148500
rect 116815 -148530 116890 -148500
rect 118315 -148530 118390 -148500
rect 119815 -148530 119890 -148500
rect 121315 -148530 121390 -148500
rect 122815 -148530 122890 -148500
rect 124315 -148530 124390 -148500
rect 125815 -148530 125890 -148500
rect 127315 -148530 127390 -148500
rect 128815 -148530 128890 -148500
rect 130315 -148530 130390 -148500
rect 131815 -148530 131890 -148500
rect 133315 -148530 133390 -148500
rect 134815 -148530 134890 -148500
rect 136315 -148530 136390 -148500
rect 137815 -148530 137890 -148500
rect 139315 -148530 139390 -148500
rect 140815 -148530 140890 -148500
rect 142315 -148530 142390 -148500
rect 143815 -148530 143890 -148500
rect 145315 -148530 145390 -148500
rect 146815 -148530 146890 -148500
rect 148315 -148530 148390 -148500
rect 149815 -148530 149890 -148500
rect 270 -148540 1390 -148530
rect 270 -148590 280 -148540
rect 1380 -148590 1390 -148540
rect 270 -148600 1390 -148590
rect 1770 -148540 2890 -148530
rect 1770 -148590 1780 -148540
rect 2880 -148590 2890 -148540
rect 1770 -148600 2890 -148590
rect 3270 -148540 4390 -148530
rect 3270 -148590 3280 -148540
rect 4380 -148590 4390 -148540
rect 3270 -148600 4390 -148590
rect 4770 -148540 5890 -148530
rect 4770 -148590 4780 -148540
rect 5880 -148590 5890 -148540
rect 4770 -148600 5890 -148590
rect 6270 -148540 7390 -148530
rect 6270 -148590 6280 -148540
rect 7380 -148590 7390 -148540
rect 6270 -148600 7390 -148590
rect 7770 -148540 8890 -148530
rect 7770 -148590 7780 -148540
rect 8880 -148590 8890 -148540
rect 7770 -148600 8890 -148590
rect 9270 -148540 10390 -148530
rect 9270 -148590 9280 -148540
rect 10380 -148590 10390 -148540
rect 9270 -148600 10390 -148590
rect 10770 -148540 11890 -148530
rect 10770 -148590 10780 -148540
rect 11880 -148590 11890 -148540
rect 10770 -148600 11890 -148590
rect 12270 -148540 13390 -148530
rect 12270 -148590 12280 -148540
rect 13380 -148590 13390 -148540
rect 12270 -148600 13390 -148590
rect 13770 -148540 14890 -148530
rect 13770 -148590 13780 -148540
rect 14880 -148590 14890 -148540
rect 13770 -148600 14890 -148590
rect 15270 -148540 16390 -148530
rect 15270 -148590 15280 -148540
rect 16380 -148590 16390 -148540
rect 15270 -148600 16390 -148590
rect 16770 -148540 17890 -148530
rect 16770 -148590 16780 -148540
rect 17880 -148590 17890 -148540
rect 16770 -148600 17890 -148590
rect 18270 -148540 19390 -148530
rect 18270 -148590 18280 -148540
rect 19380 -148590 19390 -148540
rect 18270 -148600 19390 -148590
rect 19770 -148540 20890 -148530
rect 19770 -148590 19780 -148540
rect 20880 -148590 20890 -148540
rect 19770 -148600 20890 -148590
rect 21270 -148540 22390 -148530
rect 21270 -148590 21280 -148540
rect 22380 -148590 22390 -148540
rect 21270 -148600 22390 -148590
rect 22770 -148540 23890 -148530
rect 22770 -148590 22780 -148540
rect 23880 -148590 23890 -148540
rect 22770 -148600 23890 -148590
rect 24270 -148540 25390 -148530
rect 24270 -148590 24280 -148540
rect 25380 -148590 25390 -148540
rect 24270 -148600 25390 -148590
rect 25770 -148540 26890 -148530
rect 25770 -148590 25780 -148540
rect 26880 -148590 26890 -148540
rect 25770 -148600 26890 -148590
rect 27270 -148540 28390 -148530
rect 27270 -148590 27280 -148540
rect 28380 -148590 28390 -148540
rect 27270 -148600 28390 -148590
rect 28770 -148540 29890 -148530
rect 28770 -148590 28780 -148540
rect 29880 -148590 29890 -148540
rect 28770 -148600 29890 -148590
rect 30270 -148540 31390 -148530
rect 30270 -148590 30280 -148540
rect 31380 -148590 31390 -148540
rect 30270 -148600 31390 -148590
rect 31770 -148540 32890 -148530
rect 31770 -148590 31780 -148540
rect 32880 -148590 32890 -148540
rect 31770 -148600 32890 -148590
rect 33270 -148540 34390 -148530
rect 33270 -148590 33280 -148540
rect 34380 -148590 34390 -148540
rect 33270 -148600 34390 -148590
rect 34770 -148540 35890 -148530
rect 34770 -148590 34780 -148540
rect 35880 -148590 35890 -148540
rect 34770 -148600 35890 -148590
rect 36270 -148540 37390 -148530
rect 36270 -148590 36280 -148540
rect 37380 -148590 37390 -148540
rect 36270 -148600 37390 -148590
rect 37770 -148540 38890 -148530
rect 37770 -148590 37780 -148540
rect 38880 -148590 38890 -148540
rect 37770 -148600 38890 -148590
rect 39270 -148540 40390 -148530
rect 39270 -148590 39280 -148540
rect 40380 -148590 40390 -148540
rect 39270 -148600 40390 -148590
rect 40770 -148540 41890 -148530
rect 40770 -148590 40780 -148540
rect 41880 -148590 41890 -148540
rect 40770 -148600 41890 -148590
rect 42270 -148540 43390 -148530
rect 42270 -148590 42280 -148540
rect 43380 -148590 43390 -148540
rect 42270 -148600 43390 -148590
rect 43770 -148540 44890 -148530
rect 43770 -148590 43780 -148540
rect 44880 -148590 44890 -148540
rect 43770 -148600 44890 -148590
rect 45270 -148540 46390 -148530
rect 45270 -148590 45280 -148540
rect 46380 -148590 46390 -148540
rect 45270 -148600 46390 -148590
rect 46770 -148540 47890 -148530
rect 46770 -148590 46780 -148540
rect 47880 -148590 47890 -148540
rect 46770 -148600 47890 -148590
rect 48270 -148540 49390 -148530
rect 48270 -148590 48280 -148540
rect 49380 -148590 49390 -148540
rect 48270 -148600 49390 -148590
rect 49770 -148540 50890 -148530
rect 49770 -148590 49780 -148540
rect 50880 -148590 50890 -148540
rect 49770 -148600 50890 -148590
rect 51270 -148540 52390 -148530
rect 51270 -148590 51280 -148540
rect 52380 -148590 52390 -148540
rect 51270 -148600 52390 -148590
rect 52770 -148540 53890 -148530
rect 52770 -148590 52780 -148540
rect 53880 -148590 53890 -148540
rect 52770 -148600 53890 -148590
rect 54270 -148540 55390 -148530
rect 54270 -148590 54280 -148540
rect 55380 -148590 55390 -148540
rect 54270 -148600 55390 -148590
rect 55770 -148540 56890 -148530
rect 55770 -148590 55780 -148540
rect 56880 -148590 56890 -148540
rect 55770 -148600 56890 -148590
rect 57270 -148540 58390 -148530
rect 57270 -148590 57280 -148540
rect 58380 -148590 58390 -148540
rect 57270 -148600 58390 -148590
rect 58770 -148540 59890 -148530
rect 58770 -148590 58780 -148540
rect 59880 -148590 59890 -148540
rect 58770 -148600 59890 -148590
rect 60270 -148540 61390 -148530
rect 60270 -148590 60280 -148540
rect 61380 -148590 61390 -148540
rect 60270 -148600 61390 -148590
rect 61770 -148540 62890 -148530
rect 61770 -148590 61780 -148540
rect 62880 -148590 62890 -148540
rect 61770 -148600 62890 -148590
rect 63270 -148540 64390 -148530
rect 63270 -148590 63280 -148540
rect 64380 -148590 64390 -148540
rect 63270 -148600 64390 -148590
rect 64770 -148540 65890 -148530
rect 64770 -148590 64780 -148540
rect 65880 -148590 65890 -148540
rect 64770 -148600 65890 -148590
rect 66270 -148540 67390 -148530
rect 66270 -148590 66280 -148540
rect 67380 -148590 67390 -148540
rect 66270 -148600 67390 -148590
rect 67770 -148540 68890 -148530
rect 67770 -148590 67780 -148540
rect 68880 -148590 68890 -148540
rect 67770 -148600 68890 -148590
rect 69270 -148540 70390 -148530
rect 69270 -148590 69280 -148540
rect 70380 -148590 70390 -148540
rect 69270 -148600 70390 -148590
rect 70770 -148540 71890 -148530
rect 70770 -148590 70780 -148540
rect 71880 -148590 71890 -148540
rect 70770 -148600 71890 -148590
rect 72270 -148540 73390 -148530
rect 72270 -148590 72280 -148540
rect 73380 -148590 73390 -148540
rect 72270 -148600 73390 -148590
rect 73770 -148540 74890 -148530
rect 73770 -148590 73780 -148540
rect 74880 -148590 74890 -148540
rect 73770 -148600 74890 -148590
rect 75270 -148540 76390 -148530
rect 75270 -148590 75280 -148540
rect 76380 -148590 76390 -148540
rect 75270 -148600 76390 -148590
rect 76770 -148540 77890 -148530
rect 76770 -148590 76780 -148540
rect 77880 -148590 77890 -148540
rect 76770 -148600 77890 -148590
rect 78270 -148540 79390 -148530
rect 78270 -148590 78280 -148540
rect 79380 -148590 79390 -148540
rect 78270 -148600 79390 -148590
rect 79770 -148540 80890 -148530
rect 79770 -148590 79780 -148540
rect 80880 -148590 80890 -148540
rect 79770 -148600 80890 -148590
rect 81270 -148540 82390 -148530
rect 81270 -148590 81280 -148540
rect 82380 -148590 82390 -148540
rect 81270 -148600 82390 -148590
rect 82770 -148540 83890 -148530
rect 82770 -148590 82780 -148540
rect 83880 -148590 83890 -148540
rect 82770 -148600 83890 -148590
rect 84270 -148540 85390 -148530
rect 84270 -148590 84280 -148540
rect 85380 -148590 85390 -148540
rect 84270 -148600 85390 -148590
rect 85770 -148540 86890 -148530
rect 85770 -148590 85780 -148540
rect 86880 -148590 86890 -148540
rect 85770 -148600 86890 -148590
rect 87270 -148540 88390 -148530
rect 87270 -148590 87280 -148540
rect 88380 -148590 88390 -148540
rect 87270 -148600 88390 -148590
rect 88770 -148540 89890 -148530
rect 88770 -148590 88780 -148540
rect 89880 -148590 89890 -148540
rect 88770 -148600 89890 -148590
rect 90270 -148540 91390 -148530
rect 90270 -148590 90280 -148540
rect 91380 -148590 91390 -148540
rect 90270 -148600 91390 -148590
rect 91770 -148540 92890 -148530
rect 91770 -148590 91780 -148540
rect 92880 -148590 92890 -148540
rect 91770 -148600 92890 -148590
rect 93270 -148540 94390 -148530
rect 93270 -148590 93280 -148540
rect 94380 -148590 94390 -148540
rect 93270 -148600 94390 -148590
rect 94770 -148540 95890 -148530
rect 94770 -148590 94780 -148540
rect 95880 -148590 95890 -148540
rect 94770 -148600 95890 -148590
rect 96270 -148540 97390 -148530
rect 96270 -148590 96280 -148540
rect 97380 -148590 97390 -148540
rect 96270 -148600 97390 -148590
rect 97770 -148540 98890 -148530
rect 97770 -148590 97780 -148540
rect 98880 -148590 98890 -148540
rect 97770 -148600 98890 -148590
rect 99270 -148540 100390 -148530
rect 99270 -148590 99280 -148540
rect 100380 -148590 100390 -148540
rect 99270 -148600 100390 -148590
rect 100770 -148540 101890 -148530
rect 100770 -148590 100780 -148540
rect 101880 -148590 101890 -148540
rect 100770 -148600 101890 -148590
rect 102270 -148540 103390 -148530
rect 102270 -148590 102280 -148540
rect 103380 -148590 103390 -148540
rect 102270 -148600 103390 -148590
rect 103770 -148540 104890 -148530
rect 103770 -148590 103780 -148540
rect 104880 -148590 104890 -148540
rect 103770 -148600 104890 -148590
rect 105270 -148540 106390 -148530
rect 105270 -148590 105280 -148540
rect 106380 -148590 106390 -148540
rect 105270 -148600 106390 -148590
rect 106770 -148540 107890 -148530
rect 106770 -148590 106780 -148540
rect 107880 -148590 107890 -148540
rect 106770 -148600 107890 -148590
rect 108270 -148540 109390 -148530
rect 108270 -148590 108280 -148540
rect 109380 -148590 109390 -148540
rect 108270 -148600 109390 -148590
rect 109770 -148540 110890 -148530
rect 109770 -148590 109780 -148540
rect 110880 -148590 110890 -148540
rect 109770 -148600 110890 -148590
rect 111270 -148540 112390 -148530
rect 111270 -148590 111280 -148540
rect 112380 -148590 112390 -148540
rect 111270 -148600 112390 -148590
rect 112770 -148540 113890 -148530
rect 112770 -148590 112780 -148540
rect 113880 -148590 113890 -148540
rect 112770 -148600 113890 -148590
rect 114270 -148540 115390 -148530
rect 114270 -148590 114280 -148540
rect 115380 -148590 115390 -148540
rect 114270 -148600 115390 -148590
rect 115770 -148540 116890 -148530
rect 115770 -148590 115780 -148540
rect 116880 -148590 116890 -148540
rect 115770 -148600 116890 -148590
rect 117270 -148540 118390 -148530
rect 117270 -148590 117280 -148540
rect 118380 -148590 118390 -148540
rect 117270 -148600 118390 -148590
rect 118770 -148540 119890 -148530
rect 118770 -148590 118780 -148540
rect 119880 -148590 119890 -148540
rect 118770 -148600 119890 -148590
rect 120270 -148540 121390 -148530
rect 120270 -148590 120280 -148540
rect 121380 -148590 121390 -148540
rect 120270 -148600 121390 -148590
rect 121770 -148540 122890 -148530
rect 121770 -148590 121780 -148540
rect 122880 -148590 122890 -148540
rect 121770 -148600 122890 -148590
rect 123270 -148540 124390 -148530
rect 123270 -148590 123280 -148540
rect 124380 -148590 124390 -148540
rect 123270 -148600 124390 -148590
rect 124770 -148540 125890 -148530
rect 124770 -148590 124780 -148540
rect 125880 -148590 125890 -148540
rect 124770 -148600 125890 -148590
rect 126270 -148540 127390 -148530
rect 126270 -148590 126280 -148540
rect 127380 -148590 127390 -148540
rect 126270 -148600 127390 -148590
rect 127770 -148540 128890 -148530
rect 127770 -148590 127780 -148540
rect 128880 -148590 128890 -148540
rect 127770 -148600 128890 -148590
rect 129270 -148540 130390 -148530
rect 129270 -148590 129280 -148540
rect 130380 -148590 130390 -148540
rect 129270 -148600 130390 -148590
rect 130770 -148540 131890 -148530
rect 130770 -148590 130780 -148540
rect 131880 -148590 131890 -148540
rect 130770 -148600 131890 -148590
rect 132270 -148540 133390 -148530
rect 132270 -148590 132280 -148540
rect 133380 -148590 133390 -148540
rect 132270 -148600 133390 -148590
rect 133770 -148540 134890 -148530
rect 133770 -148590 133780 -148540
rect 134880 -148590 134890 -148540
rect 133770 -148600 134890 -148590
rect 135270 -148540 136390 -148530
rect 135270 -148590 135280 -148540
rect 136380 -148590 136390 -148540
rect 135270 -148600 136390 -148590
rect 136770 -148540 137890 -148530
rect 136770 -148590 136780 -148540
rect 137880 -148590 137890 -148540
rect 136770 -148600 137890 -148590
rect 138270 -148540 139390 -148530
rect 138270 -148590 138280 -148540
rect 139380 -148590 139390 -148540
rect 138270 -148600 139390 -148590
rect 139770 -148540 140890 -148530
rect 139770 -148590 139780 -148540
rect 140880 -148590 140890 -148540
rect 139770 -148600 140890 -148590
rect 141270 -148540 142390 -148530
rect 141270 -148590 141280 -148540
rect 142380 -148590 142390 -148540
rect 141270 -148600 142390 -148590
rect 142770 -148540 143890 -148530
rect 142770 -148590 142780 -148540
rect 143880 -148590 143890 -148540
rect 142770 -148600 143890 -148590
rect 144270 -148540 145390 -148530
rect 144270 -148590 144280 -148540
rect 145380 -148590 145390 -148540
rect 144270 -148600 145390 -148590
rect 145770 -148540 146890 -148530
rect 145770 -148590 145780 -148540
rect 146880 -148590 146890 -148540
rect 145770 -148600 146890 -148590
rect 147270 -148540 148390 -148530
rect 147270 -148590 147280 -148540
rect 148380 -148590 148390 -148540
rect 147270 -148600 148390 -148590
rect 148770 -148540 149890 -148530
rect 148770 -148590 148780 -148540
rect 149880 -148590 149890 -148540
rect 148770 -148600 149890 -148590
rect 110 -148750 220 -148745
rect 110 -148850 120 -148750
rect 210 -148850 220 -148750
rect 110 -149050 220 -148850
rect 1610 -148750 1720 -148745
rect 1610 -148850 1620 -148750
rect 1710 -148850 1720 -148750
rect 1610 -149050 1720 -148850
rect 3110 -148750 3220 -148745
rect 3110 -148850 3120 -148750
rect 3210 -148850 3220 -148750
rect 3110 -149050 3220 -148850
rect 4610 -148750 4720 -148745
rect 4610 -148850 4620 -148750
rect 4710 -148850 4720 -148750
rect 4610 -149050 4720 -148850
rect 6110 -148750 6220 -148745
rect 6110 -148850 6120 -148750
rect 6210 -148850 6220 -148750
rect 6110 -149050 6220 -148850
rect 7610 -148750 7720 -148745
rect 7610 -148850 7620 -148750
rect 7710 -148850 7720 -148750
rect 7610 -149050 7720 -148850
rect 9110 -148750 9220 -148745
rect 9110 -148850 9120 -148750
rect 9210 -148850 9220 -148750
rect 9110 -149050 9220 -148850
rect 10610 -148750 10720 -148745
rect 10610 -148850 10620 -148750
rect 10710 -148850 10720 -148750
rect 10610 -149050 10720 -148850
rect 12110 -148750 12220 -148745
rect 12110 -148850 12120 -148750
rect 12210 -148850 12220 -148750
rect 12110 -149050 12220 -148850
rect 13610 -148750 13720 -148745
rect 13610 -148850 13620 -148750
rect 13710 -148850 13720 -148750
rect 13610 -149050 13720 -148850
rect 15110 -148750 15220 -148745
rect 15110 -148850 15120 -148750
rect 15210 -148850 15220 -148750
rect 15110 -149050 15220 -148850
rect 16610 -148750 16720 -148745
rect 16610 -148850 16620 -148750
rect 16710 -148850 16720 -148750
rect 16610 -149050 16720 -148850
rect 18110 -148750 18220 -148745
rect 18110 -148850 18120 -148750
rect 18210 -148850 18220 -148750
rect 18110 -149050 18220 -148850
rect 19610 -148750 19720 -148745
rect 19610 -148850 19620 -148750
rect 19710 -148850 19720 -148750
rect 19610 -149050 19720 -148850
rect 21110 -148750 21220 -148745
rect 21110 -148850 21120 -148750
rect 21210 -148850 21220 -148750
rect 21110 -149050 21220 -148850
rect 22610 -148750 22720 -148745
rect 22610 -148850 22620 -148750
rect 22710 -148850 22720 -148750
rect 22610 -149050 22720 -148850
rect 24110 -148750 24220 -148745
rect 24110 -148850 24120 -148750
rect 24210 -148850 24220 -148750
rect 24110 -149050 24220 -148850
rect 25610 -148750 25720 -148745
rect 25610 -148850 25620 -148750
rect 25710 -148850 25720 -148750
rect 25610 -149050 25720 -148850
rect 27110 -148750 27220 -148745
rect 27110 -148850 27120 -148750
rect 27210 -148850 27220 -148750
rect 27110 -149050 27220 -148850
rect 28610 -148750 28720 -148745
rect 28610 -148850 28620 -148750
rect 28710 -148850 28720 -148750
rect 28610 -149050 28720 -148850
rect 30110 -148750 30220 -148745
rect 30110 -148850 30120 -148750
rect 30210 -148850 30220 -148750
rect 30110 -149050 30220 -148850
rect 31610 -148750 31720 -148745
rect 31610 -148850 31620 -148750
rect 31710 -148850 31720 -148750
rect 31610 -149050 31720 -148850
rect 33110 -148750 33220 -148745
rect 33110 -148850 33120 -148750
rect 33210 -148850 33220 -148750
rect 33110 -149050 33220 -148850
rect 34610 -148750 34720 -148745
rect 34610 -148850 34620 -148750
rect 34710 -148850 34720 -148750
rect 34610 -149050 34720 -148850
rect 36110 -148750 36220 -148745
rect 36110 -148850 36120 -148750
rect 36210 -148850 36220 -148750
rect 36110 -149050 36220 -148850
rect 37610 -148750 37720 -148745
rect 37610 -148850 37620 -148750
rect 37710 -148850 37720 -148750
rect 37610 -149050 37720 -148850
rect 39110 -148750 39220 -148745
rect 39110 -148850 39120 -148750
rect 39210 -148850 39220 -148750
rect 39110 -149050 39220 -148850
rect 40610 -148750 40720 -148745
rect 40610 -148850 40620 -148750
rect 40710 -148850 40720 -148750
rect 40610 -149050 40720 -148850
rect 42110 -148750 42220 -148745
rect 42110 -148850 42120 -148750
rect 42210 -148850 42220 -148750
rect 42110 -149050 42220 -148850
rect 43610 -148750 43720 -148745
rect 43610 -148850 43620 -148750
rect 43710 -148850 43720 -148750
rect 43610 -149050 43720 -148850
rect 45110 -148750 45220 -148745
rect 45110 -148850 45120 -148750
rect 45210 -148850 45220 -148750
rect 45110 -149050 45220 -148850
rect 46610 -148750 46720 -148745
rect 46610 -148850 46620 -148750
rect 46710 -148850 46720 -148750
rect 46610 -149050 46720 -148850
rect 48110 -148750 48220 -148745
rect 48110 -148850 48120 -148750
rect 48210 -148850 48220 -148750
rect 48110 -149050 48220 -148850
rect 49610 -148750 49720 -148745
rect 49610 -148850 49620 -148750
rect 49710 -148850 49720 -148750
rect 49610 -149050 49720 -148850
rect 51110 -148750 51220 -148745
rect 51110 -148850 51120 -148750
rect 51210 -148850 51220 -148750
rect 51110 -149050 51220 -148850
rect 52610 -148750 52720 -148745
rect 52610 -148850 52620 -148750
rect 52710 -148850 52720 -148750
rect 52610 -149050 52720 -148850
rect 54110 -148750 54220 -148745
rect 54110 -148850 54120 -148750
rect 54210 -148850 54220 -148750
rect 54110 -149050 54220 -148850
rect 55610 -148750 55720 -148745
rect 55610 -148850 55620 -148750
rect 55710 -148850 55720 -148750
rect 55610 -149050 55720 -148850
rect 57110 -148750 57220 -148745
rect 57110 -148850 57120 -148750
rect 57210 -148850 57220 -148750
rect 57110 -149050 57220 -148850
rect 58610 -148750 58720 -148745
rect 58610 -148850 58620 -148750
rect 58710 -148850 58720 -148750
rect 58610 -149050 58720 -148850
rect 60110 -148750 60220 -148745
rect 60110 -148850 60120 -148750
rect 60210 -148850 60220 -148750
rect 60110 -149050 60220 -148850
rect 61610 -148750 61720 -148745
rect 61610 -148850 61620 -148750
rect 61710 -148850 61720 -148750
rect 61610 -149050 61720 -148850
rect 63110 -148750 63220 -148745
rect 63110 -148850 63120 -148750
rect 63210 -148850 63220 -148750
rect 63110 -149050 63220 -148850
rect 64610 -148750 64720 -148745
rect 64610 -148850 64620 -148750
rect 64710 -148850 64720 -148750
rect 64610 -149050 64720 -148850
rect 66110 -148750 66220 -148745
rect 66110 -148850 66120 -148750
rect 66210 -148850 66220 -148750
rect 66110 -149050 66220 -148850
rect 67610 -148750 67720 -148745
rect 67610 -148850 67620 -148750
rect 67710 -148850 67720 -148750
rect 67610 -149050 67720 -148850
rect 69110 -148750 69220 -148745
rect 69110 -148850 69120 -148750
rect 69210 -148850 69220 -148750
rect 69110 -149050 69220 -148850
rect 70610 -148750 70720 -148745
rect 70610 -148850 70620 -148750
rect 70710 -148850 70720 -148750
rect 70610 -149050 70720 -148850
rect 72110 -148750 72220 -148745
rect 72110 -148850 72120 -148750
rect 72210 -148850 72220 -148750
rect 72110 -149050 72220 -148850
rect 73610 -148750 73720 -148745
rect 73610 -148850 73620 -148750
rect 73710 -148850 73720 -148750
rect 73610 -149050 73720 -148850
rect 75110 -148750 75220 -148745
rect 75110 -148850 75120 -148750
rect 75210 -148850 75220 -148750
rect 75110 -149050 75220 -148850
rect 76610 -148750 76720 -148745
rect 76610 -148850 76620 -148750
rect 76710 -148850 76720 -148750
rect 76610 -149050 76720 -148850
rect 78110 -148750 78220 -148745
rect 78110 -148850 78120 -148750
rect 78210 -148850 78220 -148750
rect 78110 -149050 78220 -148850
rect 79610 -148750 79720 -148745
rect 79610 -148850 79620 -148750
rect 79710 -148850 79720 -148750
rect 79610 -149050 79720 -148850
rect 81110 -148750 81220 -148745
rect 81110 -148850 81120 -148750
rect 81210 -148850 81220 -148750
rect 81110 -149050 81220 -148850
rect 82610 -148750 82720 -148745
rect 82610 -148850 82620 -148750
rect 82710 -148850 82720 -148750
rect 82610 -149050 82720 -148850
rect 84110 -148750 84220 -148745
rect 84110 -148850 84120 -148750
rect 84210 -148850 84220 -148750
rect 84110 -149050 84220 -148850
rect 85610 -148750 85720 -148745
rect 85610 -148850 85620 -148750
rect 85710 -148850 85720 -148750
rect 85610 -149050 85720 -148850
rect 87110 -148750 87220 -148745
rect 87110 -148850 87120 -148750
rect 87210 -148850 87220 -148750
rect 87110 -149050 87220 -148850
rect 88610 -148750 88720 -148745
rect 88610 -148850 88620 -148750
rect 88710 -148850 88720 -148750
rect 88610 -149050 88720 -148850
rect 90110 -148750 90220 -148745
rect 90110 -148850 90120 -148750
rect 90210 -148850 90220 -148750
rect 90110 -149050 90220 -148850
rect 91610 -148750 91720 -148745
rect 91610 -148850 91620 -148750
rect 91710 -148850 91720 -148750
rect 91610 -149050 91720 -148850
rect 93110 -148750 93220 -148745
rect 93110 -148850 93120 -148750
rect 93210 -148850 93220 -148750
rect 93110 -149050 93220 -148850
rect 94610 -148750 94720 -148745
rect 94610 -148850 94620 -148750
rect 94710 -148850 94720 -148750
rect 94610 -149050 94720 -148850
rect 96110 -148750 96220 -148745
rect 96110 -148850 96120 -148750
rect 96210 -148850 96220 -148750
rect 96110 -149050 96220 -148850
rect 97610 -148750 97720 -148745
rect 97610 -148850 97620 -148750
rect 97710 -148850 97720 -148750
rect 97610 -149050 97720 -148850
rect 99110 -148750 99220 -148745
rect 99110 -148850 99120 -148750
rect 99210 -148850 99220 -148750
rect 99110 -149050 99220 -148850
rect 100610 -148750 100720 -148745
rect 100610 -148850 100620 -148750
rect 100710 -148850 100720 -148750
rect 100610 -149050 100720 -148850
rect 102110 -148750 102220 -148745
rect 102110 -148850 102120 -148750
rect 102210 -148850 102220 -148750
rect 102110 -149050 102220 -148850
rect 103610 -148750 103720 -148745
rect 103610 -148850 103620 -148750
rect 103710 -148850 103720 -148750
rect 103610 -149050 103720 -148850
rect 105110 -148750 105220 -148745
rect 105110 -148850 105120 -148750
rect 105210 -148850 105220 -148750
rect 105110 -149050 105220 -148850
rect 106610 -148750 106720 -148745
rect 106610 -148850 106620 -148750
rect 106710 -148850 106720 -148750
rect 106610 -149050 106720 -148850
rect 108110 -148750 108220 -148745
rect 108110 -148850 108120 -148750
rect 108210 -148850 108220 -148750
rect 108110 -149050 108220 -148850
rect 109610 -148750 109720 -148745
rect 109610 -148850 109620 -148750
rect 109710 -148850 109720 -148750
rect 109610 -149050 109720 -148850
rect 111110 -148750 111220 -148745
rect 111110 -148850 111120 -148750
rect 111210 -148850 111220 -148750
rect 111110 -149050 111220 -148850
rect 112610 -148750 112720 -148745
rect 112610 -148850 112620 -148750
rect 112710 -148850 112720 -148750
rect 112610 -149050 112720 -148850
rect 114110 -148750 114220 -148745
rect 114110 -148850 114120 -148750
rect 114210 -148850 114220 -148750
rect 114110 -149050 114220 -148850
rect 115610 -148750 115720 -148745
rect 115610 -148850 115620 -148750
rect 115710 -148850 115720 -148750
rect 115610 -149050 115720 -148850
rect 117110 -148750 117220 -148745
rect 117110 -148850 117120 -148750
rect 117210 -148850 117220 -148750
rect 117110 -149050 117220 -148850
rect 118610 -148750 118720 -148745
rect 118610 -148850 118620 -148750
rect 118710 -148850 118720 -148750
rect 118610 -149050 118720 -148850
rect 120110 -148750 120220 -148745
rect 120110 -148850 120120 -148750
rect 120210 -148850 120220 -148750
rect 120110 -149050 120220 -148850
rect 121610 -148750 121720 -148745
rect 121610 -148850 121620 -148750
rect 121710 -148850 121720 -148750
rect 121610 -149050 121720 -148850
rect 123110 -148750 123220 -148745
rect 123110 -148850 123120 -148750
rect 123210 -148850 123220 -148750
rect 123110 -149050 123220 -148850
rect 124610 -148750 124720 -148745
rect 124610 -148850 124620 -148750
rect 124710 -148850 124720 -148750
rect 124610 -149050 124720 -148850
rect 126110 -148750 126220 -148745
rect 126110 -148850 126120 -148750
rect 126210 -148850 126220 -148750
rect 126110 -149050 126220 -148850
rect 127610 -148750 127720 -148745
rect 127610 -148850 127620 -148750
rect 127710 -148850 127720 -148750
rect 127610 -149050 127720 -148850
rect 129110 -148750 129220 -148745
rect 129110 -148850 129120 -148750
rect 129210 -148850 129220 -148750
rect 129110 -149050 129220 -148850
rect 130610 -148750 130720 -148745
rect 130610 -148850 130620 -148750
rect 130710 -148850 130720 -148750
rect 130610 -149050 130720 -148850
rect 132110 -148750 132220 -148745
rect 132110 -148850 132120 -148750
rect 132210 -148850 132220 -148750
rect 132110 -149050 132220 -148850
rect 133610 -148750 133720 -148745
rect 133610 -148850 133620 -148750
rect 133710 -148850 133720 -148750
rect 133610 -149050 133720 -148850
rect 135110 -148750 135220 -148745
rect 135110 -148850 135120 -148750
rect 135210 -148850 135220 -148750
rect 135110 -149050 135220 -148850
rect 136610 -148750 136720 -148745
rect 136610 -148850 136620 -148750
rect 136710 -148850 136720 -148750
rect 136610 -149050 136720 -148850
rect 138110 -148750 138220 -148745
rect 138110 -148850 138120 -148750
rect 138210 -148850 138220 -148750
rect 138110 -149050 138220 -148850
rect 139610 -148750 139720 -148745
rect 139610 -148850 139620 -148750
rect 139710 -148850 139720 -148750
rect 139610 -149050 139720 -148850
rect 141110 -148750 141220 -148745
rect 141110 -148850 141120 -148750
rect 141210 -148850 141220 -148750
rect 141110 -149050 141220 -148850
rect 142610 -148750 142720 -148745
rect 142610 -148850 142620 -148750
rect 142710 -148850 142720 -148750
rect 142610 -149050 142720 -148850
rect 144110 -148750 144220 -148745
rect 144110 -148850 144120 -148750
rect 144210 -148850 144220 -148750
rect 144110 -149050 144220 -148850
rect 145610 -148750 145720 -148745
rect 145610 -148850 145620 -148750
rect 145710 -148850 145720 -148750
rect 145610 -149050 145720 -148850
rect 147110 -148750 147220 -148745
rect 147110 -148850 147120 -148750
rect 147210 -148850 147220 -148750
rect 147110 -149050 147220 -148850
rect 148610 -148750 148720 -148745
rect 148610 -148850 148620 -148750
rect 148710 -148850 148720 -148750
rect 148610 -149050 148720 -148850
<< metal5 >>
rect -1000 1420 0 1580
use pixel  pixel_0
timestamp 1757982896
transform 1 0 -1900 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_1
timestamp 1757982896
transform 1 0 -400 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_2
timestamp 1757982896
transform 1 0 1100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_3
timestamp 1757982896
transform 1 0 2600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_4
timestamp 1757982896
transform 1 0 4100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_5
timestamp 1757982896
transform 1 0 5600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_6
timestamp 1757982896
transform 1 0 7100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_7
timestamp 1757982896
transform 1 0 8600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_8
timestamp 1757982896
transform 1 0 10100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_9
timestamp 1757982896
transform 1 0 11600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_10
timestamp 1757982896
transform 1 0 13100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_11
timestamp 1757982896
transform 1 0 14600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_12
timestamp 1757982896
transform 1 0 16100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_13
timestamp 1757982896
transform 1 0 17600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_14
timestamp 1757982896
transform 1 0 19100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_15
timestamp 1757982896
transform 1 0 20600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_16
timestamp 1757982896
transform 1 0 22100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_17
timestamp 1757982896
transform 1 0 23600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_18
timestamp 1757982896
transform 1 0 25100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_19
timestamp 1757982896
transform 1 0 26600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_20
timestamp 1757982896
transform 1 0 28100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_21
timestamp 1757982896
transform 1 0 29600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_22
timestamp 1757982896
transform 1 0 31100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_23
timestamp 1757982896
transform 1 0 32600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_24
timestamp 1757982896
transform 1 0 34100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_25
timestamp 1757982896
transform 1 0 35600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_26
timestamp 1757982896
transform 1 0 37100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_27
timestamp 1757982896
transform 1 0 38600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_28
timestamp 1757982896
transform 1 0 40100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_29
timestamp 1757982896
transform 1 0 41600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_30
timestamp 1757982896
transform 1 0 43100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_31
timestamp 1757982896
transform 1 0 44600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_32
timestamp 1757982896
transform 1 0 46100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_33
timestamp 1757982896
transform 1 0 47600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_34
timestamp 1757982896
transform 1 0 49100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_35
timestamp 1757982896
transform 1 0 50600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_36
timestamp 1757982896
transform 1 0 52100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_37
timestamp 1757982896
transform 1 0 53600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_38
timestamp 1757982896
transform 1 0 55100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_39
timestamp 1757982896
transform 1 0 56600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_40
timestamp 1757982896
transform 1 0 58100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_41
timestamp 1757982896
transform 1 0 59600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_42
timestamp 1757982896
transform 1 0 61100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_43
timestamp 1757982896
transform 1 0 62600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_44
timestamp 1757982896
transform 1 0 64100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_45
timestamp 1757982896
transform 1 0 65600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_46
timestamp 1757982896
transform 1 0 67100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_47
timestamp 1757982896
transform 1 0 68600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_48
timestamp 1757982896
transform 1 0 70100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_49
timestamp 1757982896
transform 1 0 71600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_50
timestamp 1757982896
transform 1 0 73100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_51
timestamp 1757982896
transform 1 0 74600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_52
timestamp 1757982896
transform 1 0 76100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_53
timestamp 1757982896
transform 1 0 77600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_54
timestamp 1757982896
transform 1 0 79100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_55
timestamp 1757982896
transform 1 0 80600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_56
timestamp 1757982896
transform 1 0 82100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_57
timestamp 1757982896
transform 1 0 83600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_58
timestamp 1757982896
transform 1 0 85100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_59
timestamp 1757982896
transform 1 0 86600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_60
timestamp 1757982896
transform 1 0 88100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_61
timestamp 1757982896
transform 1 0 89600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_62
timestamp 1757982896
transform 1 0 91100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_63
timestamp 1757982896
transform 1 0 92600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_64
timestamp 1757982896
transform 1 0 94100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_65
timestamp 1757982896
transform 1 0 95600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_66
timestamp 1757982896
transform 1 0 97100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_67
timestamp 1757982896
transform 1 0 98600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_68
timestamp 1757982896
transform 1 0 100100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_69
timestamp 1757982896
transform 1 0 101600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_70
timestamp 1757982896
transform 1 0 103100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_71
timestamp 1757982896
transform 1 0 104600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_72
timestamp 1757982896
transform 1 0 106100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_73
timestamp 1757982896
transform 1 0 107600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_74
timestamp 1757982896
transform 1 0 109100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_75
timestamp 1757982896
transform 1 0 110600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_76
timestamp 1757982896
transform 1 0 112100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_77
timestamp 1757982896
transform 1 0 113600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_78
timestamp 1757982896
transform 1 0 115100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_79
timestamp 1757982896
transform 1 0 116600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_80
timestamp 1757982896
transform 1 0 118100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_81
timestamp 1757982896
transform 1 0 119600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_82
timestamp 1757982896
transform 1 0 121100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_83
timestamp 1757982896
transform 1 0 122600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_84
timestamp 1757982896
transform 1 0 124100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_85
timestamp 1757982896
transform 1 0 125600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_86
timestamp 1757982896
transform 1 0 127100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_87
timestamp 1757982896
transform 1 0 128600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_88
timestamp 1757982896
transform 1 0 130100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_89
timestamp 1757982896
transform 1 0 131600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_90
timestamp 1757982896
transform 1 0 133100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_91
timestamp 1757982896
transform 1 0 134600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_92
timestamp 1757982896
transform 1 0 136100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_93
timestamp 1757982896
transform 1 0 137600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_94
timestamp 1757982896
transform 1 0 139100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_95
timestamp 1757982896
transform 1 0 140600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_96
timestamp 1757982896
transform 1 0 142100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_97
timestamp 1757982896
transform 1 0 143600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_98
timestamp 1757982896
transform 1 0 145100 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_99
timestamp 1757982896
transform 1 0 146600 0 1 1350
box 1820 -1430 3480 230
use pixel  pixel_100
timestamp 1757982896
transform 1 0 -1900 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_101
timestamp 1757982896
transform 1 0 -400 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_102
timestamp 1757982896
transform 1 0 1100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_103
timestamp 1757982896
transform 1 0 2600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_104
timestamp 1757982896
transform 1 0 4100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_105
timestamp 1757982896
transform 1 0 5600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_106
timestamp 1757982896
transform 1 0 7100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_107
timestamp 1757982896
transform 1 0 8600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_108
timestamp 1757982896
transform 1 0 10100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_109
timestamp 1757982896
transform 1 0 11600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_110
timestamp 1757982896
transform 1 0 13100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_111
timestamp 1757982896
transform 1 0 14600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_112
timestamp 1757982896
transform 1 0 16100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_113
timestamp 1757982896
transform 1 0 17600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_114
timestamp 1757982896
transform 1 0 19100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_115
timestamp 1757982896
transform 1 0 20600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_116
timestamp 1757982896
transform 1 0 22100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_117
timestamp 1757982896
transform 1 0 23600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_118
timestamp 1757982896
transform 1 0 25100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_119
timestamp 1757982896
transform 1 0 26600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_120
timestamp 1757982896
transform 1 0 28100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_121
timestamp 1757982896
transform 1 0 29600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_122
timestamp 1757982896
transform 1 0 31100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_123
timestamp 1757982896
transform 1 0 32600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_124
timestamp 1757982896
transform 1 0 34100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_125
timestamp 1757982896
transform 1 0 35600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_126
timestamp 1757982896
transform 1 0 37100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_127
timestamp 1757982896
transform 1 0 38600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_128
timestamp 1757982896
transform 1 0 40100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_129
timestamp 1757982896
transform 1 0 41600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_130
timestamp 1757982896
transform 1 0 43100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_131
timestamp 1757982896
transform 1 0 44600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_132
timestamp 1757982896
transform 1 0 46100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_133
timestamp 1757982896
transform 1 0 47600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_134
timestamp 1757982896
transform 1 0 49100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_135
timestamp 1757982896
transform 1 0 50600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_136
timestamp 1757982896
transform 1 0 52100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_137
timestamp 1757982896
transform 1 0 53600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_138
timestamp 1757982896
transform 1 0 55100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_139
timestamp 1757982896
transform 1 0 56600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_140
timestamp 1757982896
transform 1 0 58100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_141
timestamp 1757982896
transform 1 0 59600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_142
timestamp 1757982896
transform 1 0 61100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_143
timestamp 1757982896
transform 1 0 62600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_144
timestamp 1757982896
transform 1 0 64100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_145
timestamp 1757982896
transform 1 0 65600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_146
timestamp 1757982896
transform 1 0 67100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_147
timestamp 1757982896
transform 1 0 68600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_148
timestamp 1757982896
transform 1 0 70100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_149
timestamp 1757982896
transform 1 0 71600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_150
timestamp 1757982896
transform 1 0 73100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_151
timestamp 1757982896
transform 1 0 74600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_152
timestamp 1757982896
transform 1 0 76100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_153
timestamp 1757982896
transform 1 0 77600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_154
timestamp 1757982896
transform 1 0 79100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_155
timestamp 1757982896
transform 1 0 80600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_156
timestamp 1757982896
transform 1 0 82100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_157
timestamp 1757982896
transform 1 0 83600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_158
timestamp 1757982896
transform 1 0 85100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_159
timestamp 1757982896
transform 1 0 86600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_160
timestamp 1757982896
transform 1 0 88100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_161
timestamp 1757982896
transform 1 0 89600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_162
timestamp 1757982896
transform 1 0 91100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_163
timestamp 1757982896
transform 1 0 92600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_164
timestamp 1757982896
transform 1 0 94100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_165
timestamp 1757982896
transform 1 0 95600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_166
timestamp 1757982896
transform 1 0 97100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_167
timestamp 1757982896
transform 1 0 98600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_168
timestamp 1757982896
transform 1 0 100100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_169
timestamp 1757982896
transform 1 0 101600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_170
timestamp 1757982896
transform 1 0 103100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_171
timestamp 1757982896
transform 1 0 104600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_172
timestamp 1757982896
transform 1 0 106100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_173
timestamp 1757982896
transform 1 0 107600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_174
timestamp 1757982896
transform 1 0 109100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_175
timestamp 1757982896
transform 1 0 110600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_176
timestamp 1757982896
transform 1 0 112100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_177
timestamp 1757982896
transform 1 0 113600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_178
timestamp 1757982896
transform 1 0 115100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_179
timestamp 1757982896
transform 1 0 116600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_180
timestamp 1757982896
transform 1 0 118100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_181
timestamp 1757982896
transform 1 0 119600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_182
timestamp 1757982896
transform 1 0 121100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_183
timestamp 1757982896
transform 1 0 122600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_184
timestamp 1757982896
transform 1 0 124100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_185
timestamp 1757982896
transform 1 0 125600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_186
timestamp 1757982896
transform 1 0 127100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_187
timestamp 1757982896
transform 1 0 128600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_188
timestamp 1757982896
transform 1 0 130100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_189
timestamp 1757982896
transform 1 0 131600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_190
timestamp 1757982896
transform 1 0 133100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_191
timestamp 1757982896
transform 1 0 134600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_192
timestamp 1757982896
transform 1 0 136100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_193
timestamp 1757982896
transform 1 0 137600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_194
timestamp 1757982896
transform 1 0 139100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_195
timestamp 1757982896
transform 1 0 140600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_196
timestamp 1757982896
transform 1 0 142100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_197
timestamp 1757982896
transform 1 0 143600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_198
timestamp 1757982896
transform 1 0 145100 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_199
timestamp 1757982896
transform 1 0 146600 0 1 -150
box 1820 -1430 3480 230
use pixel  pixel_200
timestamp 1757982896
transform 1 0 -1900 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_201
timestamp 1757982896
transform 1 0 -400 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_202
timestamp 1757982896
transform 1 0 1100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_203
timestamp 1757982896
transform 1 0 2600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_204
timestamp 1757982896
transform 1 0 4100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_205
timestamp 1757982896
transform 1 0 5600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_206
timestamp 1757982896
transform 1 0 7100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_207
timestamp 1757982896
transform 1 0 8600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_208
timestamp 1757982896
transform 1 0 10100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_209
timestamp 1757982896
transform 1 0 11600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_210
timestamp 1757982896
transform 1 0 13100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_211
timestamp 1757982896
transform 1 0 14600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_212
timestamp 1757982896
transform 1 0 16100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_213
timestamp 1757982896
transform 1 0 17600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_214
timestamp 1757982896
transform 1 0 19100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_215
timestamp 1757982896
transform 1 0 20600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_216
timestamp 1757982896
transform 1 0 22100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_217
timestamp 1757982896
transform 1 0 23600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_218
timestamp 1757982896
transform 1 0 25100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_219
timestamp 1757982896
transform 1 0 26600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_220
timestamp 1757982896
transform 1 0 28100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_221
timestamp 1757982896
transform 1 0 29600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_222
timestamp 1757982896
transform 1 0 31100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_223
timestamp 1757982896
transform 1 0 32600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_224
timestamp 1757982896
transform 1 0 34100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_225
timestamp 1757982896
transform 1 0 35600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_226
timestamp 1757982896
transform 1 0 37100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_227
timestamp 1757982896
transform 1 0 38600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_228
timestamp 1757982896
transform 1 0 40100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_229
timestamp 1757982896
transform 1 0 41600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_230
timestamp 1757982896
transform 1 0 43100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_231
timestamp 1757982896
transform 1 0 44600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_232
timestamp 1757982896
transform 1 0 46100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_233
timestamp 1757982896
transform 1 0 47600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_234
timestamp 1757982896
transform 1 0 49100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_235
timestamp 1757982896
transform 1 0 50600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_236
timestamp 1757982896
transform 1 0 52100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_237
timestamp 1757982896
transform 1 0 53600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_238
timestamp 1757982896
transform 1 0 55100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_239
timestamp 1757982896
transform 1 0 56600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_240
timestamp 1757982896
transform 1 0 58100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_241
timestamp 1757982896
transform 1 0 59600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_242
timestamp 1757982896
transform 1 0 61100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_243
timestamp 1757982896
transform 1 0 62600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_244
timestamp 1757982896
transform 1 0 64100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_245
timestamp 1757982896
transform 1 0 65600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_246
timestamp 1757982896
transform 1 0 67100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_247
timestamp 1757982896
transform 1 0 68600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_248
timestamp 1757982896
transform 1 0 70100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_249
timestamp 1757982896
transform 1 0 71600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_250
timestamp 1757982896
transform 1 0 73100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_251
timestamp 1757982896
transform 1 0 74600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_252
timestamp 1757982896
transform 1 0 76100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_253
timestamp 1757982896
transform 1 0 77600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_254
timestamp 1757982896
transform 1 0 79100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_255
timestamp 1757982896
transform 1 0 80600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_256
timestamp 1757982896
transform 1 0 82100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_257
timestamp 1757982896
transform 1 0 83600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_258
timestamp 1757982896
transform 1 0 85100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_259
timestamp 1757982896
transform 1 0 86600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_260
timestamp 1757982896
transform 1 0 88100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_261
timestamp 1757982896
transform 1 0 89600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_262
timestamp 1757982896
transform 1 0 91100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_263
timestamp 1757982896
transform 1 0 92600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_264
timestamp 1757982896
transform 1 0 94100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_265
timestamp 1757982896
transform 1 0 95600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_266
timestamp 1757982896
transform 1 0 97100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_267
timestamp 1757982896
transform 1 0 98600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_268
timestamp 1757982896
transform 1 0 100100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_269
timestamp 1757982896
transform 1 0 101600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_270
timestamp 1757982896
transform 1 0 103100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_271
timestamp 1757982896
transform 1 0 104600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_272
timestamp 1757982896
transform 1 0 106100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_273
timestamp 1757982896
transform 1 0 107600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_274
timestamp 1757982896
transform 1 0 109100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_275
timestamp 1757982896
transform 1 0 110600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_276
timestamp 1757982896
transform 1 0 112100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_277
timestamp 1757982896
transform 1 0 113600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_278
timestamp 1757982896
transform 1 0 115100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_279
timestamp 1757982896
transform 1 0 116600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_280
timestamp 1757982896
transform 1 0 118100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_281
timestamp 1757982896
transform 1 0 119600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_282
timestamp 1757982896
transform 1 0 121100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_283
timestamp 1757982896
transform 1 0 122600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_284
timestamp 1757982896
transform 1 0 124100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_285
timestamp 1757982896
transform 1 0 125600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_286
timestamp 1757982896
transform 1 0 127100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_287
timestamp 1757982896
transform 1 0 128600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_288
timestamp 1757982896
transform 1 0 130100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_289
timestamp 1757982896
transform 1 0 131600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_290
timestamp 1757982896
transform 1 0 133100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_291
timestamp 1757982896
transform 1 0 134600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_292
timestamp 1757982896
transform 1 0 136100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_293
timestamp 1757982896
transform 1 0 137600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_294
timestamp 1757982896
transform 1 0 139100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_295
timestamp 1757982896
transform 1 0 140600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_296
timestamp 1757982896
transform 1 0 142100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_297
timestamp 1757982896
transform 1 0 143600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_298
timestamp 1757982896
transform 1 0 145100 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_299
timestamp 1757982896
transform 1 0 146600 0 1 -1650
box 1820 -1430 3480 230
use pixel  pixel_300
timestamp 1757982896
transform 1 0 -1900 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_301
timestamp 1757982896
transform 1 0 -400 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_302
timestamp 1757982896
transform 1 0 1100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_303
timestamp 1757982896
transform 1 0 2600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_304
timestamp 1757982896
transform 1 0 4100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_305
timestamp 1757982896
transform 1 0 5600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_306
timestamp 1757982896
transform 1 0 7100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_307
timestamp 1757982896
transform 1 0 8600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_308
timestamp 1757982896
transform 1 0 10100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_309
timestamp 1757982896
transform 1 0 11600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_310
timestamp 1757982896
transform 1 0 13100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_311
timestamp 1757982896
transform 1 0 14600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_312
timestamp 1757982896
transform 1 0 16100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_313
timestamp 1757982896
transform 1 0 17600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_314
timestamp 1757982896
transform 1 0 19100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_315
timestamp 1757982896
transform 1 0 20600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_316
timestamp 1757982896
transform 1 0 22100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_317
timestamp 1757982896
transform 1 0 23600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_318
timestamp 1757982896
transform 1 0 25100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_319
timestamp 1757982896
transform 1 0 26600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_320
timestamp 1757982896
transform 1 0 28100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_321
timestamp 1757982896
transform 1 0 29600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_322
timestamp 1757982896
transform 1 0 31100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_323
timestamp 1757982896
transform 1 0 32600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_324
timestamp 1757982896
transform 1 0 34100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_325
timestamp 1757982896
transform 1 0 35600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_326
timestamp 1757982896
transform 1 0 37100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_327
timestamp 1757982896
transform 1 0 38600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_328
timestamp 1757982896
transform 1 0 40100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_329
timestamp 1757982896
transform 1 0 41600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_330
timestamp 1757982896
transform 1 0 43100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_331
timestamp 1757982896
transform 1 0 44600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_332
timestamp 1757982896
transform 1 0 46100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_333
timestamp 1757982896
transform 1 0 47600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_334
timestamp 1757982896
transform 1 0 49100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_335
timestamp 1757982896
transform 1 0 50600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_336
timestamp 1757982896
transform 1 0 52100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_337
timestamp 1757982896
transform 1 0 53600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_338
timestamp 1757982896
transform 1 0 55100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_339
timestamp 1757982896
transform 1 0 56600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_340
timestamp 1757982896
transform 1 0 58100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_341
timestamp 1757982896
transform 1 0 59600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_342
timestamp 1757982896
transform 1 0 61100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_343
timestamp 1757982896
transform 1 0 62600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_344
timestamp 1757982896
transform 1 0 64100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_345
timestamp 1757982896
transform 1 0 65600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_346
timestamp 1757982896
transform 1 0 67100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_347
timestamp 1757982896
transform 1 0 68600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_348
timestamp 1757982896
transform 1 0 70100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_349
timestamp 1757982896
transform 1 0 71600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_350
timestamp 1757982896
transform 1 0 73100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_351
timestamp 1757982896
transform 1 0 74600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_352
timestamp 1757982896
transform 1 0 76100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_353
timestamp 1757982896
transform 1 0 77600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_354
timestamp 1757982896
transform 1 0 79100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_355
timestamp 1757982896
transform 1 0 80600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_356
timestamp 1757982896
transform 1 0 82100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_357
timestamp 1757982896
transform 1 0 83600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_358
timestamp 1757982896
transform 1 0 85100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_359
timestamp 1757982896
transform 1 0 86600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_360
timestamp 1757982896
transform 1 0 88100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_361
timestamp 1757982896
transform 1 0 89600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_362
timestamp 1757982896
transform 1 0 91100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_363
timestamp 1757982896
transform 1 0 92600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_364
timestamp 1757982896
transform 1 0 94100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_365
timestamp 1757982896
transform 1 0 95600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_366
timestamp 1757982896
transform 1 0 97100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_367
timestamp 1757982896
transform 1 0 98600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_368
timestamp 1757982896
transform 1 0 100100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_369
timestamp 1757982896
transform 1 0 101600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_370
timestamp 1757982896
transform 1 0 103100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_371
timestamp 1757982896
transform 1 0 104600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_372
timestamp 1757982896
transform 1 0 106100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_373
timestamp 1757982896
transform 1 0 107600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_374
timestamp 1757982896
transform 1 0 109100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_375
timestamp 1757982896
transform 1 0 110600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_376
timestamp 1757982896
transform 1 0 112100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_377
timestamp 1757982896
transform 1 0 113600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_378
timestamp 1757982896
transform 1 0 115100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_379
timestamp 1757982896
transform 1 0 116600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_380
timestamp 1757982896
transform 1 0 118100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_381
timestamp 1757982896
transform 1 0 119600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_382
timestamp 1757982896
transform 1 0 121100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_383
timestamp 1757982896
transform 1 0 122600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_384
timestamp 1757982896
transform 1 0 124100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_385
timestamp 1757982896
transform 1 0 125600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_386
timestamp 1757982896
transform 1 0 127100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_387
timestamp 1757982896
transform 1 0 128600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_388
timestamp 1757982896
transform 1 0 130100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_389
timestamp 1757982896
transform 1 0 131600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_390
timestamp 1757982896
transform 1 0 133100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_391
timestamp 1757982896
transform 1 0 134600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_392
timestamp 1757982896
transform 1 0 136100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_393
timestamp 1757982896
transform 1 0 137600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_394
timestamp 1757982896
transform 1 0 139100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_395
timestamp 1757982896
transform 1 0 140600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_396
timestamp 1757982896
transform 1 0 142100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_397
timestamp 1757982896
transform 1 0 143600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_398
timestamp 1757982896
transform 1 0 145100 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_399
timestamp 1757982896
transform 1 0 146600 0 1 -3150
box 1820 -1430 3480 230
use pixel  pixel_400
timestamp 1757982896
transform 1 0 -1900 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_401
timestamp 1757982896
transform 1 0 -400 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_402
timestamp 1757982896
transform 1 0 1100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_403
timestamp 1757982896
transform 1 0 2600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_404
timestamp 1757982896
transform 1 0 4100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_405
timestamp 1757982896
transform 1 0 5600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_406
timestamp 1757982896
transform 1 0 7100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_407
timestamp 1757982896
transform 1 0 8600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_408
timestamp 1757982896
transform 1 0 10100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_409
timestamp 1757982896
transform 1 0 11600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_410
timestamp 1757982896
transform 1 0 13100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_411
timestamp 1757982896
transform 1 0 14600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_412
timestamp 1757982896
transform 1 0 16100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_413
timestamp 1757982896
transform 1 0 17600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_414
timestamp 1757982896
transform 1 0 19100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_415
timestamp 1757982896
transform 1 0 20600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_416
timestamp 1757982896
transform 1 0 22100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_417
timestamp 1757982896
transform 1 0 23600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_418
timestamp 1757982896
transform 1 0 25100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_419
timestamp 1757982896
transform 1 0 26600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_420
timestamp 1757982896
transform 1 0 28100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_421
timestamp 1757982896
transform 1 0 29600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_422
timestamp 1757982896
transform 1 0 31100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_423
timestamp 1757982896
transform 1 0 32600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_424
timestamp 1757982896
transform 1 0 34100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_425
timestamp 1757982896
transform 1 0 35600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_426
timestamp 1757982896
transform 1 0 37100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_427
timestamp 1757982896
transform 1 0 38600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_428
timestamp 1757982896
transform 1 0 40100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_429
timestamp 1757982896
transform 1 0 41600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_430
timestamp 1757982896
transform 1 0 43100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_431
timestamp 1757982896
transform 1 0 44600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_432
timestamp 1757982896
transform 1 0 46100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_433
timestamp 1757982896
transform 1 0 47600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_434
timestamp 1757982896
transform 1 0 49100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_435
timestamp 1757982896
transform 1 0 50600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_436
timestamp 1757982896
transform 1 0 52100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_437
timestamp 1757982896
transform 1 0 53600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_438
timestamp 1757982896
transform 1 0 55100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_439
timestamp 1757982896
transform 1 0 56600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_440
timestamp 1757982896
transform 1 0 58100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_441
timestamp 1757982896
transform 1 0 59600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_442
timestamp 1757982896
transform 1 0 61100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_443
timestamp 1757982896
transform 1 0 62600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_444
timestamp 1757982896
transform 1 0 64100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_445
timestamp 1757982896
transform 1 0 65600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_446
timestamp 1757982896
transform 1 0 67100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_447
timestamp 1757982896
transform 1 0 68600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_448
timestamp 1757982896
transform 1 0 70100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_449
timestamp 1757982896
transform 1 0 71600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_450
timestamp 1757982896
transform 1 0 73100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_451
timestamp 1757982896
transform 1 0 74600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_452
timestamp 1757982896
transform 1 0 76100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_453
timestamp 1757982896
transform 1 0 77600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_454
timestamp 1757982896
transform 1 0 79100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_455
timestamp 1757982896
transform 1 0 80600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_456
timestamp 1757982896
transform 1 0 82100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_457
timestamp 1757982896
transform 1 0 83600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_458
timestamp 1757982896
transform 1 0 85100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_459
timestamp 1757982896
transform 1 0 86600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_460
timestamp 1757982896
transform 1 0 88100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_461
timestamp 1757982896
transform 1 0 89600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_462
timestamp 1757982896
transform 1 0 91100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_463
timestamp 1757982896
transform 1 0 92600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_464
timestamp 1757982896
transform 1 0 94100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_465
timestamp 1757982896
transform 1 0 95600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_466
timestamp 1757982896
transform 1 0 97100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_467
timestamp 1757982896
transform 1 0 98600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_468
timestamp 1757982896
transform 1 0 100100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_469
timestamp 1757982896
transform 1 0 101600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_470
timestamp 1757982896
transform 1 0 103100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_471
timestamp 1757982896
transform 1 0 104600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_472
timestamp 1757982896
transform 1 0 106100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_473
timestamp 1757982896
transform 1 0 107600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_474
timestamp 1757982896
transform 1 0 109100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_475
timestamp 1757982896
transform 1 0 110600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_476
timestamp 1757982896
transform 1 0 112100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_477
timestamp 1757982896
transform 1 0 113600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_478
timestamp 1757982896
transform 1 0 115100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_479
timestamp 1757982896
transform 1 0 116600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_480
timestamp 1757982896
transform 1 0 118100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_481
timestamp 1757982896
transform 1 0 119600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_482
timestamp 1757982896
transform 1 0 121100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_483
timestamp 1757982896
transform 1 0 122600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_484
timestamp 1757982896
transform 1 0 124100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_485
timestamp 1757982896
transform 1 0 125600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_486
timestamp 1757982896
transform 1 0 127100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_487
timestamp 1757982896
transform 1 0 128600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_488
timestamp 1757982896
transform 1 0 130100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_489
timestamp 1757982896
transform 1 0 131600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_490
timestamp 1757982896
transform 1 0 133100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_491
timestamp 1757982896
transform 1 0 134600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_492
timestamp 1757982896
transform 1 0 136100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_493
timestamp 1757982896
transform 1 0 137600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_494
timestamp 1757982896
transform 1 0 139100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_495
timestamp 1757982896
transform 1 0 140600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_496
timestamp 1757982896
transform 1 0 142100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_497
timestamp 1757982896
transform 1 0 143600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_498
timestamp 1757982896
transform 1 0 145100 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_499
timestamp 1757982896
transform 1 0 146600 0 1 -4650
box 1820 -1430 3480 230
use pixel  pixel_500
timestamp 1757982896
transform 1 0 -1900 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_501
timestamp 1757982896
transform 1 0 -400 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_502
timestamp 1757982896
transform 1 0 1100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_503
timestamp 1757982896
transform 1 0 2600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_504
timestamp 1757982896
transform 1 0 4100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_505
timestamp 1757982896
transform 1 0 5600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_506
timestamp 1757982896
transform 1 0 7100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_507
timestamp 1757982896
transform 1 0 8600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_508
timestamp 1757982896
transform 1 0 10100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_509
timestamp 1757982896
transform 1 0 11600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_510
timestamp 1757982896
transform 1 0 13100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_511
timestamp 1757982896
transform 1 0 14600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_512
timestamp 1757982896
transform 1 0 16100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_513
timestamp 1757982896
transform 1 0 17600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_514
timestamp 1757982896
transform 1 0 19100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_515
timestamp 1757982896
transform 1 0 20600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_516
timestamp 1757982896
transform 1 0 22100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_517
timestamp 1757982896
transform 1 0 23600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_518
timestamp 1757982896
transform 1 0 25100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_519
timestamp 1757982896
transform 1 0 26600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_520
timestamp 1757982896
transform 1 0 28100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_521
timestamp 1757982896
transform 1 0 29600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_522
timestamp 1757982896
transform 1 0 31100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_523
timestamp 1757982896
transform 1 0 32600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_524
timestamp 1757982896
transform 1 0 34100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_525
timestamp 1757982896
transform 1 0 35600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_526
timestamp 1757982896
transform 1 0 37100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_527
timestamp 1757982896
transform 1 0 38600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_528
timestamp 1757982896
transform 1 0 40100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_529
timestamp 1757982896
transform 1 0 41600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_530
timestamp 1757982896
transform 1 0 43100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_531
timestamp 1757982896
transform 1 0 44600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_532
timestamp 1757982896
transform 1 0 46100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_533
timestamp 1757982896
transform 1 0 47600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_534
timestamp 1757982896
transform 1 0 49100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_535
timestamp 1757982896
transform 1 0 50600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_536
timestamp 1757982896
transform 1 0 52100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_537
timestamp 1757982896
transform 1 0 53600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_538
timestamp 1757982896
transform 1 0 55100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_539
timestamp 1757982896
transform 1 0 56600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_540
timestamp 1757982896
transform 1 0 58100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_541
timestamp 1757982896
transform 1 0 59600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_542
timestamp 1757982896
transform 1 0 61100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_543
timestamp 1757982896
transform 1 0 62600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_544
timestamp 1757982896
transform 1 0 64100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_545
timestamp 1757982896
transform 1 0 65600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_546
timestamp 1757982896
transform 1 0 67100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_547
timestamp 1757982896
transform 1 0 68600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_548
timestamp 1757982896
transform 1 0 70100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_549
timestamp 1757982896
transform 1 0 71600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_550
timestamp 1757982896
transform 1 0 73100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_551
timestamp 1757982896
transform 1 0 74600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_552
timestamp 1757982896
transform 1 0 76100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_553
timestamp 1757982896
transform 1 0 77600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_554
timestamp 1757982896
transform 1 0 79100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_555
timestamp 1757982896
transform 1 0 80600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_556
timestamp 1757982896
transform 1 0 82100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_557
timestamp 1757982896
transform 1 0 83600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_558
timestamp 1757982896
transform 1 0 85100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_559
timestamp 1757982896
transform 1 0 86600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_560
timestamp 1757982896
transform 1 0 88100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_561
timestamp 1757982896
transform 1 0 89600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_562
timestamp 1757982896
transform 1 0 91100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_563
timestamp 1757982896
transform 1 0 92600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_564
timestamp 1757982896
transform 1 0 94100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_565
timestamp 1757982896
transform 1 0 95600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_566
timestamp 1757982896
transform 1 0 97100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_567
timestamp 1757982896
transform 1 0 98600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_568
timestamp 1757982896
transform 1 0 100100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_569
timestamp 1757982896
transform 1 0 101600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_570
timestamp 1757982896
transform 1 0 103100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_571
timestamp 1757982896
transform 1 0 104600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_572
timestamp 1757982896
transform 1 0 106100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_573
timestamp 1757982896
transform 1 0 107600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_574
timestamp 1757982896
transform 1 0 109100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_575
timestamp 1757982896
transform 1 0 110600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_576
timestamp 1757982896
transform 1 0 112100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_577
timestamp 1757982896
transform 1 0 113600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_578
timestamp 1757982896
transform 1 0 115100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_579
timestamp 1757982896
transform 1 0 116600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_580
timestamp 1757982896
transform 1 0 118100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_581
timestamp 1757982896
transform 1 0 119600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_582
timestamp 1757982896
transform 1 0 121100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_583
timestamp 1757982896
transform 1 0 122600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_584
timestamp 1757982896
transform 1 0 124100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_585
timestamp 1757982896
transform 1 0 125600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_586
timestamp 1757982896
transform 1 0 127100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_587
timestamp 1757982896
transform 1 0 128600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_588
timestamp 1757982896
transform 1 0 130100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_589
timestamp 1757982896
transform 1 0 131600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_590
timestamp 1757982896
transform 1 0 133100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_591
timestamp 1757982896
transform 1 0 134600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_592
timestamp 1757982896
transform 1 0 136100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_593
timestamp 1757982896
transform 1 0 137600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_594
timestamp 1757982896
transform 1 0 139100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_595
timestamp 1757982896
transform 1 0 140600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_596
timestamp 1757982896
transform 1 0 142100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_597
timestamp 1757982896
transform 1 0 143600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_598
timestamp 1757982896
transform 1 0 145100 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_599
timestamp 1757982896
transform 1 0 146600 0 1 -6150
box 1820 -1430 3480 230
use pixel  pixel_600
timestamp 1757982896
transform 1 0 -1900 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_601
timestamp 1757982896
transform 1 0 -400 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_602
timestamp 1757982896
transform 1 0 1100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_603
timestamp 1757982896
transform 1 0 2600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_604
timestamp 1757982896
transform 1 0 4100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_605
timestamp 1757982896
transform 1 0 5600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_606
timestamp 1757982896
transform 1 0 7100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_607
timestamp 1757982896
transform 1 0 8600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_608
timestamp 1757982896
transform 1 0 10100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_609
timestamp 1757982896
transform 1 0 11600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_610
timestamp 1757982896
transform 1 0 13100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_611
timestamp 1757982896
transform 1 0 14600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_612
timestamp 1757982896
transform 1 0 16100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_613
timestamp 1757982896
transform 1 0 17600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_614
timestamp 1757982896
transform 1 0 19100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_615
timestamp 1757982896
transform 1 0 20600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_616
timestamp 1757982896
transform 1 0 22100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_617
timestamp 1757982896
transform 1 0 23600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_618
timestamp 1757982896
transform 1 0 25100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_619
timestamp 1757982896
transform 1 0 26600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_620
timestamp 1757982896
transform 1 0 28100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_621
timestamp 1757982896
transform 1 0 29600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_622
timestamp 1757982896
transform 1 0 31100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_623
timestamp 1757982896
transform 1 0 32600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_624
timestamp 1757982896
transform 1 0 34100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_625
timestamp 1757982896
transform 1 0 35600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_626
timestamp 1757982896
transform 1 0 37100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_627
timestamp 1757982896
transform 1 0 38600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_628
timestamp 1757982896
transform 1 0 40100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_629
timestamp 1757982896
transform 1 0 41600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_630
timestamp 1757982896
transform 1 0 43100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_631
timestamp 1757982896
transform 1 0 44600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_632
timestamp 1757982896
transform 1 0 46100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_633
timestamp 1757982896
transform 1 0 47600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_634
timestamp 1757982896
transform 1 0 49100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_635
timestamp 1757982896
transform 1 0 50600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_636
timestamp 1757982896
transform 1 0 52100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_637
timestamp 1757982896
transform 1 0 53600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_638
timestamp 1757982896
transform 1 0 55100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_639
timestamp 1757982896
transform 1 0 56600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_640
timestamp 1757982896
transform 1 0 58100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_641
timestamp 1757982896
transform 1 0 59600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_642
timestamp 1757982896
transform 1 0 61100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_643
timestamp 1757982896
transform 1 0 62600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_644
timestamp 1757982896
transform 1 0 64100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_645
timestamp 1757982896
transform 1 0 65600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_646
timestamp 1757982896
transform 1 0 67100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_647
timestamp 1757982896
transform 1 0 68600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_648
timestamp 1757982896
transform 1 0 70100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_649
timestamp 1757982896
transform 1 0 71600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_650
timestamp 1757982896
transform 1 0 73100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_651
timestamp 1757982896
transform 1 0 74600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_652
timestamp 1757982896
transform 1 0 76100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_653
timestamp 1757982896
transform 1 0 77600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_654
timestamp 1757982896
transform 1 0 79100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_655
timestamp 1757982896
transform 1 0 80600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_656
timestamp 1757982896
transform 1 0 82100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_657
timestamp 1757982896
transform 1 0 83600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_658
timestamp 1757982896
transform 1 0 85100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_659
timestamp 1757982896
transform 1 0 86600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_660
timestamp 1757982896
transform 1 0 88100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_661
timestamp 1757982896
transform 1 0 89600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_662
timestamp 1757982896
transform 1 0 91100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_663
timestamp 1757982896
transform 1 0 92600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_664
timestamp 1757982896
transform 1 0 94100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_665
timestamp 1757982896
transform 1 0 95600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_666
timestamp 1757982896
transform 1 0 97100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_667
timestamp 1757982896
transform 1 0 98600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_668
timestamp 1757982896
transform 1 0 100100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_669
timestamp 1757982896
transform 1 0 101600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_670
timestamp 1757982896
transform 1 0 103100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_671
timestamp 1757982896
transform 1 0 104600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_672
timestamp 1757982896
transform 1 0 106100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_673
timestamp 1757982896
transform 1 0 107600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_674
timestamp 1757982896
transform 1 0 109100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_675
timestamp 1757982896
transform 1 0 110600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_676
timestamp 1757982896
transform 1 0 112100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_677
timestamp 1757982896
transform 1 0 113600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_678
timestamp 1757982896
transform 1 0 115100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_679
timestamp 1757982896
transform 1 0 116600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_680
timestamp 1757982896
transform 1 0 118100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_681
timestamp 1757982896
transform 1 0 119600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_682
timestamp 1757982896
transform 1 0 121100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_683
timestamp 1757982896
transform 1 0 122600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_684
timestamp 1757982896
transform 1 0 124100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_685
timestamp 1757982896
transform 1 0 125600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_686
timestamp 1757982896
transform 1 0 127100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_687
timestamp 1757982896
transform 1 0 128600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_688
timestamp 1757982896
transform 1 0 130100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_689
timestamp 1757982896
transform 1 0 131600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_690
timestamp 1757982896
transform 1 0 133100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_691
timestamp 1757982896
transform 1 0 134600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_692
timestamp 1757982896
transform 1 0 136100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_693
timestamp 1757982896
transform 1 0 137600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_694
timestamp 1757982896
transform 1 0 139100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_695
timestamp 1757982896
transform 1 0 140600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_696
timestamp 1757982896
transform 1 0 142100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_697
timestamp 1757982896
transform 1 0 143600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_698
timestamp 1757982896
transform 1 0 145100 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_699
timestamp 1757982896
transform 1 0 146600 0 1 -7650
box 1820 -1430 3480 230
use pixel  pixel_700
timestamp 1757982896
transform 1 0 -1900 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_701
timestamp 1757982896
transform 1 0 -400 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_702
timestamp 1757982896
transform 1 0 1100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_703
timestamp 1757982896
transform 1 0 2600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_704
timestamp 1757982896
transform 1 0 4100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_705
timestamp 1757982896
transform 1 0 5600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_706
timestamp 1757982896
transform 1 0 7100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_707
timestamp 1757982896
transform 1 0 8600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_708
timestamp 1757982896
transform 1 0 10100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_709
timestamp 1757982896
transform 1 0 11600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_710
timestamp 1757982896
transform 1 0 13100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_711
timestamp 1757982896
transform 1 0 14600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_712
timestamp 1757982896
transform 1 0 16100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_713
timestamp 1757982896
transform 1 0 17600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_714
timestamp 1757982896
transform 1 0 19100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_715
timestamp 1757982896
transform 1 0 20600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_716
timestamp 1757982896
transform 1 0 22100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_717
timestamp 1757982896
transform 1 0 23600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_718
timestamp 1757982896
transform 1 0 25100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_719
timestamp 1757982896
transform 1 0 26600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_720
timestamp 1757982896
transform 1 0 28100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_721
timestamp 1757982896
transform 1 0 29600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_722
timestamp 1757982896
transform 1 0 31100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_723
timestamp 1757982896
transform 1 0 32600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_724
timestamp 1757982896
transform 1 0 34100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_725
timestamp 1757982896
transform 1 0 35600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_726
timestamp 1757982896
transform 1 0 37100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_727
timestamp 1757982896
transform 1 0 38600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_728
timestamp 1757982896
transform 1 0 40100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_729
timestamp 1757982896
transform 1 0 41600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_730
timestamp 1757982896
transform 1 0 43100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_731
timestamp 1757982896
transform 1 0 44600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_732
timestamp 1757982896
transform 1 0 46100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_733
timestamp 1757982896
transform 1 0 47600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_734
timestamp 1757982896
transform 1 0 49100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_735
timestamp 1757982896
transform 1 0 50600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_736
timestamp 1757982896
transform 1 0 52100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_737
timestamp 1757982896
transform 1 0 53600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_738
timestamp 1757982896
transform 1 0 55100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_739
timestamp 1757982896
transform 1 0 56600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_740
timestamp 1757982896
transform 1 0 58100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_741
timestamp 1757982896
transform 1 0 59600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_742
timestamp 1757982896
transform 1 0 61100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_743
timestamp 1757982896
transform 1 0 62600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_744
timestamp 1757982896
transform 1 0 64100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_745
timestamp 1757982896
transform 1 0 65600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_746
timestamp 1757982896
transform 1 0 67100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_747
timestamp 1757982896
transform 1 0 68600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_748
timestamp 1757982896
transform 1 0 70100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_749
timestamp 1757982896
transform 1 0 71600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_750
timestamp 1757982896
transform 1 0 73100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_751
timestamp 1757982896
transform 1 0 74600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_752
timestamp 1757982896
transform 1 0 76100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_753
timestamp 1757982896
transform 1 0 77600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_754
timestamp 1757982896
transform 1 0 79100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_755
timestamp 1757982896
transform 1 0 80600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_756
timestamp 1757982896
transform 1 0 82100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_757
timestamp 1757982896
transform 1 0 83600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_758
timestamp 1757982896
transform 1 0 85100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_759
timestamp 1757982896
transform 1 0 86600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_760
timestamp 1757982896
transform 1 0 88100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_761
timestamp 1757982896
transform 1 0 89600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_762
timestamp 1757982896
transform 1 0 91100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_763
timestamp 1757982896
transform 1 0 92600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_764
timestamp 1757982896
transform 1 0 94100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_765
timestamp 1757982896
transform 1 0 95600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_766
timestamp 1757982896
transform 1 0 97100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_767
timestamp 1757982896
transform 1 0 98600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_768
timestamp 1757982896
transform 1 0 100100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_769
timestamp 1757982896
transform 1 0 101600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_770
timestamp 1757982896
transform 1 0 103100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_771
timestamp 1757982896
transform 1 0 104600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_772
timestamp 1757982896
transform 1 0 106100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_773
timestamp 1757982896
transform 1 0 107600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_774
timestamp 1757982896
transform 1 0 109100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_775
timestamp 1757982896
transform 1 0 110600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_776
timestamp 1757982896
transform 1 0 112100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_777
timestamp 1757982896
transform 1 0 113600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_778
timestamp 1757982896
transform 1 0 115100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_779
timestamp 1757982896
transform 1 0 116600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_780
timestamp 1757982896
transform 1 0 118100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_781
timestamp 1757982896
transform 1 0 119600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_782
timestamp 1757982896
transform 1 0 121100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_783
timestamp 1757982896
transform 1 0 122600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_784
timestamp 1757982896
transform 1 0 124100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_785
timestamp 1757982896
transform 1 0 125600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_786
timestamp 1757982896
transform 1 0 127100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_787
timestamp 1757982896
transform 1 0 128600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_788
timestamp 1757982896
transform 1 0 130100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_789
timestamp 1757982896
transform 1 0 131600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_790
timestamp 1757982896
transform 1 0 133100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_791
timestamp 1757982896
transform 1 0 134600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_792
timestamp 1757982896
transform 1 0 136100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_793
timestamp 1757982896
transform 1 0 137600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_794
timestamp 1757982896
transform 1 0 139100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_795
timestamp 1757982896
transform 1 0 140600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_796
timestamp 1757982896
transform 1 0 142100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_797
timestamp 1757982896
transform 1 0 143600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_798
timestamp 1757982896
transform 1 0 145100 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_799
timestamp 1757982896
transform 1 0 146600 0 1 -9150
box 1820 -1430 3480 230
use pixel  pixel_800
timestamp 1757982896
transform 1 0 -1900 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_801
timestamp 1757982896
transform 1 0 -400 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_802
timestamp 1757982896
transform 1 0 1100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_803
timestamp 1757982896
transform 1 0 2600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_804
timestamp 1757982896
transform 1 0 4100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_805
timestamp 1757982896
transform 1 0 5600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_806
timestamp 1757982896
transform 1 0 7100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_807
timestamp 1757982896
transform 1 0 8600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_808
timestamp 1757982896
transform 1 0 10100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_809
timestamp 1757982896
transform 1 0 11600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_810
timestamp 1757982896
transform 1 0 13100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_811
timestamp 1757982896
transform 1 0 14600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_812
timestamp 1757982896
transform 1 0 16100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_813
timestamp 1757982896
transform 1 0 17600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_814
timestamp 1757982896
transform 1 0 19100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_815
timestamp 1757982896
transform 1 0 20600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_816
timestamp 1757982896
transform 1 0 22100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_817
timestamp 1757982896
transform 1 0 23600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_818
timestamp 1757982896
transform 1 0 25100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_819
timestamp 1757982896
transform 1 0 26600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_820
timestamp 1757982896
transform 1 0 28100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_821
timestamp 1757982896
transform 1 0 29600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_822
timestamp 1757982896
transform 1 0 31100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_823
timestamp 1757982896
transform 1 0 32600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_824
timestamp 1757982896
transform 1 0 34100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_825
timestamp 1757982896
transform 1 0 35600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_826
timestamp 1757982896
transform 1 0 37100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_827
timestamp 1757982896
transform 1 0 38600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_828
timestamp 1757982896
transform 1 0 40100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_829
timestamp 1757982896
transform 1 0 41600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_830
timestamp 1757982896
transform 1 0 43100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_831
timestamp 1757982896
transform 1 0 44600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_832
timestamp 1757982896
transform 1 0 46100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_833
timestamp 1757982896
transform 1 0 47600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_834
timestamp 1757982896
transform 1 0 49100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_835
timestamp 1757982896
transform 1 0 50600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_836
timestamp 1757982896
transform 1 0 52100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_837
timestamp 1757982896
transform 1 0 53600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_838
timestamp 1757982896
transform 1 0 55100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_839
timestamp 1757982896
transform 1 0 56600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_840
timestamp 1757982896
transform 1 0 58100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_841
timestamp 1757982896
transform 1 0 59600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_842
timestamp 1757982896
transform 1 0 61100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_843
timestamp 1757982896
transform 1 0 62600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_844
timestamp 1757982896
transform 1 0 64100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_845
timestamp 1757982896
transform 1 0 65600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_846
timestamp 1757982896
transform 1 0 67100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_847
timestamp 1757982896
transform 1 0 68600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_848
timestamp 1757982896
transform 1 0 70100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_849
timestamp 1757982896
transform 1 0 71600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_850
timestamp 1757982896
transform 1 0 73100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_851
timestamp 1757982896
transform 1 0 74600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_852
timestamp 1757982896
transform 1 0 76100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_853
timestamp 1757982896
transform 1 0 77600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_854
timestamp 1757982896
transform 1 0 79100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_855
timestamp 1757982896
transform 1 0 80600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_856
timestamp 1757982896
transform 1 0 82100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_857
timestamp 1757982896
transform 1 0 83600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_858
timestamp 1757982896
transform 1 0 85100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_859
timestamp 1757982896
transform 1 0 86600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_860
timestamp 1757982896
transform 1 0 88100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_861
timestamp 1757982896
transform 1 0 89600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_862
timestamp 1757982896
transform 1 0 91100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_863
timestamp 1757982896
transform 1 0 92600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_864
timestamp 1757982896
transform 1 0 94100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_865
timestamp 1757982896
transform 1 0 95600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_866
timestamp 1757982896
transform 1 0 97100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_867
timestamp 1757982896
transform 1 0 98600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_868
timestamp 1757982896
transform 1 0 100100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_869
timestamp 1757982896
transform 1 0 101600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_870
timestamp 1757982896
transform 1 0 103100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_871
timestamp 1757982896
transform 1 0 104600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_872
timestamp 1757982896
transform 1 0 106100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_873
timestamp 1757982896
transform 1 0 107600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_874
timestamp 1757982896
transform 1 0 109100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_875
timestamp 1757982896
transform 1 0 110600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_876
timestamp 1757982896
transform 1 0 112100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_877
timestamp 1757982896
transform 1 0 113600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_878
timestamp 1757982896
transform 1 0 115100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_879
timestamp 1757982896
transform 1 0 116600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_880
timestamp 1757982896
transform 1 0 118100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_881
timestamp 1757982896
transform 1 0 119600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_882
timestamp 1757982896
transform 1 0 121100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_883
timestamp 1757982896
transform 1 0 122600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_884
timestamp 1757982896
transform 1 0 124100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_885
timestamp 1757982896
transform 1 0 125600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_886
timestamp 1757982896
transform 1 0 127100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_887
timestamp 1757982896
transform 1 0 128600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_888
timestamp 1757982896
transform 1 0 130100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_889
timestamp 1757982896
transform 1 0 131600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_890
timestamp 1757982896
transform 1 0 133100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_891
timestamp 1757982896
transform 1 0 134600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_892
timestamp 1757982896
transform 1 0 136100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_893
timestamp 1757982896
transform 1 0 137600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_894
timestamp 1757982896
transform 1 0 139100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_895
timestamp 1757982896
transform 1 0 140600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_896
timestamp 1757982896
transform 1 0 142100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_897
timestamp 1757982896
transform 1 0 143600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_898
timestamp 1757982896
transform 1 0 145100 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_899
timestamp 1757982896
transform 1 0 146600 0 1 -10650
box 1820 -1430 3480 230
use pixel  pixel_900
timestamp 1757982896
transform 1 0 -1900 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_901
timestamp 1757982896
transform 1 0 -400 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_902
timestamp 1757982896
transform 1 0 1100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_903
timestamp 1757982896
transform 1 0 2600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_904
timestamp 1757982896
transform 1 0 4100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_905
timestamp 1757982896
transform 1 0 5600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_906
timestamp 1757982896
transform 1 0 7100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_907
timestamp 1757982896
transform 1 0 8600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_908
timestamp 1757982896
transform 1 0 10100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_909
timestamp 1757982896
transform 1 0 11600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_910
timestamp 1757982896
transform 1 0 13100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_911
timestamp 1757982896
transform 1 0 14600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_912
timestamp 1757982896
transform 1 0 16100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_913
timestamp 1757982896
transform 1 0 17600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_914
timestamp 1757982896
transform 1 0 19100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_915
timestamp 1757982896
transform 1 0 20600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_916
timestamp 1757982896
transform 1 0 22100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_917
timestamp 1757982896
transform 1 0 23600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_918
timestamp 1757982896
transform 1 0 25100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_919
timestamp 1757982896
transform 1 0 26600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_920
timestamp 1757982896
transform 1 0 28100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_921
timestamp 1757982896
transform 1 0 29600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_922
timestamp 1757982896
transform 1 0 31100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_923
timestamp 1757982896
transform 1 0 32600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_924
timestamp 1757982896
transform 1 0 34100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_925
timestamp 1757982896
transform 1 0 35600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_926
timestamp 1757982896
transform 1 0 37100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_927
timestamp 1757982896
transform 1 0 38600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_928
timestamp 1757982896
transform 1 0 40100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_929
timestamp 1757982896
transform 1 0 41600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_930
timestamp 1757982896
transform 1 0 43100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_931
timestamp 1757982896
transform 1 0 44600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_932
timestamp 1757982896
transform 1 0 46100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_933
timestamp 1757982896
transform 1 0 47600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_934
timestamp 1757982896
transform 1 0 49100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_935
timestamp 1757982896
transform 1 0 50600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_936
timestamp 1757982896
transform 1 0 52100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_937
timestamp 1757982896
transform 1 0 53600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_938
timestamp 1757982896
transform 1 0 55100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_939
timestamp 1757982896
transform 1 0 56600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_940
timestamp 1757982896
transform 1 0 58100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_941
timestamp 1757982896
transform 1 0 59600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_942
timestamp 1757982896
transform 1 0 61100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_943
timestamp 1757982896
transform 1 0 62600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_944
timestamp 1757982896
transform 1 0 64100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_945
timestamp 1757982896
transform 1 0 65600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_946
timestamp 1757982896
transform 1 0 67100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_947
timestamp 1757982896
transform 1 0 68600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_948
timestamp 1757982896
transform 1 0 70100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_949
timestamp 1757982896
transform 1 0 71600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_950
timestamp 1757982896
transform 1 0 73100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_951
timestamp 1757982896
transform 1 0 74600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_952
timestamp 1757982896
transform 1 0 76100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_953
timestamp 1757982896
transform 1 0 77600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_954
timestamp 1757982896
transform 1 0 79100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_955
timestamp 1757982896
transform 1 0 80600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_956
timestamp 1757982896
transform 1 0 82100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_957
timestamp 1757982896
transform 1 0 83600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_958
timestamp 1757982896
transform 1 0 85100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_959
timestamp 1757982896
transform 1 0 86600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_960
timestamp 1757982896
transform 1 0 88100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_961
timestamp 1757982896
transform 1 0 89600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_962
timestamp 1757982896
transform 1 0 91100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_963
timestamp 1757982896
transform 1 0 92600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_964
timestamp 1757982896
transform 1 0 94100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_965
timestamp 1757982896
transform 1 0 95600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_966
timestamp 1757982896
transform 1 0 97100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_967
timestamp 1757982896
transform 1 0 98600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_968
timestamp 1757982896
transform 1 0 100100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_969
timestamp 1757982896
transform 1 0 101600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_970
timestamp 1757982896
transform 1 0 103100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_971
timestamp 1757982896
transform 1 0 104600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_972
timestamp 1757982896
transform 1 0 106100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_973
timestamp 1757982896
transform 1 0 107600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_974
timestamp 1757982896
transform 1 0 109100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_975
timestamp 1757982896
transform 1 0 110600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_976
timestamp 1757982896
transform 1 0 112100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_977
timestamp 1757982896
transform 1 0 113600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_978
timestamp 1757982896
transform 1 0 115100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_979
timestamp 1757982896
transform 1 0 116600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_980
timestamp 1757982896
transform 1 0 118100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_981
timestamp 1757982896
transform 1 0 119600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_982
timestamp 1757982896
transform 1 0 121100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_983
timestamp 1757982896
transform 1 0 122600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_984
timestamp 1757982896
transform 1 0 124100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_985
timestamp 1757982896
transform 1 0 125600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_986
timestamp 1757982896
transform 1 0 127100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_987
timestamp 1757982896
transform 1 0 128600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_988
timestamp 1757982896
transform 1 0 130100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_989
timestamp 1757982896
transform 1 0 131600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_990
timestamp 1757982896
transform 1 0 133100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_991
timestamp 1757982896
transform 1 0 134600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_992
timestamp 1757982896
transform 1 0 136100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_993
timestamp 1757982896
transform 1 0 137600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_994
timestamp 1757982896
transform 1 0 139100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_995
timestamp 1757982896
transform 1 0 140600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_996
timestamp 1757982896
transform 1 0 142100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_997
timestamp 1757982896
transform 1 0 143600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_998
timestamp 1757982896
transform 1 0 145100 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_999
timestamp 1757982896
transform 1 0 146600 0 1 -12150
box 1820 -1430 3480 230
use pixel  pixel_1000
timestamp 1757982896
transform 1 0 -1900 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1001
timestamp 1757982896
transform 1 0 -400 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1002
timestamp 1757982896
transform 1 0 1100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1003
timestamp 1757982896
transform 1 0 2600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1004
timestamp 1757982896
transform 1 0 4100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1005
timestamp 1757982896
transform 1 0 5600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1006
timestamp 1757982896
transform 1 0 7100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1007
timestamp 1757982896
transform 1 0 8600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1008
timestamp 1757982896
transform 1 0 10100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1009
timestamp 1757982896
transform 1 0 11600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1010
timestamp 1757982896
transform 1 0 13100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1011
timestamp 1757982896
transform 1 0 14600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1012
timestamp 1757982896
transform 1 0 16100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1013
timestamp 1757982896
transform 1 0 17600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1014
timestamp 1757982896
transform 1 0 19100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1015
timestamp 1757982896
transform 1 0 20600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1016
timestamp 1757982896
transform 1 0 22100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1017
timestamp 1757982896
transform 1 0 23600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1018
timestamp 1757982896
transform 1 0 25100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1019
timestamp 1757982896
transform 1 0 26600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1020
timestamp 1757982896
transform 1 0 28100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1021
timestamp 1757982896
transform 1 0 29600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1022
timestamp 1757982896
transform 1 0 31100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1023
timestamp 1757982896
transform 1 0 32600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1024
timestamp 1757982896
transform 1 0 34100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1025
timestamp 1757982896
transform 1 0 35600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1026
timestamp 1757982896
transform 1 0 37100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1027
timestamp 1757982896
transform 1 0 38600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1028
timestamp 1757982896
transform 1 0 40100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1029
timestamp 1757982896
transform 1 0 41600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1030
timestamp 1757982896
transform 1 0 43100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1031
timestamp 1757982896
transform 1 0 44600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1032
timestamp 1757982896
transform 1 0 46100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1033
timestamp 1757982896
transform 1 0 47600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1034
timestamp 1757982896
transform 1 0 49100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1035
timestamp 1757982896
transform 1 0 50600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1036
timestamp 1757982896
transform 1 0 52100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1037
timestamp 1757982896
transform 1 0 53600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1038
timestamp 1757982896
transform 1 0 55100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1039
timestamp 1757982896
transform 1 0 56600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1040
timestamp 1757982896
transform 1 0 58100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1041
timestamp 1757982896
transform 1 0 59600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1042
timestamp 1757982896
transform 1 0 61100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1043
timestamp 1757982896
transform 1 0 62600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1044
timestamp 1757982896
transform 1 0 64100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1045
timestamp 1757982896
transform 1 0 65600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1046
timestamp 1757982896
transform 1 0 67100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1047
timestamp 1757982896
transform 1 0 68600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1048
timestamp 1757982896
transform 1 0 70100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1049
timestamp 1757982896
transform 1 0 71600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1050
timestamp 1757982896
transform 1 0 73100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1051
timestamp 1757982896
transform 1 0 74600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1052
timestamp 1757982896
transform 1 0 76100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1053
timestamp 1757982896
transform 1 0 77600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1054
timestamp 1757982896
transform 1 0 79100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1055
timestamp 1757982896
transform 1 0 80600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1056
timestamp 1757982896
transform 1 0 82100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1057
timestamp 1757982896
transform 1 0 83600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1058
timestamp 1757982896
transform 1 0 85100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1059
timestamp 1757982896
transform 1 0 86600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1060
timestamp 1757982896
transform 1 0 88100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1061
timestamp 1757982896
transform 1 0 89600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1062
timestamp 1757982896
transform 1 0 91100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1063
timestamp 1757982896
transform 1 0 92600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1064
timestamp 1757982896
transform 1 0 94100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1065
timestamp 1757982896
transform 1 0 95600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1066
timestamp 1757982896
transform 1 0 97100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1067
timestamp 1757982896
transform 1 0 98600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1068
timestamp 1757982896
transform 1 0 100100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1069
timestamp 1757982896
transform 1 0 101600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1070
timestamp 1757982896
transform 1 0 103100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1071
timestamp 1757982896
transform 1 0 104600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1072
timestamp 1757982896
transform 1 0 106100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1073
timestamp 1757982896
transform 1 0 107600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1074
timestamp 1757982896
transform 1 0 109100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1075
timestamp 1757982896
transform 1 0 110600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1076
timestamp 1757982896
transform 1 0 112100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1077
timestamp 1757982896
transform 1 0 113600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1078
timestamp 1757982896
transform 1 0 115100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1079
timestamp 1757982896
transform 1 0 116600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1080
timestamp 1757982896
transform 1 0 118100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1081
timestamp 1757982896
transform 1 0 119600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1082
timestamp 1757982896
transform 1 0 121100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1083
timestamp 1757982896
transform 1 0 122600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1084
timestamp 1757982896
transform 1 0 124100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1085
timestamp 1757982896
transform 1 0 125600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1086
timestamp 1757982896
transform 1 0 127100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1087
timestamp 1757982896
transform 1 0 128600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1088
timestamp 1757982896
transform 1 0 130100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1089
timestamp 1757982896
transform 1 0 131600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1090
timestamp 1757982896
transform 1 0 133100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1091
timestamp 1757982896
transform 1 0 134600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1092
timestamp 1757982896
transform 1 0 136100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1093
timestamp 1757982896
transform 1 0 137600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1094
timestamp 1757982896
transform 1 0 139100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1095
timestamp 1757982896
transform 1 0 140600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1096
timestamp 1757982896
transform 1 0 142100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1097
timestamp 1757982896
transform 1 0 143600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1098
timestamp 1757982896
transform 1 0 145100 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1099
timestamp 1757982896
transform 1 0 146600 0 1 -13650
box 1820 -1430 3480 230
use pixel  pixel_1100
timestamp 1757982896
transform 1 0 -1900 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1101
timestamp 1757982896
transform 1 0 -400 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1102
timestamp 1757982896
transform 1 0 1100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1103
timestamp 1757982896
transform 1 0 2600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1104
timestamp 1757982896
transform 1 0 4100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1105
timestamp 1757982896
transform 1 0 5600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1106
timestamp 1757982896
transform 1 0 7100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1107
timestamp 1757982896
transform 1 0 8600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1108
timestamp 1757982896
transform 1 0 10100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1109
timestamp 1757982896
transform 1 0 11600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1110
timestamp 1757982896
transform 1 0 13100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1111
timestamp 1757982896
transform 1 0 14600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1112
timestamp 1757982896
transform 1 0 16100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1113
timestamp 1757982896
transform 1 0 17600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1114
timestamp 1757982896
transform 1 0 19100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1115
timestamp 1757982896
transform 1 0 20600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1116
timestamp 1757982896
transform 1 0 22100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1117
timestamp 1757982896
transform 1 0 23600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1118
timestamp 1757982896
transform 1 0 25100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1119
timestamp 1757982896
transform 1 0 26600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1120
timestamp 1757982896
transform 1 0 28100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1121
timestamp 1757982896
transform 1 0 29600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1122
timestamp 1757982896
transform 1 0 31100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1123
timestamp 1757982896
transform 1 0 32600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1124
timestamp 1757982896
transform 1 0 34100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1125
timestamp 1757982896
transform 1 0 35600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1126
timestamp 1757982896
transform 1 0 37100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1127
timestamp 1757982896
transform 1 0 38600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1128
timestamp 1757982896
transform 1 0 40100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1129
timestamp 1757982896
transform 1 0 41600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1130
timestamp 1757982896
transform 1 0 43100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1131
timestamp 1757982896
transform 1 0 44600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1132
timestamp 1757982896
transform 1 0 46100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1133
timestamp 1757982896
transform 1 0 47600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1134
timestamp 1757982896
transform 1 0 49100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1135
timestamp 1757982896
transform 1 0 50600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1136
timestamp 1757982896
transform 1 0 52100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1137
timestamp 1757982896
transform 1 0 53600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1138
timestamp 1757982896
transform 1 0 55100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1139
timestamp 1757982896
transform 1 0 56600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1140
timestamp 1757982896
transform 1 0 58100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1141
timestamp 1757982896
transform 1 0 59600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1142
timestamp 1757982896
transform 1 0 61100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1143
timestamp 1757982896
transform 1 0 62600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1144
timestamp 1757982896
transform 1 0 64100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1145
timestamp 1757982896
transform 1 0 65600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1146
timestamp 1757982896
transform 1 0 67100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1147
timestamp 1757982896
transform 1 0 68600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1148
timestamp 1757982896
transform 1 0 70100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1149
timestamp 1757982896
transform 1 0 71600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1150
timestamp 1757982896
transform 1 0 73100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1151
timestamp 1757982896
transform 1 0 74600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1152
timestamp 1757982896
transform 1 0 76100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1153
timestamp 1757982896
transform 1 0 77600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1154
timestamp 1757982896
transform 1 0 79100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1155
timestamp 1757982896
transform 1 0 80600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1156
timestamp 1757982896
transform 1 0 82100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1157
timestamp 1757982896
transform 1 0 83600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1158
timestamp 1757982896
transform 1 0 85100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1159
timestamp 1757982896
transform 1 0 86600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1160
timestamp 1757982896
transform 1 0 88100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1161
timestamp 1757982896
transform 1 0 89600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1162
timestamp 1757982896
transform 1 0 91100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1163
timestamp 1757982896
transform 1 0 92600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1164
timestamp 1757982896
transform 1 0 94100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1165
timestamp 1757982896
transform 1 0 95600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1166
timestamp 1757982896
transform 1 0 97100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1167
timestamp 1757982896
transform 1 0 98600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1168
timestamp 1757982896
transform 1 0 100100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1169
timestamp 1757982896
transform 1 0 101600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1170
timestamp 1757982896
transform 1 0 103100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1171
timestamp 1757982896
transform 1 0 104600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1172
timestamp 1757982896
transform 1 0 106100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1173
timestamp 1757982896
transform 1 0 107600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1174
timestamp 1757982896
transform 1 0 109100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1175
timestamp 1757982896
transform 1 0 110600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1176
timestamp 1757982896
transform 1 0 112100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1177
timestamp 1757982896
transform 1 0 113600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1178
timestamp 1757982896
transform 1 0 115100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1179
timestamp 1757982896
transform 1 0 116600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1180
timestamp 1757982896
transform 1 0 118100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1181
timestamp 1757982896
transform 1 0 119600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1182
timestamp 1757982896
transform 1 0 121100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1183
timestamp 1757982896
transform 1 0 122600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1184
timestamp 1757982896
transform 1 0 124100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1185
timestamp 1757982896
transform 1 0 125600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1186
timestamp 1757982896
transform 1 0 127100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1187
timestamp 1757982896
transform 1 0 128600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1188
timestamp 1757982896
transform 1 0 130100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1189
timestamp 1757982896
transform 1 0 131600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1190
timestamp 1757982896
transform 1 0 133100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1191
timestamp 1757982896
transform 1 0 134600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1192
timestamp 1757982896
transform 1 0 136100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1193
timestamp 1757982896
transform 1 0 137600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1194
timestamp 1757982896
transform 1 0 139100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1195
timestamp 1757982896
transform 1 0 140600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1196
timestamp 1757982896
transform 1 0 142100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1197
timestamp 1757982896
transform 1 0 143600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1198
timestamp 1757982896
transform 1 0 145100 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1199
timestamp 1757982896
transform 1 0 146600 0 1 -15150
box 1820 -1430 3480 230
use pixel  pixel_1200
timestamp 1757982896
transform 1 0 -1900 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1201
timestamp 1757982896
transform 1 0 -400 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1202
timestamp 1757982896
transform 1 0 1100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1203
timestamp 1757982896
transform 1 0 2600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1204
timestamp 1757982896
transform 1 0 4100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1205
timestamp 1757982896
transform 1 0 5600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1206
timestamp 1757982896
transform 1 0 7100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1207
timestamp 1757982896
transform 1 0 8600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1208
timestamp 1757982896
transform 1 0 10100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1209
timestamp 1757982896
transform 1 0 11600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1210
timestamp 1757982896
transform 1 0 13100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1211
timestamp 1757982896
transform 1 0 14600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1212
timestamp 1757982896
transform 1 0 16100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1213
timestamp 1757982896
transform 1 0 17600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1214
timestamp 1757982896
transform 1 0 19100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1215
timestamp 1757982896
transform 1 0 20600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1216
timestamp 1757982896
transform 1 0 22100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1217
timestamp 1757982896
transform 1 0 23600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1218
timestamp 1757982896
transform 1 0 25100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1219
timestamp 1757982896
transform 1 0 26600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1220
timestamp 1757982896
transform 1 0 28100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1221
timestamp 1757982896
transform 1 0 29600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1222
timestamp 1757982896
transform 1 0 31100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1223
timestamp 1757982896
transform 1 0 32600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1224
timestamp 1757982896
transform 1 0 34100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1225
timestamp 1757982896
transform 1 0 35600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1226
timestamp 1757982896
transform 1 0 37100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1227
timestamp 1757982896
transform 1 0 38600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1228
timestamp 1757982896
transform 1 0 40100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1229
timestamp 1757982896
transform 1 0 41600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1230
timestamp 1757982896
transform 1 0 43100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1231
timestamp 1757982896
transform 1 0 44600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1232
timestamp 1757982896
transform 1 0 46100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1233
timestamp 1757982896
transform 1 0 47600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1234
timestamp 1757982896
transform 1 0 49100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1235
timestamp 1757982896
transform 1 0 50600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1236
timestamp 1757982896
transform 1 0 52100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1237
timestamp 1757982896
transform 1 0 53600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1238
timestamp 1757982896
transform 1 0 55100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1239
timestamp 1757982896
transform 1 0 56600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1240
timestamp 1757982896
transform 1 0 58100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1241
timestamp 1757982896
transform 1 0 59600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1242
timestamp 1757982896
transform 1 0 61100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1243
timestamp 1757982896
transform 1 0 62600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1244
timestamp 1757982896
transform 1 0 64100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1245
timestamp 1757982896
transform 1 0 65600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1246
timestamp 1757982896
transform 1 0 67100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1247
timestamp 1757982896
transform 1 0 68600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1248
timestamp 1757982896
transform 1 0 70100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1249
timestamp 1757982896
transform 1 0 71600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1250
timestamp 1757982896
transform 1 0 73100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1251
timestamp 1757982896
transform 1 0 74600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1252
timestamp 1757982896
transform 1 0 76100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1253
timestamp 1757982896
transform 1 0 77600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1254
timestamp 1757982896
transform 1 0 79100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1255
timestamp 1757982896
transform 1 0 80600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1256
timestamp 1757982896
transform 1 0 82100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1257
timestamp 1757982896
transform 1 0 83600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1258
timestamp 1757982896
transform 1 0 85100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1259
timestamp 1757982896
transform 1 0 86600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1260
timestamp 1757982896
transform 1 0 88100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1261
timestamp 1757982896
transform 1 0 89600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1262
timestamp 1757982896
transform 1 0 91100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1263
timestamp 1757982896
transform 1 0 92600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1264
timestamp 1757982896
transform 1 0 94100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1265
timestamp 1757982896
transform 1 0 95600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1266
timestamp 1757982896
transform 1 0 97100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1267
timestamp 1757982896
transform 1 0 98600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1268
timestamp 1757982896
transform 1 0 100100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1269
timestamp 1757982896
transform 1 0 101600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1270
timestamp 1757982896
transform 1 0 103100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1271
timestamp 1757982896
transform 1 0 104600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1272
timestamp 1757982896
transform 1 0 106100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1273
timestamp 1757982896
transform 1 0 107600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1274
timestamp 1757982896
transform 1 0 109100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1275
timestamp 1757982896
transform 1 0 110600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1276
timestamp 1757982896
transform 1 0 112100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1277
timestamp 1757982896
transform 1 0 113600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1278
timestamp 1757982896
transform 1 0 115100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1279
timestamp 1757982896
transform 1 0 116600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1280
timestamp 1757982896
transform 1 0 118100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1281
timestamp 1757982896
transform 1 0 119600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1282
timestamp 1757982896
transform 1 0 121100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1283
timestamp 1757982896
transform 1 0 122600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1284
timestamp 1757982896
transform 1 0 124100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1285
timestamp 1757982896
transform 1 0 125600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1286
timestamp 1757982896
transform 1 0 127100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1287
timestamp 1757982896
transform 1 0 128600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1288
timestamp 1757982896
transform 1 0 130100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1289
timestamp 1757982896
transform 1 0 131600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1290
timestamp 1757982896
transform 1 0 133100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1291
timestamp 1757982896
transform 1 0 134600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1292
timestamp 1757982896
transform 1 0 136100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1293
timestamp 1757982896
transform 1 0 137600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1294
timestamp 1757982896
transform 1 0 139100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1295
timestamp 1757982896
transform 1 0 140600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1296
timestamp 1757982896
transform 1 0 142100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1297
timestamp 1757982896
transform 1 0 143600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1298
timestamp 1757982896
transform 1 0 145100 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1299
timestamp 1757982896
transform 1 0 146600 0 1 -16650
box 1820 -1430 3480 230
use pixel  pixel_1300
timestamp 1757982896
transform 1 0 -1900 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1301
timestamp 1757982896
transform 1 0 -400 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1302
timestamp 1757982896
transform 1 0 1100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1303
timestamp 1757982896
transform 1 0 2600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1304
timestamp 1757982896
transform 1 0 4100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1305
timestamp 1757982896
transform 1 0 5600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1306
timestamp 1757982896
transform 1 0 7100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1307
timestamp 1757982896
transform 1 0 8600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1308
timestamp 1757982896
transform 1 0 10100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1309
timestamp 1757982896
transform 1 0 11600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1310
timestamp 1757982896
transform 1 0 13100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1311
timestamp 1757982896
transform 1 0 14600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1312
timestamp 1757982896
transform 1 0 16100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1313
timestamp 1757982896
transform 1 0 17600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1314
timestamp 1757982896
transform 1 0 19100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1315
timestamp 1757982896
transform 1 0 20600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1316
timestamp 1757982896
transform 1 0 22100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1317
timestamp 1757982896
transform 1 0 23600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1318
timestamp 1757982896
transform 1 0 25100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1319
timestamp 1757982896
transform 1 0 26600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1320
timestamp 1757982896
transform 1 0 28100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1321
timestamp 1757982896
transform 1 0 29600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1322
timestamp 1757982896
transform 1 0 31100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1323
timestamp 1757982896
transform 1 0 32600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1324
timestamp 1757982896
transform 1 0 34100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1325
timestamp 1757982896
transform 1 0 35600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1326
timestamp 1757982896
transform 1 0 37100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1327
timestamp 1757982896
transform 1 0 38600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1328
timestamp 1757982896
transform 1 0 40100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1329
timestamp 1757982896
transform 1 0 41600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1330
timestamp 1757982896
transform 1 0 43100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1331
timestamp 1757982896
transform 1 0 44600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1332
timestamp 1757982896
transform 1 0 46100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1333
timestamp 1757982896
transform 1 0 47600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1334
timestamp 1757982896
transform 1 0 49100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1335
timestamp 1757982896
transform 1 0 50600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1336
timestamp 1757982896
transform 1 0 52100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1337
timestamp 1757982896
transform 1 0 53600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1338
timestamp 1757982896
transform 1 0 55100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1339
timestamp 1757982896
transform 1 0 56600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1340
timestamp 1757982896
transform 1 0 58100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1341
timestamp 1757982896
transform 1 0 59600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1342
timestamp 1757982896
transform 1 0 61100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1343
timestamp 1757982896
transform 1 0 62600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1344
timestamp 1757982896
transform 1 0 64100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1345
timestamp 1757982896
transform 1 0 65600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1346
timestamp 1757982896
transform 1 0 67100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1347
timestamp 1757982896
transform 1 0 68600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1348
timestamp 1757982896
transform 1 0 70100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1349
timestamp 1757982896
transform 1 0 71600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1350
timestamp 1757982896
transform 1 0 73100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1351
timestamp 1757982896
transform 1 0 74600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1352
timestamp 1757982896
transform 1 0 76100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1353
timestamp 1757982896
transform 1 0 77600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1354
timestamp 1757982896
transform 1 0 79100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1355
timestamp 1757982896
transform 1 0 80600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1356
timestamp 1757982896
transform 1 0 82100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1357
timestamp 1757982896
transform 1 0 83600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1358
timestamp 1757982896
transform 1 0 85100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1359
timestamp 1757982896
transform 1 0 86600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1360
timestamp 1757982896
transform 1 0 88100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1361
timestamp 1757982896
transform 1 0 89600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1362
timestamp 1757982896
transform 1 0 91100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1363
timestamp 1757982896
transform 1 0 92600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1364
timestamp 1757982896
transform 1 0 94100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1365
timestamp 1757982896
transform 1 0 95600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1366
timestamp 1757982896
transform 1 0 97100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1367
timestamp 1757982896
transform 1 0 98600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1368
timestamp 1757982896
transform 1 0 100100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1369
timestamp 1757982896
transform 1 0 101600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1370
timestamp 1757982896
transform 1 0 103100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1371
timestamp 1757982896
transform 1 0 104600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1372
timestamp 1757982896
transform 1 0 106100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1373
timestamp 1757982896
transform 1 0 107600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1374
timestamp 1757982896
transform 1 0 109100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1375
timestamp 1757982896
transform 1 0 110600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1376
timestamp 1757982896
transform 1 0 112100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1377
timestamp 1757982896
transform 1 0 113600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1378
timestamp 1757982896
transform 1 0 115100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1379
timestamp 1757982896
transform 1 0 116600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1380
timestamp 1757982896
transform 1 0 118100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1381
timestamp 1757982896
transform 1 0 119600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1382
timestamp 1757982896
transform 1 0 121100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1383
timestamp 1757982896
transform 1 0 122600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1384
timestamp 1757982896
transform 1 0 124100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1385
timestamp 1757982896
transform 1 0 125600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1386
timestamp 1757982896
transform 1 0 127100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1387
timestamp 1757982896
transform 1 0 128600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1388
timestamp 1757982896
transform 1 0 130100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1389
timestamp 1757982896
transform 1 0 131600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1390
timestamp 1757982896
transform 1 0 133100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1391
timestamp 1757982896
transform 1 0 134600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1392
timestamp 1757982896
transform 1 0 136100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1393
timestamp 1757982896
transform 1 0 137600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1394
timestamp 1757982896
transform 1 0 139100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1395
timestamp 1757982896
transform 1 0 140600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1396
timestamp 1757982896
transform 1 0 142100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1397
timestamp 1757982896
transform 1 0 143600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1398
timestamp 1757982896
transform 1 0 145100 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1399
timestamp 1757982896
transform 1 0 146600 0 1 -18150
box 1820 -1430 3480 230
use pixel  pixel_1400
timestamp 1757982896
transform 1 0 -1900 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1401
timestamp 1757982896
transform 1 0 -400 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1402
timestamp 1757982896
transform 1 0 1100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1403
timestamp 1757982896
transform 1 0 2600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1404
timestamp 1757982896
transform 1 0 4100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1405
timestamp 1757982896
transform 1 0 5600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1406
timestamp 1757982896
transform 1 0 7100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1407
timestamp 1757982896
transform 1 0 8600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1408
timestamp 1757982896
transform 1 0 10100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1409
timestamp 1757982896
transform 1 0 11600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1410
timestamp 1757982896
transform 1 0 13100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1411
timestamp 1757982896
transform 1 0 14600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1412
timestamp 1757982896
transform 1 0 16100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1413
timestamp 1757982896
transform 1 0 17600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1414
timestamp 1757982896
transform 1 0 19100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1415
timestamp 1757982896
transform 1 0 20600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1416
timestamp 1757982896
transform 1 0 22100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1417
timestamp 1757982896
transform 1 0 23600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1418
timestamp 1757982896
transform 1 0 25100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1419
timestamp 1757982896
transform 1 0 26600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1420
timestamp 1757982896
transform 1 0 28100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1421
timestamp 1757982896
transform 1 0 29600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1422
timestamp 1757982896
transform 1 0 31100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1423
timestamp 1757982896
transform 1 0 32600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1424
timestamp 1757982896
transform 1 0 34100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1425
timestamp 1757982896
transform 1 0 35600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1426
timestamp 1757982896
transform 1 0 37100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1427
timestamp 1757982896
transform 1 0 38600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1428
timestamp 1757982896
transform 1 0 40100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1429
timestamp 1757982896
transform 1 0 41600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1430
timestamp 1757982896
transform 1 0 43100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1431
timestamp 1757982896
transform 1 0 44600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1432
timestamp 1757982896
transform 1 0 46100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1433
timestamp 1757982896
transform 1 0 47600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1434
timestamp 1757982896
transform 1 0 49100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1435
timestamp 1757982896
transform 1 0 50600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1436
timestamp 1757982896
transform 1 0 52100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1437
timestamp 1757982896
transform 1 0 53600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1438
timestamp 1757982896
transform 1 0 55100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1439
timestamp 1757982896
transform 1 0 56600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1440
timestamp 1757982896
transform 1 0 58100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1441
timestamp 1757982896
transform 1 0 59600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1442
timestamp 1757982896
transform 1 0 61100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1443
timestamp 1757982896
transform 1 0 62600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1444
timestamp 1757982896
transform 1 0 64100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1445
timestamp 1757982896
transform 1 0 65600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1446
timestamp 1757982896
transform 1 0 67100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1447
timestamp 1757982896
transform 1 0 68600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1448
timestamp 1757982896
transform 1 0 70100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1449
timestamp 1757982896
transform 1 0 71600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1450
timestamp 1757982896
transform 1 0 73100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1451
timestamp 1757982896
transform 1 0 74600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1452
timestamp 1757982896
transform 1 0 76100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1453
timestamp 1757982896
transform 1 0 77600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1454
timestamp 1757982896
transform 1 0 79100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1455
timestamp 1757982896
transform 1 0 80600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1456
timestamp 1757982896
transform 1 0 82100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1457
timestamp 1757982896
transform 1 0 83600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1458
timestamp 1757982896
transform 1 0 85100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1459
timestamp 1757982896
transform 1 0 86600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1460
timestamp 1757982896
transform 1 0 88100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1461
timestamp 1757982896
transform 1 0 89600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1462
timestamp 1757982896
transform 1 0 91100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1463
timestamp 1757982896
transform 1 0 92600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1464
timestamp 1757982896
transform 1 0 94100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1465
timestamp 1757982896
transform 1 0 95600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1466
timestamp 1757982896
transform 1 0 97100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1467
timestamp 1757982896
transform 1 0 98600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1468
timestamp 1757982896
transform 1 0 100100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1469
timestamp 1757982896
transform 1 0 101600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1470
timestamp 1757982896
transform 1 0 103100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1471
timestamp 1757982896
transform 1 0 104600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1472
timestamp 1757982896
transform 1 0 106100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1473
timestamp 1757982896
transform 1 0 107600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1474
timestamp 1757982896
transform 1 0 109100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1475
timestamp 1757982896
transform 1 0 110600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1476
timestamp 1757982896
transform 1 0 112100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1477
timestamp 1757982896
transform 1 0 113600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1478
timestamp 1757982896
transform 1 0 115100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1479
timestamp 1757982896
transform 1 0 116600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1480
timestamp 1757982896
transform 1 0 118100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1481
timestamp 1757982896
transform 1 0 119600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1482
timestamp 1757982896
transform 1 0 121100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1483
timestamp 1757982896
transform 1 0 122600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1484
timestamp 1757982896
transform 1 0 124100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1485
timestamp 1757982896
transform 1 0 125600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1486
timestamp 1757982896
transform 1 0 127100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1487
timestamp 1757982896
transform 1 0 128600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1488
timestamp 1757982896
transform 1 0 130100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1489
timestamp 1757982896
transform 1 0 131600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1490
timestamp 1757982896
transform 1 0 133100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1491
timestamp 1757982896
transform 1 0 134600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1492
timestamp 1757982896
transform 1 0 136100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1493
timestamp 1757982896
transform 1 0 137600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1494
timestamp 1757982896
transform 1 0 139100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1495
timestamp 1757982896
transform 1 0 140600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1496
timestamp 1757982896
transform 1 0 142100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1497
timestamp 1757982896
transform 1 0 143600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1498
timestamp 1757982896
transform 1 0 145100 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1499
timestamp 1757982896
transform 1 0 146600 0 1 -19650
box 1820 -1430 3480 230
use pixel  pixel_1500
timestamp 1757982896
transform 1 0 -1900 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1501
timestamp 1757982896
transform 1 0 -400 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1502
timestamp 1757982896
transform 1 0 1100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1503
timestamp 1757982896
transform 1 0 2600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1504
timestamp 1757982896
transform 1 0 4100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1505
timestamp 1757982896
transform 1 0 5600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1506
timestamp 1757982896
transform 1 0 7100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1507
timestamp 1757982896
transform 1 0 8600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1508
timestamp 1757982896
transform 1 0 10100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1509
timestamp 1757982896
transform 1 0 11600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1510
timestamp 1757982896
transform 1 0 13100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1511
timestamp 1757982896
transform 1 0 14600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1512
timestamp 1757982896
transform 1 0 16100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1513
timestamp 1757982896
transform 1 0 17600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1514
timestamp 1757982896
transform 1 0 19100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1515
timestamp 1757982896
transform 1 0 20600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1516
timestamp 1757982896
transform 1 0 22100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1517
timestamp 1757982896
transform 1 0 23600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1518
timestamp 1757982896
transform 1 0 25100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1519
timestamp 1757982896
transform 1 0 26600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1520
timestamp 1757982896
transform 1 0 28100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1521
timestamp 1757982896
transform 1 0 29600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1522
timestamp 1757982896
transform 1 0 31100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1523
timestamp 1757982896
transform 1 0 32600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1524
timestamp 1757982896
transform 1 0 34100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1525
timestamp 1757982896
transform 1 0 35600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1526
timestamp 1757982896
transform 1 0 37100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1527
timestamp 1757982896
transform 1 0 38600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1528
timestamp 1757982896
transform 1 0 40100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1529
timestamp 1757982896
transform 1 0 41600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1530
timestamp 1757982896
transform 1 0 43100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1531
timestamp 1757982896
transform 1 0 44600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1532
timestamp 1757982896
transform 1 0 46100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1533
timestamp 1757982896
transform 1 0 47600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1534
timestamp 1757982896
transform 1 0 49100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1535
timestamp 1757982896
transform 1 0 50600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1536
timestamp 1757982896
transform 1 0 52100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1537
timestamp 1757982896
transform 1 0 53600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1538
timestamp 1757982896
transform 1 0 55100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1539
timestamp 1757982896
transform 1 0 56600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1540
timestamp 1757982896
transform 1 0 58100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1541
timestamp 1757982896
transform 1 0 59600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1542
timestamp 1757982896
transform 1 0 61100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1543
timestamp 1757982896
transform 1 0 62600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1544
timestamp 1757982896
transform 1 0 64100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1545
timestamp 1757982896
transform 1 0 65600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1546
timestamp 1757982896
transform 1 0 67100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1547
timestamp 1757982896
transform 1 0 68600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1548
timestamp 1757982896
transform 1 0 70100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1549
timestamp 1757982896
transform 1 0 71600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1550
timestamp 1757982896
transform 1 0 73100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1551
timestamp 1757982896
transform 1 0 74600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1552
timestamp 1757982896
transform 1 0 76100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1553
timestamp 1757982896
transform 1 0 77600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1554
timestamp 1757982896
transform 1 0 79100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1555
timestamp 1757982896
transform 1 0 80600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1556
timestamp 1757982896
transform 1 0 82100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1557
timestamp 1757982896
transform 1 0 83600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1558
timestamp 1757982896
transform 1 0 85100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1559
timestamp 1757982896
transform 1 0 86600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1560
timestamp 1757982896
transform 1 0 88100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1561
timestamp 1757982896
transform 1 0 89600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1562
timestamp 1757982896
transform 1 0 91100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1563
timestamp 1757982896
transform 1 0 92600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1564
timestamp 1757982896
transform 1 0 94100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1565
timestamp 1757982896
transform 1 0 95600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1566
timestamp 1757982896
transform 1 0 97100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1567
timestamp 1757982896
transform 1 0 98600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1568
timestamp 1757982896
transform 1 0 100100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1569
timestamp 1757982896
transform 1 0 101600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1570
timestamp 1757982896
transform 1 0 103100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1571
timestamp 1757982896
transform 1 0 104600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1572
timestamp 1757982896
transform 1 0 106100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1573
timestamp 1757982896
transform 1 0 107600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1574
timestamp 1757982896
transform 1 0 109100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1575
timestamp 1757982896
transform 1 0 110600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1576
timestamp 1757982896
transform 1 0 112100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1577
timestamp 1757982896
transform 1 0 113600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1578
timestamp 1757982896
transform 1 0 115100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1579
timestamp 1757982896
transform 1 0 116600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1580
timestamp 1757982896
transform 1 0 118100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1581
timestamp 1757982896
transform 1 0 119600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1582
timestamp 1757982896
transform 1 0 121100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1583
timestamp 1757982896
transform 1 0 122600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1584
timestamp 1757982896
transform 1 0 124100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1585
timestamp 1757982896
transform 1 0 125600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1586
timestamp 1757982896
transform 1 0 127100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1587
timestamp 1757982896
transform 1 0 128600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1588
timestamp 1757982896
transform 1 0 130100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1589
timestamp 1757982896
transform 1 0 131600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1590
timestamp 1757982896
transform 1 0 133100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1591
timestamp 1757982896
transform 1 0 134600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1592
timestamp 1757982896
transform 1 0 136100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1593
timestamp 1757982896
transform 1 0 137600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1594
timestamp 1757982896
transform 1 0 139100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1595
timestamp 1757982896
transform 1 0 140600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1596
timestamp 1757982896
transform 1 0 142100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1597
timestamp 1757982896
transform 1 0 143600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1598
timestamp 1757982896
transform 1 0 145100 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1599
timestamp 1757982896
transform 1 0 146600 0 1 -21150
box 1820 -1430 3480 230
use pixel  pixel_1600
timestamp 1757982896
transform 1 0 -1900 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1601
timestamp 1757982896
transform 1 0 -400 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1602
timestamp 1757982896
transform 1 0 1100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1603
timestamp 1757982896
transform 1 0 2600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1604
timestamp 1757982896
transform 1 0 4100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1605
timestamp 1757982896
transform 1 0 5600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1606
timestamp 1757982896
transform 1 0 7100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1607
timestamp 1757982896
transform 1 0 8600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1608
timestamp 1757982896
transform 1 0 10100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1609
timestamp 1757982896
transform 1 0 11600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1610
timestamp 1757982896
transform 1 0 13100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1611
timestamp 1757982896
transform 1 0 14600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1612
timestamp 1757982896
transform 1 0 16100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1613
timestamp 1757982896
transform 1 0 17600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1614
timestamp 1757982896
transform 1 0 19100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1615
timestamp 1757982896
transform 1 0 20600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1616
timestamp 1757982896
transform 1 0 22100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1617
timestamp 1757982896
transform 1 0 23600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1618
timestamp 1757982896
transform 1 0 25100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1619
timestamp 1757982896
transform 1 0 26600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1620
timestamp 1757982896
transform 1 0 28100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1621
timestamp 1757982896
transform 1 0 29600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1622
timestamp 1757982896
transform 1 0 31100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1623
timestamp 1757982896
transform 1 0 32600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1624
timestamp 1757982896
transform 1 0 34100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1625
timestamp 1757982896
transform 1 0 35600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1626
timestamp 1757982896
transform 1 0 37100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1627
timestamp 1757982896
transform 1 0 38600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1628
timestamp 1757982896
transform 1 0 40100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1629
timestamp 1757982896
transform 1 0 41600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1630
timestamp 1757982896
transform 1 0 43100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1631
timestamp 1757982896
transform 1 0 44600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1632
timestamp 1757982896
transform 1 0 46100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1633
timestamp 1757982896
transform 1 0 47600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1634
timestamp 1757982896
transform 1 0 49100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1635
timestamp 1757982896
transform 1 0 50600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1636
timestamp 1757982896
transform 1 0 52100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1637
timestamp 1757982896
transform 1 0 53600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1638
timestamp 1757982896
transform 1 0 55100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1639
timestamp 1757982896
transform 1 0 56600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1640
timestamp 1757982896
transform 1 0 58100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1641
timestamp 1757982896
transform 1 0 59600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1642
timestamp 1757982896
transform 1 0 61100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1643
timestamp 1757982896
transform 1 0 62600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1644
timestamp 1757982896
transform 1 0 64100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1645
timestamp 1757982896
transform 1 0 65600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1646
timestamp 1757982896
transform 1 0 67100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1647
timestamp 1757982896
transform 1 0 68600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1648
timestamp 1757982896
transform 1 0 70100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1649
timestamp 1757982896
transform 1 0 71600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1650
timestamp 1757982896
transform 1 0 73100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1651
timestamp 1757982896
transform 1 0 74600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1652
timestamp 1757982896
transform 1 0 76100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1653
timestamp 1757982896
transform 1 0 77600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1654
timestamp 1757982896
transform 1 0 79100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1655
timestamp 1757982896
transform 1 0 80600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1656
timestamp 1757982896
transform 1 0 82100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1657
timestamp 1757982896
transform 1 0 83600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1658
timestamp 1757982896
transform 1 0 85100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1659
timestamp 1757982896
transform 1 0 86600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1660
timestamp 1757982896
transform 1 0 88100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1661
timestamp 1757982896
transform 1 0 89600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1662
timestamp 1757982896
transform 1 0 91100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1663
timestamp 1757982896
transform 1 0 92600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1664
timestamp 1757982896
transform 1 0 94100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1665
timestamp 1757982896
transform 1 0 95600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1666
timestamp 1757982896
transform 1 0 97100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1667
timestamp 1757982896
transform 1 0 98600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1668
timestamp 1757982896
transform 1 0 100100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1669
timestamp 1757982896
transform 1 0 101600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1670
timestamp 1757982896
transform 1 0 103100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1671
timestamp 1757982896
transform 1 0 104600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1672
timestamp 1757982896
transform 1 0 106100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1673
timestamp 1757982896
transform 1 0 107600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1674
timestamp 1757982896
transform 1 0 109100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1675
timestamp 1757982896
transform 1 0 110600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1676
timestamp 1757982896
transform 1 0 112100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1677
timestamp 1757982896
transform 1 0 113600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1678
timestamp 1757982896
transform 1 0 115100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1679
timestamp 1757982896
transform 1 0 116600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1680
timestamp 1757982896
transform 1 0 118100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1681
timestamp 1757982896
transform 1 0 119600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1682
timestamp 1757982896
transform 1 0 121100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1683
timestamp 1757982896
transform 1 0 122600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1684
timestamp 1757982896
transform 1 0 124100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1685
timestamp 1757982896
transform 1 0 125600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1686
timestamp 1757982896
transform 1 0 127100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1687
timestamp 1757982896
transform 1 0 128600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1688
timestamp 1757982896
transform 1 0 130100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1689
timestamp 1757982896
transform 1 0 131600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1690
timestamp 1757982896
transform 1 0 133100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1691
timestamp 1757982896
transform 1 0 134600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1692
timestamp 1757982896
transform 1 0 136100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1693
timestamp 1757982896
transform 1 0 137600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1694
timestamp 1757982896
transform 1 0 139100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1695
timestamp 1757982896
transform 1 0 140600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1696
timestamp 1757982896
transform 1 0 142100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1697
timestamp 1757982896
transform 1 0 143600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1698
timestamp 1757982896
transform 1 0 145100 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1699
timestamp 1757982896
transform 1 0 146600 0 1 -22650
box 1820 -1430 3480 230
use pixel  pixel_1700
timestamp 1757982896
transform 1 0 -1900 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1701
timestamp 1757982896
transform 1 0 -400 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1702
timestamp 1757982896
transform 1 0 1100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1703
timestamp 1757982896
transform 1 0 2600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1704
timestamp 1757982896
transform 1 0 4100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1705
timestamp 1757982896
transform 1 0 5600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1706
timestamp 1757982896
transform 1 0 7100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1707
timestamp 1757982896
transform 1 0 8600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1708
timestamp 1757982896
transform 1 0 10100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1709
timestamp 1757982896
transform 1 0 11600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1710
timestamp 1757982896
transform 1 0 13100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1711
timestamp 1757982896
transform 1 0 14600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1712
timestamp 1757982896
transform 1 0 16100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1713
timestamp 1757982896
transform 1 0 17600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1714
timestamp 1757982896
transform 1 0 19100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1715
timestamp 1757982896
transform 1 0 20600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1716
timestamp 1757982896
transform 1 0 22100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1717
timestamp 1757982896
transform 1 0 23600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1718
timestamp 1757982896
transform 1 0 25100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1719
timestamp 1757982896
transform 1 0 26600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1720
timestamp 1757982896
transform 1 0 28100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1721
timestamp 1757982896
transform 1 0 29600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1722
timestamp 1757982896
transform 1 0 31100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1723
timestamp 1757982896
transform 1 0 32600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1724
timestamp 1757982896
transform 1 0 34100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1725
timestamp 1757982896
transform 1 0 35600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1726
timestamp 1757982896
transform 1 0 37100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1727
timestamp 1757982896
transform 1 0 38600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1728
timestamp 1757982896
transform 1 0 40100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1729
timestamp 1757982896
transform 1 0 41600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1730
timestamp 1757982896
transform 1 0 43100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1731
timestamp 1757982896
transform 1 0 44600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1732
timestamp 1757982896
transform 1 0 46100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1733
timestamp 1757982896
transform 1 0 47600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1734
timestamp 1757982896
transform 1 0 49100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1735
timestamp 1757982896
transform 1 0 50600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1736
timestamp 1757982896
transform 1 0 52100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1737
timestamp 1757982896
transform 1 0 53600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1738
timestamp 1757982896
transform 1 0 55100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1739
timestamp 1757982896
transform 1 0 56600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1740
timestamp 1757982896
transform 1 0 58100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1741
timestamp 1757982896
transform 1 0 59600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1742
timestamp 1757982896
transform 1 0 61100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1743
timestamp 1757982896
transform 1 0 62600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1744
timestamp 1757982896
transform 1 0 64100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1745
timestamp 1757982896
transform 1 0 65600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1746
timestamp 1757982896
transform 1 0 67100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1747
timestamp 1757982896
transform 1 0 68600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1748
timestamp 1757982896
transform 1 0 70100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1749
timestamp 1757982896
transform 1 0 71600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1750
timestamp 1757982896
transform 1 0 73100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1751
timestamp 1757982896
transform 1 0 74600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1752
timestamp 1757982896
transform 1 0 76100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1753
timestamp 1757982896
transform 1 0 77600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1754
timestamp 1757982896
transform 1 0 79100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1755
timestamp 1757982896
transform 1 0 80600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1756
timestamp 1757982896
transform 1 0 82100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1757
timestamp 1757982896
transform 1 0 83600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1758
timestamp 1757982896
transform 1 0 85100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1759
timestamp 1757982896
transform 1 0 86600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1760
timestamp 1757982896
transform 1 0 88100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1761
timestamp 1757982896
transform 1 0 89600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1762
timestamp 1757982896
transform 1 0 91100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1763
timestamp 1757982896
transform 1 0 92600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1764
timestamp 1757982896
transform 1 0 94100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1765
timestamp 1757982896
transform 1 0 95600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1766
timestamp 1757982896
transform 1 0 97100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1767
timestamp 1757982896
transform 1 0 98600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1768
timestamp 1757982896
transform 1 0 100100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1769
timestamp 1757982896
transform 1 0 101600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1770
timestamp 1757982896
transform 1 0 103100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1771
timestamp 1757982896
transform 1 0 104600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1772
timestamp 1757982896
transform 1 0 106100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1773
timestamp 1757982896
transform 1 0 107600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1774
timestamp 1757982896
transform 1 0 109100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1775
timestamp 1757982896
transform 1 0 110600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1776
timestamp 1757982896
transform 1 0 112100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1777
timestamp 1757982896
transform 1 0 113600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1778
timestamp 1757982896
transform 1 0 115100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1779
timestamp 1757982896
transform 1 0 116600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1780
timestamp 1757982896
transform 1 0 118100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1781
timestamp 1757982896
transform 1 0 119600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1782
timestamp 1757982896
transform 1 0 121100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1783
timestamp 1757982896
transform 1 0 122600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1784
timestamp 1757982896
transform 1 0 124100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1785
timestamp 1757982896
transform 1 0 125600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1786
timestamp 1757982896
transform 1 0 127100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1787
timestamp 1757982896
transform 1 0 128600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1788
timestamp 1757982896
transform 1 0 130100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1789
timestamp 1757982896
transform 1 0 131600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1790
timestamp 1757982896
transform 1 0 133100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1791
timestamp 1757982896
transform 1 0 134600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1792
timestamp 1757982896
transform 1 0 136100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1793
timestamp 1757982896
transform 1 0 137600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1794
timestamp 1757982896
transform 1 0 139100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1795
timestamp 1757982896
transform 1 0 140600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1796
timestamp 1757982896
transform 1 0 142100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1797
timestamp 1757982896
transform 1 0 143600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1798
timestamp 1757982896
transform 1 0 145100 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1799
timestamp 1757982896
transform 1 0 146600 0 1 -24150
box 1820 -1430 3480 230
use pixel  pixel_1800
timestamp 1757982896
transform 1 0 -1900 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1801
timestamp 1757982896
transform 1 0 -400 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1802
timestamp 1757982896
transform 1 0 1100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1803
timestamp 1757982896
transform 1 0 2600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1804
timestamp 1757982896
transform 1 0 4100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1805
timestamp 1757982896
transform 1 0 5600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1806
timestamp 1757982896
transform 1 0 7100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1807
timestamp 1757982896
transform 1 0 8600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1808
timestamp 1757982896
transform 1 0 10100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1809
timestamp 1757982896
transform 1 0 11600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1810
timestamp 1757982896
transform 1 0 13100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1811
timestamp 1757982896
transform 1 0 14600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1812
timestamp 1757982896
transform 1 0 16100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1813
timestamp 1757982896
transform 1 0 17600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1814
timestamp 1757982896
transform 1 0 19100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1815
timestamp 1757982896
transform 1 0 20600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1816
timestamp 1757982896
transform 1 0 22100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1817
timestamp 1757982896
transform 1 0 23600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1818
timestamp 1757982896
transform 1 0 25100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1819
timestamp 1757982896
transform 1 0 26600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1820
timestamp 1757982896
transform 1 0 28100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1821
timestamp 1757982896
transform 1 0 29600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1822
timestamp 1757982896
transform 1 0 31100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1823
timestamp 1757982896
transform 1 0 32600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1824
timestamp 1757982896
transform 1 0 34100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1825
timestamp 1757982896
transform 1 0 35600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1826
timestamp 1757982896
transform 1 0 37100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1827
timestamp 1757982896
transform 1 0 38600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1828
timestamp 1757982896
transform 1 0 40100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1829
timestamp 1757982896
transform 1 0 41600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1830
timestamp 1757982896
transform 1 0 43100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1831
timestamp 1757982896
transform 1 0 44600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1832
timestamp 1757982896
transform 1 0 46100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1833
timestamp 1757982896
transform 1 0 47600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1834
timestamp 1757982896
transform 1 0 49100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1835
timestamp 1757982896
transform 1 0 50600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1836
timestamp 1757982896
transform 1 0 52100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1837
timestamp 1757982896
transform 1 0 53600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1838
timestamp 1757982896
transform 1 0 55100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1839
timestamp 1757982896
transform 1 0 56600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1840
timestamp 1757982896
transform 1 0 58100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1841
timestamp 1757982896
transform 1 0 59600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1842
timestamp 1757982896
transform 1 0 61100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1843
timestamp 1757982896
transform 1 0 62600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1844
timestamp 1757982896
transform 1 0 64100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1845
timestamp 1757982896
transform 1 0 65600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1846
timestamp 1757982896
transform 1 0 67100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1847
timestamp 1757982896
transform 1 0 68600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1848
timestamp 1757982896
transform 1 0 70100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1849
timestamp 1757982896
transform 1 0 71600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1850
timestamp 1757982896
transform 1 0 73100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1851
timestamp 1757982896
transform 1 0 74600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1852
timestamp 1757982896
transform 1 0 76100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1853
timestamp 1757982896
transform 1 0 77600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1854
timestamp 1757982896
transform 1 0 79100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1855
timestamp 1757982896
transform 1 0 80600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1856
timestamp 1757982896
transform 1 0 82100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1857
timestamp 1757982896
transform 1 0 83600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1858
timestamp 1757982896
transform 1 0 85100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1859
timestamp 1757982896
transform 1 0 86600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1860
timestamp 1757982896
transform 1 0 88100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1861
timestamp 1757982896
transform 1 0 89600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1862
timestamp 1757982896
transform 1 0 91100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1863
timestamp 1757982896
transform 1 0 92600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1864
timestamp 1757982896
transform 1 0 94100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1865
timestamp 1757982896
transform 1 0 95600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1866
timestamp 1757982896
transform 1 0 97100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1867
timestamp 1757982896
transform 1 0 98600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1868
timestamp 1757982896
transform 1 0 100100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1869
timestamp 1757982896
transform 1 0 101600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1870
timestamp 1757982896
transform 1 0 103100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1871
timestamp 1757982896
transform 1 0 104600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1872
timestamp 1757982896
transform 1 0 106100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1873
timestamp 1757982896
transform 1 0 107600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1874
timestamp 1757982896
transform 1 0 109100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1875
timestamp 1757982896
transform 1 0 110600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1876
timestamp 1757982896
transform 1 0 112100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1877
timestamp 1757982896
transform 1 0 113600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1878
timestamp 1757982896
transform 1 0 115100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1879
timestamp 1757982896
transform 1 0 116600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1880
timestamp 1757982896
transform 1 0 118100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1881
timestamp 1757982896
transform 1 0 119600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1882
timestamp 1757982896
transform 1 0 121100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1883
timestamp 1757982896
transform 1 0 122600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1884
timestamp 1757982896
transform 1 0 124100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1885
timestamp 1757982896
transform 1 0 125600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1886
timestamp 1757982896
transform 1 0 127100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1887
timestamp 1757982896
transform 1 0 128600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1888
timestamp 1757982896
transform 1 0 130100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1889
timestamp 1757982896
transform 1 0 131600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1890
timestamp 1757982896
transform 1 0 133100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1891
timestamp 1757982896
transform 1 0 134600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1892
timestamp 1757982896
transform 1 0 136100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1893
timestamp 1757982896
transform 1 0 137600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1894
timestamp 1757982896
transform 1 0 139100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1895
timestamp 1757982896
transform 1 0 140600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1896
timestamp 1757982896
transform 1 0 142100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1897
timestamp 1757982896
transform 1 0 143600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1898
timestamp 1757982896
transform 1 0 145100 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1899
timestamp 1757982896
transform 1 0 146600 0 1 -25650
box 1820 -1430 3480 230
use pixel  pixel_1900
timestamp 1757982896
transform 1 0 -1900 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1901
timestamp 1757982896
transform 1 0 -400 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1902
timestamp 1757982896
transform 1 0 1100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1903
timestamp 1757982896
transform 1 0 2600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1904
timestamp 1757982896
transform 1 0 4100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1905
timestamp 1757982896
transform 1 0 5600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1906
timestamp 1757982896
transform 1 0 7100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1907
timestamp 1757982896
transform 1 0 8600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1908
timestamp 1757982896
transform 1 0 10100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1909
timestamp 1757982896
transform 1 0 11600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1910
timestamp 1757982896
transform 1 0 13100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1911
timestamp 1757982896
transform 1 0 14600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1912
timestamp 1757982896
transform 1 0 16100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1913
timestamp 1757982896
transform 1 0 17600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1914
timestamp 1757982896
transform 1 0 19100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1915
timestamp 1757982896
transform 1 0 20600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1916
timestamp 1757982896
transform 1 0 22100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1917
timestamp 1757982896
transform 1 0 23600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1918
timestamp 1757982896
transform 1 0 25100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1919
timestamp 1757982896
transform 1 0 26600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1920
timestamp 1757982896
transform 1 0 28100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1921
timestamp 1757982896
transform 1 0 29600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1922
timestamp 1757982896
transform 1 0 31100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1923
timestamp 1757982896
transform 1 0 32600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1924
timestamp 1757982896
transform 1 0 34100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1925
timestamp 1757982896
transform 1 0 35600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1926
timestamp 1757982896
transform 1 0 37100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1927
timestamp 1757982896
transform 1 0 38600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1928
timestamp 1757982896
transform 1 0 40100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1929
timestamp 1757982896
transform 1 0 41600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1930
timestamp 1757982896
transform 1 0 43100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1931
timestamp 1757982896
transform 1 0 44600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1932
timestamp 1757982896
transform 1 0 46100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1933
timestamp 1757982896
transform 1 0 47600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1934
timestamp 1757982896
transform 1 0 49100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1935
timestamp 1757982896
transform 1 0 50600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1936
timestamp 1757982896
transform 1 0 52100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1937
timestamp 1757982896
transform 1 0 53600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1938
timestamp 1757982896
transform 1 0 55100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1939
timestamp 1757982896
transform 1 0 56600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1940
timestamp 1757982896
transform 1 0 58100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1941
timestamp 1757982896
transform 1 0 59600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1942
timestamp 1757982896
transform 1 0 61100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1943
timestamp 1757982896
transform 1 0 62600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1944
timestamp 1757982896
transform 1 0 64100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1945
timestamp 1757982896
transform 1 0 65600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1946
timestamp 1757982896
transform 1 0 67100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1947
timestamp 1757982896
transform 1 0 68600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1948
timestamp 1757982896
transform 1 0 70100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1949
timestamp 1757982896
transform 1 0 71600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1950
timestamp 1757982896
transform 1 0 73100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1951
timestamp 1757982896
transform 1 0 74600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1952
timestamp 1757982896
transform 1 0 76100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1953
timestamp 1757982896
transform 1 0 77600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1954
timestamp 1757982896
transform 1 0 79100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1955
timestamp 1757982896
transform 1 0 80600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1956
timestamp 1757982896
transform 1 0 82100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1957
timestamp 1757982896
transform 1 0 83600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1958
timestamp 1757982896
transform 1 0 85100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1959
timestamp 1757982896
transform 1 0 86600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1960
timestamp 1757982896
transform 1 0 88100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1961
timestamp 1757982896
transform 1 0 89600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1962
timestamp 1757982896
transform 1 0 91100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1963
timestamp 1757982896
transform 1 0 92600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1964
timestamp 1757982896
transform 1 0 94100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1965
timestamp 1757982896
transform 1 0 95600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1966
timestamp 1757982896
transform 1 0 97100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1967
timestamp 1757982896
transform 1 0 98600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1968
timestamp 1757982896
transform 1 0 100100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1969
timestamp 1757982896
transform 1 0 101600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1970
timestamp 1757982896
transform 1 0 103100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1971
timestamp 1757982896
transform 1 0 104600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1972
timestamp 1757982896
transform 1 0 106100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1973
timestamp 1757982896
transform 1 0 107600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1974
timestamp 1757982896
transform 1 0 109100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1975
timestamp 1757982896
transform 1 0 110600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1976
timestamp 1757982896
transform 1 0 112100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1977
timestamp 1757982896
transform 1 0 113600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1978
timestamp 1757982896
transform 1 0 115100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1979
timestamp 1757982896
transform 1 0 116600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1980
timestamp 1757982896
transform 1 0 118100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1981
timestamp 1757982896
transform 1 0 119600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1982
timestamp 1757982896
transform 1 0 121100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1983
timestamp 1757982896
transform 1 0 122600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1984
timestamp 1757982896
transform 1 0 124100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1985
timestamp 1757982896
transform 1 0 125600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1986
timestamp 1757982896
transform 1 0 127100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1987
timestamp 1757982896
transform 1 0 128600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1988
timestamp 1757982896
transform 1 0 130100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1989
timestamp 1757982896
transform 1 0 131600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1990
timestamp 1757982896
transform 1 0 133100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1991
timestamp 1757982896
transform 1 0 134600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1992
timestamp 1757982896
transform 1 0 136100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1993
timestamp 1757982896
transform 1 0 137600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1994
timestamp 1757982896
transform 1 0 139100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1995
timestamp 1757982896
transform 1 0 140600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1996
timestamp 1757982896
transform 1 0 142100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1997
timestamp 1757982896
transform 1 0 143600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1998
timestamp 1757982896
transform 1 0 145100 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_1999
timestamp 1757982896
transform 1 0 146600 0 1 -27150
box 1820 -1430 3480 230
use pixel  pixel_2000
timestamp 1757982896
transform 1 0 -1900 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2001
timestamp 1757982896
transform 1 0 -400 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2002
timestamp 1757982896
transform 1 0 1100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2003
timestamp 1757982896
transform 1 0 2600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2004
timestamp 1757982896
transform 1 0 4100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2005
timestamp 1757982896
transform 1 0 5600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2006
timestamp 1757982896
transform 1 0 7100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2007
timestamp 1757982896
transform 1 0 8600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2008
timestamp 1757982896
transform 1 0 10100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2009
timestamp 1757982896
transform 1 0 11600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2010
timestamp 1757982896
transform 1 0 13100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2011
timestamp 1757982896
transform 1 0 14600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2012
timestamp 1757982896
transform 1 0 16100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2013
timestamp 1757982896
transform 1 0 17600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2014
timestamp 1757982896
transform 1 0 19100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2015
timestamp 1757982896
transform 1 0 20600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2016
timestamp 1757982896
transform 1 0 22100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2017
timestamp 1757982896
transform 1 0 23600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2018
timestamp 1757982896
transform 1 0 25100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2019
timestamp 1757982896
transform 1 0 26600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2020
timestamp 1757982896
transform 1 0 28100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2021
timestamp 1757982896
transform 1 0 29600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2022
timestamp 1757982896
transform 1 0 31100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2023
timestamp 1757982896
transform 1 0 32600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2024
timestamp 1757982896
transform 1 0 34100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2025
timestamp 1757982896
transform 1 0 35600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2026
timestamp 1757982896
transform 1 0 37100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2027
timestamp 1757982896
transform 1 0 38600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2028
timestamp 1757982896
transform 1 0 40100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2029
timestamp 1757982896
transform 1 0 41600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2030
timestamp 1757982896
transform 1 0 43100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2031
timestamp 1757982896
transform 1 0 44600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2032
timestamp 1757982896
transform 1 0 46100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2033
timestamp 1757982896
transform 1 0 47600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2034
timestamp 1757982896
transform 1 0 49100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2035
timestamp 1757982896
transform 1 0 50600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2036
timestamp 1757982896
transform 1 0 52100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2037
timestamp 1757982896
transform 1 0 53600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2038
timestamp 1757982896
transform 1 0 55100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2039
timestamp 1757982896
transform 1 0 56600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2040
timestamp 1757982896
transform 1 0 58100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2041
timestamp 1757982896
transform 1 0 59600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2042
timestamp 1757982896
transform 1 0 61100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2043
timestamp 1757982896
transform 1 0 62600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2044
timestamp 1757982896
transform 1 0 64100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2045
timestamp 1757982896
transform 1 0 65600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2046
timestamp 1757982896
transform 1 0 67100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2047
timestamp 1757982896
transform 1 0 68600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2048
timestamp 1757982896
transform 1 0 70100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2049
timestamp 1757982896
transform 1 0 71600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2050
timestamp 1757982896
transform 1 0 73100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2051
timestamp 1757982896
transform 1 0 74600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2052
timestamp 1757982896
transform 1 0 76100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2053
timestamp 1757982896
transform 1 0 77600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2054
timestamp 1757982896
transform 1 0 79100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2055
timestamp 1757982896
transform 1 0 80600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2056
timestamp 1757982896
transform 1 0 82100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2057
timestamp 1757982896
transform 1 0 83600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2058
timestamp 1757982896
transform 1 0 85100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2059
timestamp 1757982896
transform 1 0 86600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2060
timestamp 1757982896
transform 1 0 88100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2061
timestamp 1757982896
transform 1 0 89600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2062
timestamp 1757982896
transform 1 0 91100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2063
timestamp 1757982896
transform 1 0 92600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2064
timestamp 1757982896
transform 1 0 94100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2065
timestamp 1757982896
transform 1 0 95600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2066
timestamp 1757982896
transform 1 0 97100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2067
timestamp 1757982896
transform 1 0 98600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2068
timestamp 1757982896
transform 1 0 100100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2069
timestamp 1757982896
transform 1 0 101600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2070
timestamp 1757982896
transform 1 0 103100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2071
timestamp 1757982896
transform 1 0 104600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2072
timestamp 1757982896
transform 1 0 106100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2073
timestamp 1757982896
transform 1 0 107600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2074
timestamp 1757982896
transform 1 0 109100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2075
timestamp 1757982896
transform 1 0 110600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2076
timestamp 1757982896
transform 1 0 112100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2077
timestamp 1757982896
transform 1 0 113600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2078
timestamp 1757982896
transform 1 0 115100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2079
timestamp 1757982896
transform 1 0 116600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2080
timestamp 1757982896
transform 1 0 118100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2081
timestamp 1757982896
transform 1 0 119600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2082
timestamp 1757982896
transform 1 0 121100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2083
timestamp 1757982896
transform 1 0 122600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2084
timestamp 1757982896
transform 1 0 124100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2085
timestamp 1757982896
transform 1 0 125600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2086
timestamp 1757982896
transform 1 0 127100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2087
timestamp 1757982896
transform 1 0 128600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2088
timestamp 1757982896
transform 1 0 130100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2089
timestamp 1757982896
transform 1 0 131600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2090
timestamp 1757982896
transform 1 0 133100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2091
timestamp 1757982896
transform 1 0 134600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2092
timestamp 1757982896
transform 1 0 136100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2093
timestamp 1757982896
transform 1 0 137600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2094
timestamp 1757982896
transform 1 0 139100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2095
timestamp 1757982896
transform 1 0 140600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2096
timestamp 1757982896
transform 1 0 142100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2097
timestamp 1757982896
transform 1 0 143600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2098
timestamp 1757982896
transform 1 0 145100 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2099
timestamp 1757982896
transform 1 0 146600 0 1 -28650
box 1820 -1430 3480 230
use pixel  pixel_2100
timestamp 1757982896
transform 1 0 -1900 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2101
timestamp 1757982896
transform 1 0 -400 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2102
timestamp 1757982896
transform 1 0 1100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2103
timestamp 1757982896
transform 1 0 2600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2104
timestamp 1757982896
transform 1 0 4100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2105
timestamp 1757982896
transform 1 0 5600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2106
timestamp 1757982896
transform 1 0 7100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2107
timestamp 1757982896
transform 1 0 8600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2108
timestamp 1757982896
transform 1 0 10100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2109
timestamp 1757982896
transform 1 0 11600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2110
timestamp 1757982896
transform 1 0 13100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2111
timestamp 1757982896
transform 1 0 14600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2112
timestamp 1757982896
transform 1 0 16100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2113
timestamp 1757982896
transform 1 0 17600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2114
timestamp 1757982896
transform 1 0 19100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2115
timestamp 1757982896
transform 1 0 20600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2116
timestamp 1757982896
transform 1 0 22100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2117
timestamp 1757982896
transform 1 0 23600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2118
timestamp 1757982896
transform 1 0 25100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2119
timestamp 1757982896
transform 1 0 26600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2120
timestamp 1757982896
transform 1 0 28100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2121
timestamp 1757982896
transform 1 0 29600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2122
timestamp 1757982896
transform 1 0 31100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2123
timestamp 1757982896
transform 1 0 32600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2124
timestamp 1757982896
transform 1 0 34100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2125
timestamp 1757982896
transform 1 0 35600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2126
timestamp 1757982896
transform 1 0 37100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2127
timestamp 1757982896
transform 1 0 38600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2128
timestamp 1757982896
transform 1 0 40100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2129
timestamp 1757982896
transform 1 0 41600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2130
timestamp 1757982896
transform 1 0 43100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2131
timestamp 1757982896
transform 1 0 44600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2132
timestamp 1757982896
transform 1 0 46100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2133
timestamp 1757982896
transform 1 0 47600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2134
timestamp 1757982896
transform 1 0 49100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2135
timestamp 1757982896
transform 1 0 50600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2136
timestamp 1757982896
transform 1 0 52100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2137
timestamp 1757982896
transform 1 0 53600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2138
timestamp 1757982896
transform 1 0 55100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2139
timestamp 1757982896
transform 1 0 56600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2140
timestamp 1757982896
transform 1 0 58100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2141
timestamp 1757982896
transform 1 0 59600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2142
timestamp 1757982896
transform 1 0 61100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2143
timestamp 1757982896
transform 1 0 62600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2144
timestamp 1757982896
transform 1 0 64100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2145
timestamp 1757982896
transform 1 0 65600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2146
timestamp 1757982896
transform 1 0 67100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2147
timestamp 1757982896
transform 1 0 68600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2148
timestamp 1757982896
transform 1 0 70100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2149
timestamp 1757982896
transform 1 0 71600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2150
timestamp 1757982896
transform 1 0 73100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2151
timestamp 1757982896
transform 1 0 74600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2152
timestamp 1757982896
transform 1 0 76100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2153
timestamp 1757982896
transform 1 0 77600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2154
timestamp 1757982896
transform 1 0 79100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2155
timestamp 1757982896
transform 1 0 80600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2156
timestamp 1757982896
transform 1 0 82100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2157
timestamp 1757982896
transform 1 0 83600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2158
timestamp 1757982896
transform 1 0 85100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2159
timestamp 1757982896
transform 1 0 86600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2160
timestamp 1757982896
transform 1 0 88100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2161
timestamp 1757982896
transform 1 0 89600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2162
timestamp 1757982896
transform 1 0 91100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2163
timestamp 1757982896
transform 1 0 92600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2164
timestamp 1757982896
transform 1 0 94100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2165
timestamp 1757982896
transform 1 0 95600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2166
timestamp 1757982896
transform 1 0 97100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2167
timestamp 1757982896
transform 1 0 98600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2168
timestamp 1757982896
transform 1 0 100100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2169
timestamp 1757982896
transform 1 0 101600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2170
timestamp 1757982896
transform 1 0 103100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2171
timestamp 1757982896
transform 1 0 104600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2172
timestamp 1757982896
transform 1 0 106100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2173
timestamp 1757982896
transform 1 0 107600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2174
timestamp 1757982896
transform 1 0 109100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2175
timestamp 1757982896
transform 1 0 110600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2176
timestamp 1757982896
transform 1 0 112100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2177
timestamp 1757982896
transform 1 0 113600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2178
timestamp 1757982896
transform 1 0 115100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2179
timestamp 1757982896
transform 1 0 116600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2180
timestamp 1757982896
transform 1 0 118100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2181
timestamp 1757982896
transform 1 0 119600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2182
timestamp 1757982896
transform 1 0 121100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2183
timestamp 1757982896
transform 1 0 122600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2184
timestamp 1757982896
transform 1 0 124100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2185
timestamp 1757982896
transform 1 0 125600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2186
timestamp 1757982896
transform 1 0 127100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2187
timestamp 1757982896
transform 1 0 128600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2188
timestamp 1757982896
transform 1 0 130100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2189
timestamp 1757982896
transform 1 0 131600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2190
timestamp 1757982896
transform 1 0 133100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2191
timestamp 1757982896
transform 1 0 134600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2192
timestamp 1757982896
transform 1 0 136100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2193
timestamp 1757982896
transform 1 0 137600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2194
timestamp 1757982896
transform 1 0 139100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2195
timestamp 1757982896
transform 1 0 140600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2196
timestamp 1757982896
transform 1 0 142100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2197
timestamp 1757982896
transform 1 0 143600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2198
timestamp 1757982896
transform 1 0 145100 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2199
timestamp 1757982896
transform 1 0 146600 0 1 -30150
box 1820 -1430 3480 230
use pixel  pixel_2200
timestamp 1757982896
transform 1 0 -1900 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2201
timestamp 1757982896
transform 1 0 -400 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2202
timestamp 1757982896
transform 1 0 1100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2203
timestamp 1757982896
transform 1 0 2600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2204
timestamp 1757982896
transform 1 0 4100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2205
timestamp 1757982896
transform 1 0 5600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2206
timestamp 1757982896
transform 1 0 7100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2207
timestamp 1757982896
transform 1 0 8600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2208
timestamp 1757982896
transform 1 0 10100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2209
timestamp 1757982896
transform 1 0 11600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2210
timestamp 1757982896
transform 1 0 13100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2211
timestamp 1757982896
transform 1 0 14600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2212
timestamp 1757982896
transform 1 0 16100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2213
timestamp 1757982896
transform 1 0 17600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2214
timestamp 1757982896
transform 1 0 19100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2215
timestamp 1757982896
transform 1 0 20600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2216
timestamp 1757982896
transform 1 0 22100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2217
timestamp 1757982896
transform 1 0 23600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2218
timestamp 1757982896
transform 1 0 25100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2219
timestamp 1757982896
transform 1 0 26600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2220
timestamp 1757982896
transform 1 0 28100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2221
timestamp 1757982896
transform 1 0 29600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2222
timestamp 1757982896
transform 1 0 31100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2223
timestamp 1757982896
transform 1 0 32600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2224
timestamp 1757982896
transform 1 0 34100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2225
timestamp 1757982896
transform 1 0 35600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2226
timestamp 1757982896
transform 1 0 37100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2227
timestamp 1757982896
transform 1 0 38600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2228
timestamp 1757982896
transform 1 0 40100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2229
timestamp 1757982896
transform 1 0 41600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2230
timestamp 1757982896
transform 1 0 43100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2231
timestamp 1757982896
transform 1 0 44600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2232
timestamp 1757982896
transform 1 0 46100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2233
timestamp 1757982896
transform 1 0 47600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2234
timestamp 1757982896
transform 1 0 49100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2235
timestamp 1757982896
transform 1 0 50600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2236
timestamp 1757982896
transform 1 0 52100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2237
timestamp 1757982896
transform 1 0 53600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2238
timestamp 1757982896
transform 1 0 55100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2239
timestamp 1757982896
transform 1 0 56600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2240
timestamp 1757982896
transform 1 0 58100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2241
timestamp 1757982896
transform 1 0 59600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2242
timestamp 1757982896
transform 1 0 61100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2243
timestamp 1757982896
transform 1 0 62600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2244
timestamp 1757982896
transform 1 0 64100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2245
timestamp 1757982896
transform 1 0 65600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2246
timestamp 1757982896
transform 1 0 67100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2247
timestamp 1757982896
transform 1 0 68600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2248
timestamp 1757982896
transform 1 0 70100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2249
timestamp 1757982896
transform 1 0 71600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2250
timestamp 1757982896
transform 1 0 73100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2251
timestamp 1757982896
transform 1 0 74600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2252
timestamp 1757982896
transform 1 0 76100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2253
timestamp 1757982896
transform 1 0 77600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2254
timestamp 1757982896
transform 1 0 79100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2255
timestamp 1757982896
transform 1 0 80600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2256
timestamp 1757982896
transform 1 0 82100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2257
timestamp 1757982896
transform 1 0 83600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2258
timestamp 1757982896
transform 1 0 85100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2259
timestamp 1757982896
transform 1 0 86600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2260
timestamp 1757982896
transform 1 0 88100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2261
timestamp 1757982896
transform 1 0 89600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2262
timestamp 1757982896
transform 1 0 91100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2263
timestamp 1757982896
transform 1 0 92600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2264
timestamp 1757982896
transform 1 0 94100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2265
timestamp 1757982896
transform 1 0 95600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2266
timestamp 1757982896
transform 1 0 97100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2267
timestamp 1757982896
transform 1 0 98600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2268
timestamp 1757982896
transform 1 0 100100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2269
timestamp 1757982896
transform 1 0 101600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2270
timestamp 1757982896
transform 1 0 103100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2271
timestamp 1757982896
transform 1 0 104600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2272
timestamp 1757982896
transform 1 0 106100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2273
timestamp 1757982896
transform 1 0 107600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2274
timestamp 1757982896
transform 1 0 109100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2275
timestamp 1757982896
transform 1 0 110600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2276
timestamp 1757982896
transform 1 0 112100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2277
timestamp 1757982896
transform 1 0 113600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2278
timestamp 1757982896
transform 1 0 115100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2279
timestamp 1757982896
transform 1 0 116600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2280
timestamp 1757982896
transform 1 0 118100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2281
timestamp 1757982896
transform 1 0 119600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2282
timestamp 1757982896
transform 1 0 121100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2283
timestamp 1757982896
transform 1 0 122600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2284
timestamp 1757982896
transform 1 0 124100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2285
timestamp 1757982896
transform 1 0 125600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2286
timestamp 1757982896
transform 1 0 127100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2287
timestamp 1757982896
transform 1 0 128600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2288
timestamp 1757982896
transform 1 0 130100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2289
timestamp 1757982896
transform 1 0 131600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2290
timestamp 1757982896
transform 1 0 133100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2291
timestamp 1757982896
transform 1 0 134600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2292
timestamp 1757982896
transform 1 0 136100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2293
timestamp 1757982896
transform 1 0 137600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2294
timestamp 1757982896
transform 1 0 139100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2295
timestamp 1757982896
transform 1 0 140600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2296
timestamp 1757982896
transform 1 0 142100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2297
timestamp 1757982896
transform 1 0 143600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2298
timestamp 1757982896
transform 1 0 145100 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2299
timestamp 1757982896
transform 1 0 146600 0 1 -31650
box 1820 -1430 3480 230
use pixel  pixel_2300
timestamp 1757982896
transform 1 0 -1900 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2301
timestamp 1757982896
transform 1 0 -400 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2302
timestamp 1757982896
transform 1 0 1100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2303
timestamp 1757982896
transform 1 0 2600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2304
timestamp 1757982896
transform 1 0 4100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2305
timestamp 1757982896
transform 1 0 5600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2306
timestamp 1757982896
transform 1 0 7100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2307
timestamp 1757982896
transform 1 0 8600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2308
timestamp 1757982896
transform 1 0 10100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2309
timestamp 1757982896
transform 1 0 11600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2310
timestamp 1757982896
transform 1 0 13100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2311
timestamp 1757982896
transform 1 0 14600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2312
timestamp 1757982896
transform 1 0 16100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2313
timestamp 1757982896
transform 1 0 17600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2314
timestamp 1757982896
transform 1 0 19100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2315
timestamp 1757982896
transform 1 0 20600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2316
timestamp 1757982896
transform 1 0 22100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2317
timestamp 1757982896
transform 1 0 23600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2318
timestamp 1757982896
transform 1 0 25100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2319
timestamp 1757982896
transform 1 0 26600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2320
timestamp 1757982896
transform 1 0 28100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2321
timestamp 1757982896
transform 1 0 29600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2322
timestamp 1757982896
transform 1 0 31100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2323
timestamp 1757982896
transform 1 0 32600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2324
timestamp 1757982896
transform 1 0 34100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2325
timestamp 1757982896
transform 1 0 35600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2326
timestamp 1757982896
transform 1 0 37100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2327
timestamp 1757982896
transform 1 0 38600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2328
timestamp 1757982896
transform 1 0 40100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2329
timestamp 1757982896
transform 1 0 41600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2330
timestamp 1757982896
transform 1 0 43100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2331
timestamp 1757982896
transform 1 0 44600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2332
timestamp 1757982896
transform 1 0 46100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2333
timestamp 1757982896
transform 1 0 47600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2334
timestamp 1757982896
transform 1 0 49100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2335
timestamp 1757982896
transform 1 0 50600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2336
timestamp 1757982896
transform 1 0 52100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2337
timestamp 1757982896
transform 1 0 53600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2338
timestamp 1757982896
transform 1 0 55100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2339
timestamp 1757982896
transform 1 0 56600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2340
timestamp 1757982896
transform 1 0 58100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2341
timestamp 1757982896
transform 1 0 59600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2342
timestamp 1757982896
transform 1 0 61100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2343
timestamp 1757982896
transform 1 0 62600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2344
timestamp 1757982896
transform 1 0 64100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2345
timestamp 1757982896
transform 1 0 65600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2346
timestamp 1757982896
transform 1 0 67100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2347
timestamp 1757982896
transform 1 0 68600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2348
timestamp 1757982896
transform 1 0 70100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2349
timestamp 1757982896
transform 1 0 71600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2350
timestamp 1757982896
transform 1 0 73100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2351
timestamp 1757982896
transform 1 0 74600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2352
timestamp 1757982896
transform 1 0 76100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2353
timestamp 1757982896
transform 1 0 77600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2354
timestamp 1757982896
transform 1 0 79100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2355
timestamp 1757982896
transform 1 0 80600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2356
timestamp 1757982896
transform 1 0 82100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2357
timestamp 1757982896
transform 1 0 83600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2358
timestamp 1757982896
transform 1 0 85100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2359
timestamp 1757982896
transform 1 0 86600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2360
timestamp 1757982896
transform 1 0 88100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2361
timestamp 1757982896
transform 1 0 89600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2362
timestamp 1757982896
transform 1 0 91100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2363
timestamp 1757982896
transform 1 0 92600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2364
timestamp 1757982896
transform 1 0 94100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2365
timestamp 1757982896
transform 1 0 95600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2366
timestamp 1757982896
transform 1 0 97100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2367
timestamp 1757982896
transform 1 0 98600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2368
timestamp 1757982896
transform 1 0 100100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2369
timestamp 1757982896
transform 1 0 101600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2370
timestamp 1757982896
transform 1 0 103100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2371
timestamp 1757982896
transform 1 0 104600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2372
timestamp 1757982896
transform 1 0 106100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2373
timestamp 1757982896
transform 1 0 107600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2374
timestamp 1757982896
transform 1 0 109100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2375
timestamp 1757982896
transform 1 0 110600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2376
timestamp 1757982896
transform 1 0 112100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2377
timestamp 1757982896
transform 1 0 113600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2378
timestamp 1757982896
transform 1 0 115100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2379
timestamp 1757982896
transform 1 0 116600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2380
timestamp 1757982896
transform 1 0 118100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2381
timestamp 1757982896
transform 1 0 119600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2382
timestamp 1757982896
transform 1 0 121100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2383
timestamp 1757982896
transform 1 0 122600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2384
timestamp 1757982896
transform 1 0 124100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2385
timestamp 1757982896
transform 1 0 125600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2386
timestamp 1757982896
transform 1 0 127100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2387
timestamp 1757982896
transform 1 0 128600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2388
timestamp 1757982896
transform 1 0 130100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2389
timestamp 1757982896
transform 1 0 131600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2390
timestamp 1757982896
transform 1 0 133100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2391
timestamp 1757982896
transform 1 0 134600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2392
timestamp 1757982896
transform 1 0 136100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2393
timestamp 1757982896
transform 1 0 137600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2394
timestamp 1757982896
transform 1 0 139100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2395
timestamp 1757982896
transform 1 0 140600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2396
timestamp 1757982896
transform 1 0 142100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2397
timestamp 1757982896
transform 1 0 143600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2398
timestamp 1757982896
transform 1 0 145100 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2399
timestamp 1757982896
transform 1 0 146600 0 1 -33150
box 1820 -1430 3480 230
use pixel  pixel_2400
timestamp 1757982896
transform 1 0 -1900 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2401
timestamp 1757982896
transform 1 0 -400 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2402
timestamp 1757982896
transform 1 0 1100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2403
timestamp 1757982896
transform 1 0 2600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2404
timestamp 1757982896
transform 1 0 4100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2405
timestamp 1757982896
transform 1 0 5600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2406
timestamp 1757982896
transform 1 0 7100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2407
timestamp 1757982896
transform 1 0 8600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2408
timestamp 1757982896
transform 1 0 10100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2409
timestamp 1757982896
transform 1 0 11600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2410
timestamp 1757982896
transform 1 0 13100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2411
timestamp 1757982896
transform 1 0 14600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2412
timestamp 1757982896
transform 1 0 16100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2413
timestamp 1757982896
transform 1 0 17600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2414
timestamp 1757982896
transform 1 0 19100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2415
timestamp 1757982896
transform 1 0 20600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2416
timestamp 1757982896
transform 1 0 22100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2417
timestamp 1757982896
transform 1 0 23600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2418
timestamp 1757982896
transform 1 0 25100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2419
timestamp 1757982896
transform 1 0 26600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2420
timestamp 1757982896
transform 1 0 28100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2421
timestamp 1757982896
transform 1 0 29600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2422
timestamp 1757982896
transform 1 0 31100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2423
timestamp 1757982896
transform 1 0 32600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2424
timestamp 1757982896
transform 1 0 34100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2425
timestamp 1757982896
transform 1 0 35600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2426
timestamp 1757982896
transform 1 0 37100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2427
timestamp 1757982896
transform 1 0 38600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2428
timestamp 1757982896
transform 1 0 40100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2429
timestamp 1757982896
transform 1 0 41600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2430
timestamp 1757982896
transform 1 0 43100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2431
timestamp 1757982896
transform 1 0 44600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2432
timestamp 1757982896
transform 1 0 46100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2433
timestamp 1757982896
transform 1 0 47600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2434
timestamp 1757982896
transform 1 0 49100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2435
timestamp 1757982896
transform 1 0 50600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2436
timestamp 1757982896
transform 1 0 52100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2437
timestamp 1757982896
transform 1 0 53600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2438
timestamp 1757982896
transform 1 0 55100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2439
timestamp 1757982896
transform 1 0 56600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2440
timestamp 1757982896
transform 1 0 58100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2441
timestamp 1757982896
transform 1 0 59600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2442
timestamp 1757982896
transform 1 0 61100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2443
timestamp 1757982896
transform 1 0 62600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2444
timestamp 1757982896
transform 1 0 64100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2445
timestamp 1757982896
transform 1 0 65600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2446
timestamp 1757982896
transform 1 0 67100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2447
timestamp 1757982896
transform 1 0 68600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2448
timestamp 1757982896
transform 1 0 70100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2449
timestamp 1757982896
transform 1 0 71600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2450
timestamp 1757982896
transform 1 0 73100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2451
timestamp 1757982896
transform 1 0 74600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2452
timestamp 1757982896
transform 1 0 76100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2453
timestamp 1757982896
transform 1 0 77600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2454
timestamp 1757982896
transform 1 0 79100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2455
timestamp 1757982896
transform 1 0 80600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2456
timestamp 1757982896
transform 1 0 82100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2457
timestamp 1757982896
transform 1 0 83600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2458
timestamp 1757982896
transform 1 0 85100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2459
timestamp 1757982896
transform 1 0 86600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2460
timestamp 1757982896
transform 1 0 88100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2461
timestamp 1757982896
transform 1 0 89600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2462
timestamp 1757982896
transform 1 0 91100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2463
timestamp 1757982896
transform 1 0 92600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2464
timestamp 1757982896
transform 1 0 94100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2465
timestamp 1757982896
transform 1 0 95600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2466
timestamp 1757982896
transform 1 0 97100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2467
timestamp 1757982896
transform 1 0 98600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2468
timestamp 1757982896
transform 1 0 100100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2469
timestamp 1757982896
transform 1 0 101600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2470
timestamp 1757982896
transform 1 0 103100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2471
timestamp 1757982896
transform 1 0 104600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2472
timestamp 1757982896
transform 1 0 106100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2473
timestamp 1757982896
transform 1 0 107600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2474
timestamp 1757982896
transform 1 0 109100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2475
timestamp 1757982896
transform 1 0 110600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2476
timestamp 1757982896
transform 1 0 112100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2477
timestamp 1757982896
transform 1 0 113600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2478
timestamp 1757982896
transform 1 0 115100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2479
timestamp 1757982896
transform 1 0 116600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2480
timestamp 1757982896
transform 1 0 118100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2481
timestamp 1757982896
transform 1 0 119600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2482
timestamp 1757982896
transform 1 0 121100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2483
timestamp 1757982896
transform 1 0 122600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2484
timestamp 1757982896
transform 1 0 124100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2485
timestamp 1757982896
transform 1 0 125600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2486
timestamp 1757982896
transform 1 0 127100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2487
timestamp 1757982896
transform 1 0 128600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2488
timestamp 1757982896
transform 1 0 130100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2489
timestamp 1757982896
transform 1 0 131600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2490
timestamp 1757982896
transform 1 0 133100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2491
timestamp 1757982896
transform 1 0 134600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2492
timestamp 1757982896
transform 1 0 136100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2493
timestamp 1757982896
transform 1 0 137600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2494
timestamp 1757982896
transform 1 0 139100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2495
timestamp 1757982896
transform 1 0 140600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2496
timestamp 1757982896
transform 1 0 142100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2497
timestamp 1757982896
transform 1 0 143600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2498
timestamp 1757982896
transform 1 0 145100 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2499
timestamp 1757982896
transform 1 0 146600 0 1 -34650
box 1820 -1430 3480 230
use pixel  pixel_2500
timestamp 1757982896
transform 1 0 -1900 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2501
timestamp 1757982896
transform 1 0 -400 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2502
timestamp 1757982896
transform 1 0 1100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2503
timestamp 1757982896
transform 1 0 2600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2504
timestamp 1757982896
transform 1 0 4100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2505
timestamp 1757982896
transform 1 0 5600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2506
timestamp 1757982896
transform 1 0 7100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2507
timestamp 1757982896
transform 1 0 8600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2508
timestamp 1757982896
transform 1 0 10100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2509
timestamp 1757982896
transform 1 0 11600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2510
timestamp 1757982896
transform 1 0 13100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2511
timestamp 1757982896
transform 1 0 14600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2512
timestamp 1757982896
transform 1 0 16100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2513
timestamp 1757982896
transform 1 0 17600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2514
timestamp 1757982896
transform 1 0 19100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2515
timestamp 1757982896
transform 1 0 20600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2516
timestamp 1757982896
transform 1 0 22100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2517
timestamp 1757982896
transform 1 0 23600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2518
timestamp 1757982896
transform 1 0 25100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2519
timestamp 1757982896
transform 1 0 26600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2520
timestamp 1757982896
transform 1 0 28100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2521
timestamp 1757982896
transform 1 0 29600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2522
timestamp 1757982896
transform 1 0 31100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2523
timestamp 1757982896
transform 1 0 32600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2524
timestamp 1757982896
transform 1 0 34100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2525
timestamp 1757982896
transform 1 0 35600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2526
timestamp 1757982896
transform 1 0 37100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2527
timestamp 1757982896
transform 1 0 38600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2528
timestamp 1757982896
transform 1 0 40100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2529
timestamp 1757982896
transform 1 0 41600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2530
timestamp 1757982896
transform 1 0 43100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2531
timestamp 1757982896
transform 1 0 44600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2532
timestamp 1757982896
transform 1 0 46100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2533
timestamp 1757982896
transform 1 0 47600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2534
timestamp 1757982896
transform 1 0 49100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2535
timestamp 1757982896
transform 1 0 50600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2536
timestamp 1757982896
transform 1 0 52100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2537
timestamp 1757982896
transform 1 0 53600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2538
timestamp 1757982896
transform 1 0 55100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2539
timestamp 1757982896
transform 1 0 56600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2540
timestamp 1757982896
transform 1 0 58100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2541
timestamp 1757982896
transform 1 0 59600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2542
timestamp 1757982896
transform 1 0 61100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2543
timestamp 1757982896
transform 1 0 62600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2544
timestamp 1757982896
transform 1 0 64100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2545
timestamp 1757982896
transform 1 0 65600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2546
timestamp 1757982896
transform 1 0 67100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2547
timestamp 1757982896
transform 1 0 68600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2548
timestamp 1757982896
transform 1 0 70100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2549
timestamp 1757982896
transform 1 0 71600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2550
timestamp 1757982896
transform 1 0 73100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2551
timestamp 1757982896
transform 1 0 74600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2552
timestamp 1757982896
transform 1 0 76100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2553
timestamp 1757982896
transform 1 0 77600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2554
timestamp 1757982896
transform 1 0 79100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2555
timestamp 1757982896
transform 1 0 80600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2556
timestamp 1757982896
transform 1 0 82100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2557
timestamp 1757982896
transform 1 0 83600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2558
timestamp 1757982896
transform 1 0 85100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2559
timestamp 1757982896
transform 1 0 86600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2560
timestamp 1757982896
transform 1 0 88100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2561
timestamp 1757982896
transform 1 0 89600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2562
timestamp 1757982896
transform 1 0 91100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2563
timestamp 1757982896
transform 1 0 92600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2564
timestamp 1757982896
transform 1 0 94100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2565
timestamp 1757982896
transform 1 0 95600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2566
timestamp 1757982896
transform 1 0 97100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2567
timestamp 1757982896
transform 1 0 98600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2568
timestamp 1757982896
transform 1 0 100100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2569
timestamp 1757982896
transform 1 0 101600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2570
timestamp 1757982896
transform 1 0 103100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2571
timestamp 1757982896
transform 1 0 104600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2572
timestamp 1757982896
transform 1 0 106100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2573
timestamp 1757982896
transform 1 0 107600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2574
timestamp 1757982896
transform 1 0 109100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2575
timestamp 1757982896
transform 1 0 110600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2576
timestamp 1757982896
transform 1 0 112100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2577
timestamp 1757982896
transform 1 0 113600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2578
timestamp 1757982896
transform 1 0 115100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2579
timestamp 1757982896
transform 1 0 116600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2580
timestamp 1757982896
transform 1 0 118100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2581
timestamp 1757982896
transform 1 0 119600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2582
timestamp 1757982896
transform 1 0 121100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2583
timestamp 1757982896
transform 1 0 122600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2584
timestamp 1757982896
transform 1 0 124100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2585
timestamp 1757982896
transform 1 0 125600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2586
timestamp 1757982896
transform 1 0 127100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2587
timestamp 1757982896
transform 1 0 128600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2588
timestamp 1757982896
transform 1 0 130100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2589
timestamp 1757982896
transform 1 0 131600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2590
timestamp 1757982896
transform 1 0 133100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2591
timestamp 1757982896
transform 1 0 134600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2592
timestamp 1757982896
transform 1 0 136100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2593
timestamp 1757982896
transform 1 0 137600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2594
timestamp 1757982896
transform 1 0 139100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2595
timestamp 1757982896
transform 1 0 140600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2596
timestamp 1757982896
transform 1 0 142100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2597
timestamp 1757982896
transform 1 0 143600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2598
timestamp 1757982896
transform 1 0 145100 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2599
timestamp 1757982896
transform 1 0 146600 0 1 -36150
box 1820 -1430 3480 230
use pixel  pixel_2600
timestamp 1757982896
transform 1 0 -1900 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2601
timestamp 1757982896
transform 1 0 -400 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2602
timestamp 1757982896
transform 1 0 1100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2603
timestamp 1757982896
transform 1 0 2600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2604
timestamp 1757982896
transform 1 0 4100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2605
timestamp 1757982896
transform 1 0 5600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2606
timestamp 1757982896
transform 1 0 7100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2607
timestamp 1757982896
transform 1 0 8600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2608
timestamp 1757982896
transform 1 0 10100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2609
timestamp 1757982896
transform 1 0 11600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2610
timestamp 1757982896
transform 1 0 13100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2611
timestamp 1757982896
transform 1 0 14600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2612
timestamp 1757982896
transform 1 0 16100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2613
timestamp 1757982896
transform 1 0 17600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2614
timestamp 1757982896
transform 1 0 19100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2615
timestamp 1757982896
transform 1 0 20600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2616
timestamp 1757982896
transform 1 0 22100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2617
timestamp 1757982896
transform 1 0 23600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2618
timestamp 1757982896
transform 1 0 25100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2619
timestamp 1757982896
transform 1 0 26600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2620
timestamp 1757982896
transform 1 0 28100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2621
timestamp 1757982896
transform 1 0 29600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2622
timestamp 1757982896
transform 1 0 31100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2623
timestamp 1757982896
transform 1 0 32600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2624
timestamp 1757982896
transform 1 0 34100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2625
timestamp 1757982896
transform 1 0 35600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2626
timestamp 1757982896
transform 1 0 37100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2627
timestamp 1757982896
transform 1 0 38600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2628
timestamp 1757982896
transform 1 0 40100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2629
timestamp 1757982896
transform 1 0 41600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2630
timestamp 1757982896
transform 1 0 43100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2631
timestamp 1757982896
transform 1 0 44600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2632
timestamp 1757982896
transform 1 0 46100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2633
timestamp 1757982896
transform 1 0 47600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2634
timestamp 1757982896
transform 1 0 49100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2635
timestamp 1757982896
transform 1 0 50600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2636
timestamp 1757982896
transform 1 0 52100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2637
timestamp 1757982896
transform 1 0 53600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2638
timestamp 1757982896
transform 1 0 55100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2639
timestamp 1757982896
transform 1 0 56600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2640
timestamp 1757982896
transform 1 0 58100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2641
timestamp 1757982896
transform 1 0 59600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2642
timestamp 1757982896
transform 1 0 61100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2643
timestamp 1757982896
transform 1 0 62600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2644
timestamp 1757982896
transform 1 0 64100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2645
timestamp 1757982896
transform 1 0 65600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2646
timestamp 1757982896
transform 1 0 67100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2647
timestamp 1757982896
transform 1 0 68600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2648
timestamp 1757982896
transform 1 0 70100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2649
timestamp 1757982896
transform 1 0 71600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2650
timestamp 1757982896
transform 1 0 73100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2651
timestamp 1757982896
transform 1 0 74600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2652
timestamp 1757982896
transform 1 0 76100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2653
timestamp 1757982896
transform 1 0 77600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2654
timestamp 1757982896
transform 1 0 79100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2655
timestamp 1757982896
transform 1 0 80600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2656
timestamp 1757982896
transform 1 0 82100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2657
timestamp 1757982896
transform 1 0 83600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2658
timestamp 1757982896
transform 1 0 85100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2659
timestamp 1757982896
transform 1 0 86600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2660
timestamp 1757982896
transform 1 0 88100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2661
timestamp 1757982896
transform 1 0 89600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2662
timestamp 1757982896
transform 1 0 91100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2663
timestamp 1757982896
transform 1 0 92600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2664
timestamp 1757982896
transform 1 0 94100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2665
timestamp 1757982896
transform 1 0 95600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2666
timestamp 1757982896
transform 1 0 97100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2667
timestamp 1757982896
transform 1 0 98600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2668
timestamp 1757982896
transform 1 0 100100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2669
timestamp 1757982896
transform 1 0 101600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2670
timestamp 1757982896
transform 1 0 103100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2671
timestamp 1757982896
transform 1 0 104600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2672
timestamp 1757982896
transform 1 0 106100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2673
timestamp 1757982896
transform 1 0 107600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2674
timestamp 1757982896
transform 1 0 109100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2675
timestamp 1757982896
transform 1 0 110600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2676
timestamp 1757982896
transform 1 0 112100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2677
timestamp 1757982896
transform 1 0 113600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2678
timestamp 1757982896
transform 1 0 115100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2679
timestamp 1757982896
transform 1 0 116600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2680
timestamp 1757982896
transform 1 0 118100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2681
timestamp 1757982896
transform 1 0 119600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2682
timestamp 1757982896
transform 1 0 121100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2683
timestamp 1757982896
transform 1 0 122600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2684
timestamp 1757982896
transform 1 0 124100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2685
timestamp 1757982896
transform 1 0 125600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2686
timestamp 1757982896
transform 1 0 127100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2687
timestamp 1757982896
transform 1 0 128600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2688
timestamp 1757982896
transform 1 0 130100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2689
timestamp 1757982896
transform 1 0 131600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2690
timestamp 1757982896
transform 1 0 133100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2691
timestamp 1757982896
transform 1 0 134600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2692
timestamp 1757982896
transform 1 0 136100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2693
timestamp 1757982896
transform 1 0 137600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2694
timestamp 1757982896
transform 1 0 139100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2695
timestamp 1757982896
transform 1 0 140600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2696
timestamp 1757982896
transform 1 0 142100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2697
timestamp 1757982896
transform 1 0 143600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2698
timestamp 1757982896
transform 1 0 145100 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2699
timestamp 1757982896
transform 1 0 146600 0 1 -37650
box 1820 -1430 3480 230
use pixel  pixel_2700
timestamp 1757982896
transform 1 0 -1900 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2701
timestamp 1757982896
transform 1 0 -400 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2702
timestamp 1757982896
transform 1 0 1100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2703
timestamp 1757982896
transform 1 0 2600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2704
timestamp 1757982896
transform 1 0 4100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2705
timestamp 1757982896
transform 1 0 5600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2706
timestamp 1757982896
transform 1 0 7100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2707
timestamp 1757982896
transform 1 0 8600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2708
timestamp 1757982896
transform 1 0 10100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2709
timestamp 1757982896
transform 1 0 11600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2710
timestamp 1757982896
transform 1 0 13100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2711
timestamp 1757982896
transform 1 0 14600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2712
timestamp 1757982896
transform 1 0 16100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2713
timestamp 1757982896
transform 1 0 17600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2714
timestamp 1757982896
transform 1 0 19100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2715
timestamp 1757982896
transform 1 0 20600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2716
timestamp 1757982896
transform 1 0 22100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2717
timestamp 1757982896
transform 1 0 23600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2718
timestamp 1757982896
transform 1 0 25100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2719
timestamp 1757982896
transform 1 0 26600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2720
timestamp 1757982896
transform 1 0 28100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2721
timestamp 1757982896
transform 1 0 29600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2722
timestamp 1757982896
transform 1 0 31100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2723
timestamp 1757982896
transform 1 0 32600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2724
timestamp 1757982896
transform 1 0 34100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2725
timestamp 1757982896
transform 1 0 35600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2726
timestamp 1757982896
transform 1 0 37100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2727
timestamp 1757982896
transform 1 0 38600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2728
timestamp 1757982896
transform 1 0 40100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2729
timestamp 1757982896
transform 1 0 41600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2730
timestamp 1757982896
transform 1 0 43100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2731
timestamp 1757982896
transform 1 0 44600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2732
timestamp 1757982896
transform 1 0 46100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2733
timestamp 1757982896
transform 1 0 47600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2734
timestamp 1757982896
transform 1 0 49100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2735
timestamp 1757982896
transform 1 0 50600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2736
timestamp 1757982896
transform 1 0 52100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2737
timestamp 1757982896
transform 1 0 53600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2738
timestamp 1757982896
transform 1 0 55100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2739
timestamp 1757982896
transform 1 0 56600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2740
timestamp 1757982896
transform 1 0 58100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2741
timestamp 1757982896
transform 1 0 59600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2742
timestamp 1757982896
transform 1 0 61100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2743
timestamp 1757982896
transform 1 0 62600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2744
timestamp 1757982896
transform 1 0 64100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2745
timestamp 1757982896
transform 1 0 65600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2746
timestamp 1757982896
transform 1 0 67100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2747
timestamp 1757982896
transform 1 0 68600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2748
timestamp 1757982896
transform 1 0 70100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2749
timestamp 1757982896
transform 1 0 71600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2750
timestamp 1757982896
transform 1 0 73100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2751
timestamp 1757982896
transform 1 0 74600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2752
timestamp 1757982896
transform 1 0 76100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2753
timestamp 1757982896
transform 1 0 77600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2754
timestamp 1757982896
transform 1 0 79100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2755
timestamp 1757982896
transform 1 0 80600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2756
timestamp 1757982896
transform 1 0 82100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2757
timestamp 1757982896
transform 1 0 83600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2758
timestamp 1757982896
transform 1 0 85100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2759
timestamp 1757982896
transform 1 0 86600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2760
timestamp 1757982896
transform 1 0 88100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2761
timestamp 1757982896
transform 1 0 89600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2762
timestamp 1757982896
transform 1 0 91100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2763
timestamp 1757982896
transform 1 0 92600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2764
timestamp 1757982896
transform 1 0 94100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2765
timestamp 1757982896
transform 1 0 95600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2766
timestamp 1757982896
transform 1 0 97100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2767
timestamp 1757982896
transform 1 0 98600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2768
timestamp 1757982896
transform 1 0 100100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2769
timestamp 1757982896
transform 1 0 101600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2770
timestamp 1757982896
transform 1 0 103100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2771
timestamp 1757982896
transform 1 0 104600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2772
timestamp 1757982896
transform 1 0 106100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2773
timestamp 1757982896
transform 1 0 107600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2774
timestamp 1757982896
transform 1 0 109100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2775
timestamp 1757982896
transform 1 0 110600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2776
timestamp 1757982896
transform 1 0 112100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2777
timestamp 1757982896
transform 1 0 113600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2778
timestamp 1757982896
transform 1 0 115100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2779
timestamp 1757982896
transform 1 0 116600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2780
timestamp 1757982896
transform 1 0 118100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2781
timestamp 1757982896
transform 1 0 119600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2782
timestamp 1757982896
transform 1 0 121100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2783
timestamp 1757982896
transform 1 0 122600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2784
timestamp 1757982896
transform 1 0 124100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2785
timestamp 1757982896
transform 1 0 125600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2786
timestamp 1757982896
transform 1 0 127100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2787
timestamp 1757982896
transform 1 0 128600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2788
timestamp 1757982896
transform 1 0 130100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2789
timestamp 1757982896
transform 1 0 131600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2790
timestamp 1757982896
transform 1 0 133100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2791
timestamp 1757982896
transform 1 0 134600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2792
timestamp 1757982896
transform 1 0 136100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2793
timestamp 1757982896
transform 1 0 137600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2794
timestamp 1757982896
transform 1 0 139100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2795
timestamp 1757982896
transform 1 0 140600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2796
timestamp 1757982896
transform 1 0 142100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2797
timestamp 1757982896
transform 1 0 143600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2798
timestamp 1757982896
transform 1 0 145100 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2799
timestamp 1757982896
transform 1 0 146600 0 1 -39150
box 1820 -1430 3480 230
use pixel  pixel_2800
timestamp 1757982896
transform 1 0 -1900 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2801
timestamp 1757982896
transform 1 0 -400 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2802
timestamp 1757982896
transform 1 0 1100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2803
timestamp 1757982896
transform 1 0 2600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2804
timestamp 1757982896
transform 1 0 4100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2805
timestamp 1757982896
transform 1 0 5600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2806
timestamp 1757982896
transform 1 0 7100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2807
timestamp 1757982896
transform 1 0 8600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2808
timestamp 1757982896
transform 1 0 10100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2809
timestamp 1757982896
transform 1 0 11600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2810
timestamp 1757982896
transform 1 0 13100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2811
timestamp 1757982896
transform 1 0 14600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2812
timestamp 1757982896
transform 1 0 16100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2813
timestamp 1757982896
transform 1 0 17600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2814
timestamp 1757982896
transform 1 0 19100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2815
timestamp 1757982896
transform 1 0 20600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2816
timestamp 1757982896
transform 1 0 22100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2817
timestamp 1757982896
transform 1 0 23600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2818
timestamp 1757982896
transform 1 0 25100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2819
timestamp 1757982896
transform 1 0 26600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2820
timestamp 1757982896
transform 1 0 28100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2821
timestamp 1757982896
transform 1 0 29600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2822
timestamp 1757982896
transform 1 0 31100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2823
timestamp 1757982896
transform 1 0 32600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2824
timestamp 1757982896
transform 1 0 34100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2825
timestamp 1757982896
transform 1 0 35600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2826
timestamp 1757982896
transform 1 0 37100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2827
timestamp 1757982896
transform 1 0 38600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2828
timestamp 1757982896
transform 1 0 40100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2829
timestamp 1757982896
transform 1 0 41600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2830
timestamp 1757982896
transform 1 0 43100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2831
timestamp 1757982896
transform 1 0 44600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2832
timestamp 1757982896
transform 1 0 46100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2833
timestamp 1757982896
transform 1 0 47600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2834
timestamp 1757982896
transform 1 0 49100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2835
timestamp 1757982896
transform 1 0 50600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2836
timestamp 1757982896
transform 1 0 52100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2837
timestamp 1757982896
transform 1 0 53600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2838
timestamp 1757982896
transform 1 0 55100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2839
timestamp 1757982896
transform 1 0 56600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2840
timestamp 1757982896
transform 1 0 58100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2841
timestamp 1757982896
transform 1 0 59600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2842
timestamp 1757982896
transform 1 0 61100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2843
timestamp 1757982896
transform 1 0 62600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2844
timestamp 1757982896
transform 1 0 64100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2845
timestamp 1757982896
transform 1 0 65600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2846
timestamp 1757982896
transform 1 0 67100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2847
timestamp 1757982896
transform 1 0 68600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2848
timestamp 1757982896
transform 1 0 70100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2849
timestamp 1757982896
transform 1 0 71600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2850
timestamp 1757982896
transform 1 0 73100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2851
timestamp 1757982896
transform 1 0 74600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2852
timestamp 1757982896
transform 1 0 76100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2853
timestamp 1757982896
transform 1 0 77600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2854
timestamp 1757982896
transform 1 0 79100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2855
timestamp 1757982896
transform 1 0 80600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2856
timestamp 1757982896
transform 1 0 82100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2857
timestamp 1757982896
transform 1 0 83600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2858
timestamp 1757982896
transform 1 0 85100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2859
timestamp 1757982896
transform 1 0 86600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2860
timestamp 1757982896
transform 1 0 88100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2861
timestamp 1757982896
transform 1 0 89600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2862
timestamp 1757982896
transform 1 0 91100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2863
timestamp 1757982896
transform 1 0 92600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2864
timestamp 1757982896
transform 1 0 94100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2865
timestamp 1757982896
transform 1 0 95600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2866
timestamp 1757982896
transform 1 0 97100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2867
timestamp 1757982896
transform 1 0 98600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2868
timestamp 1757982896
transform 1 0 100100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2869
timestamp 1757982896
transform 1 0 101600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2870
timestamp 1757982896
transform 1 0 103100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2871
timestamp 1757982896
transform 1 0 104600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2872
timestamp 1757982896
transform 1 0 106100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2873
timestamp 1757982896
transform 1 0 107600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2874
timestamp 1757982896
transform 1 0 109100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2875
timestamp 1757982896
transform 1 0 110600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2876
timestamp 1757982896
transform 1 0 112100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2877
timestamp 1757982896
transform 1 0 113600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2878
timestamp 1757982896
transform 1 0 115100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2879
timestamp 1757982896
transform 1 0 116600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2880
timestamp 1757982896
transform 1 0 118100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2881
timestamp 1757982896
transform 1 0 119600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2882
timestamp 1757982896
transform 1 0 121100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2883
timestamp 1757982896
transform 1 0 122600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2884
timestamp 1757982896
transform 1 0 124100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2885
timestamp 1757982896
transform 1 0 125600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2886
timestamp 1757982896
transform 1 0 127100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2887
timestamp 1757982896
transform 1 0 128600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2888
timestamp 1757982896
transform 1 0 130100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2889
timestamp 1757982896
transform 1 0 131600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2890
timestamp 1757982896
transform 1 0 133100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2891
timestamp 1757982896
transform 1 0 134600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2892
timestamp 1757982896
transform 1 0 136100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2893
timestamp 1757982896
transform 1 0 137600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2894
timestamp 1757982896
transform 1 0 139100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2895
timestamp 1757982896
transform 1 0 140600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2896
timestamp 1757982896
transform 1 0 142100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2897
timestamp 1757982896
transform 1 0 143600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2898
timestamp 1757982896
transform 1 0 145100 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2899
timestamp 1757982896
transform 1 0 146600 0 1 -40650
box 1820 -1430 3480 230
use pixel  pixel_2900
timestamp 1757982896
transform 1 0 -1900 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2901
timestamp 1757982896
transform 1 0 -400 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2902
timestamp 1757982896
transform 1 0 1100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2903
timestamp 1757982896
transform 1 0 2600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2904
timestamp 1757982896
transform 1 0 4100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2905
timestamp 1757982896
transform 1 0 5600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2906
timestamp 1757982896
transform 1 0 7100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2907
timestamp 1757982896
transform 1 0 8600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2908
timestamp 1757982896
transform 1 0 10100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2909
timestamp 1757982896
transform 1 0 11600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2910
timestamp 1757982896
transform 1 0 13100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2911
timestamp 1757982896
transform 1 0 14600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2912
timestamp 1757982896
transform 1 0 16100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2913
timestamp 1757982896
transform 1 0 17600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2914
timestamp 1757982896
transform 1 0 19100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2915
timestamp 1757982896
transform 1 0 20600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2916
timestamp 1757982896
transform 1 0 22100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2917
timestamp 1757982896
transform 1 0 23600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2918
timestamp 1757982896
transform 1 0 25100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2919
timestamp 1757982896
transform 1 0 26600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2920
timestamp 1757982896
transform 1 0 28100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2921
timestamp 1757982896
transform 1 0 29600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2922
timestamp 1757982896
transform 1 0 31100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2923
timestamp 1757982896
transform 1 0 32600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2924
timestamp 1757982896
transform 1 0 34100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2925
timestamp 1757982896
transform 1 0 35600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2926
timestamp 1757982896
transform 1 0 37100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2927
timestamp 1757982896
transform 1 0 38600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2928
timestamp 1757982896
transform 1 0 40100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2929
timestamp 1757982896
transform 1 0 41600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2930
timestamp 1757982896
transform 1 0 43100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2931
timestamp 1757982896
transform 1 0 44600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2932
timestamp 1757982896
transform 1 0 46100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2933
timestamp 1757982896
transform 1 0 47600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2934
timestamp 1757982896
transform 1 0 49100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2935
timestamp 1757982896
transform 1 0 50600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2936
timestamp 1757982896
transform 1 0 52100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2937
timestamp 1757982896
transform 1 0 53600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2938
timestamp 1757982896
transform 1 0 55100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2939
timestamp 1757982896
transform 1 0 56600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2940
timestamp 1757982896
transform 1 0 58100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2941
timestamp 1757982896
transform 1 0 59600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2942
timestamp 1757982896
transform 1 0 61100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2943
timestamp 1757982896
transform 1 0 62600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2944
timestamp 1757982896
transform 1 0 64100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2945
timestamp 1757982896
transform 1 0 65600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2946
timestamp 1757982896
transform 1 0 67100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2947
timestamp 1757982896
transform 1 0 68600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2948
timestamp 1757982896
transform 1 0 70100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2949
timestamp 1757982896
transform 1 0 71600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2950
timestamp 1757982896
transform 1 0 73100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2951
timestamp 1757982896
transform 1 0 74600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2952
timestamp 1757982896
transform 1 0 76100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2953
timestamp 1757982896
transform 1 0 77600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2954
timestamp 1757982896
transform 1 0 79100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2955
timestamp 1757982896
transform 1 0 80600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2956
timestamp 1757982896
transform 1 0 82100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2957
timestamp 1757982896
transform 1 0 83600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2958
timestamp 1757982896
transform 1 0 85100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2959
timestamp 1757982896
transform 1 0 86600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2960
timestamp 1757982896
transform 1 0 88100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2961
timestamp 1757982896
transform 1 0 89600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2962
timestamp 1757982896
transform 1 0 91100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2963
timestamp 1757982896
transform 1 0 92600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2964
timestamp 1757982896
transform 1 0 94100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2965
timestamp 1757982896
transform 1 0 95600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2966
timestamp 1757982896
transform 1 0 97100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2967
timestamp 1757982896
transform 1 0 98600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2968
timestamp 1757982896
transform 1 0 100100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2969
timestamp 1757982896
transform 1 0 101600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2970
timestamp 1757982896
transform 1 0 103100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2971
timestamp 1757982896
transform 1 0 104600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2972
timestamp 1757982896
transform 1 0 106100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2973
timestamp 1757982896
transform 1 0 107600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2974
timestamp 1757982896
transform 1 0 109100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2975
timestamp 1757982896
transform 1 0 110600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2976
timestamp 1757982896
transform 1 0 112100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2977
timestamp 1757982896
transform 1 0 113600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2978
timestamp 1757982896
transform 1 0 115100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2979
timestamp 1757982896
transform 1 0 116600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2980
timestamp 1757982896
transform 1 0 118100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2981
timestamp 1757982896
transform 1 0 119600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2982
timestamp 1757982896
transform 1 0 121100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2983
timestamp 1757982896
transform 1 0 122600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2984
timestamp 1757982896
transform 1 0 124100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2985
timestamp 1757982896
transform 1 0 125600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2986
timestamp 1757982896
transform 1 0 127100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2987
timestamp 1757982896
transform 1 0 128600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2988
timestamp 1757982896
transform 1 0 130100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2989
timestamp 1757982896
transform 1 0 131600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2990
timestamp 1757982896
transform 1 0 133100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2991
timestamp 1757982896
transform 1 0 134600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2992
timestamp 1757982896
transform 1 0 136100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2993
timestamp 1757982896
transform 1 0 137600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2994
timestamp 1757982896
transform 1 0 139100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2995
timestamp 1757982896
transform 1 0 140600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2996
timestamp 1757982896
transform 1 0 142100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2997
timestamp 1757982896
transform 1 0 143600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2998
timestamp 1757982896
transform 1 0 145100 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_2999
timestamp 1757982896
transform 1 0 146600 0 1 -42150
box 1820 -1430 3480 230
use pixel  pixel_3000
timestamp 1757982896
transform 1 0 -1900 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3001
timestamp 1757982896
transform 1 0 -400 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3002
timestamp 1757982896
transform 1 0 1100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3003
timestamp 1757982896
transform 1 0 2600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3004
timestamp 1757982896
transform 1 0 4100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3005
timestamp 1757982896
transform 1 0 5600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3006
timestamp 1757982896
transform 1 0 7100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3007
timestamp 1757982896
transform 1 0 8600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3008
timestamp 1757982896
transform 1 0 10100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3009
timestamp 1757982896
transform 1 0 11600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3010
timestamp 1757982896
transform 1 0 13100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3011
timestamp 1757982896
transform 1 0 14600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3012
timestamp 1757982896
transform 1 0 16100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3013
timestamp 1757982896
transform 1 0 17600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3014
timestamp 1757982896
transform 1 0 19100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3015
timestamp 1757982896
transform 1 0 20600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3016
timestamp 1757982896
transform 1 0 22100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3017
timestamp 1757982896
transform 1 0 23600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3018
timestamp 1757982896
transform 1 0 25100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3019
timestamp 1757982896
transform 1 0 26600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3020
timestamp 1757982896
transform 1 0 28100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3021
timestamp 1757982896
transform 1 0 29600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3022
timestamp 1757982896
transform 1 0 31100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3023
timestamp 1757982896
transform 1 0 32600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3024
timestamp 1757982896
transform 1 0 34100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3025
timestamp 1757982896
transform 1 0 35600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3026
timestamp 1757982896
transform 1 0 37100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3027
timestamp 1757982896
transform 1 0 38600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3028
timestamp 1757982896
transform 1 0 40100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3029
timestamp 1757982896
transform 1 0 41600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3030
timestamp 1757982896
transform 1 0 43100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3031
timestamp 1757982896
transform 1 0 44600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3032
timestamp 1757982896
transform 1 0 46100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3033
timestamp 1757982896
transform 1 0 47600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3034
timestamp 1757982896
transform 1 0 49100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3035
timestamp 1757982896
transform 1 0 50600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3036
timestamp 1757982896
transform 1 0 52100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3037
timestamp 1757982896
transform 1 0 53600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3038
timestamp 1757982896
transform 1 0 55100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3039
timestamp 1757982896
transform 1 0 56600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3040
timestamp 1757982896
transform 1 0 58100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3041
timestamp 1757982896
transform 1 0 59600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3042
timestamp 1757982896
transform 1 0 61100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3043
timestamp 1757982896
transform 1 0 62600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3044
timestamp 1757982896
transform 1 0 64100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3045
timestamp 1757982896
transform 1 0 65600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3046
timestamp 1757982896
transform 1 0 67100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3047
timestamp 1757982896
transform 1 0 68600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3048
timestamp 1757982896
transform 1 0 70100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3049
timestamp 1757982896
transform 1 0 71600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3050
timestamp 1757982896
transform 1 0 73100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3051
timestamp 1757982896
transform 1 0 74600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3052
timestamp 1757982896
transform 1 0 76100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3053
timestamp 1757982896
transform 1 0 77600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3054
timestamp 1757982896
transform 1 0 79100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3055
timestamp 1757982896
transform 1 0 80600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3056
timestamp 1757982896
transform 1 0 82100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3057
timestamp 1757982896
transform 1 0 83600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3058
timestamp 1757982896
transform 1 0 85100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3059
timestamp 1757982896
transform 1 0 86600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3060
timestamp 1757982896
transform 1 0 88100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3061
timestamp 1757982896
transform 1 0 89600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3062
timestamp 1757982896
transform 1 0 91100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3063
timestamp 1757982896
transform 1 0 92600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3064
timestamp 1757982896
transform 1 0 94100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3065
timestamp 1757982896
transform 1 0 95600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3066
timestamp 1757982896
transform 1 0 97100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3067
timestamp 1757982896
transform 1 0 98600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3068
timestamp 1757982896
transform 1 0 100100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3069
timestamp 1757982896
transform 1 0 101600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3070
timestamp 1757982896
transform 1 0 103100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3071
timestamp 1757982896
transform 1 0 104600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3072
timestamp 1757982896
transform 1 0 106100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3073
timestamp 1757982896
transform 1 0 107600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3074
timestamp 1757982896
transform 1 0 109100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3075
timestamp 1757982896
transform 1 0 110600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3076
timestamp 1757982896
transform 1 0 112100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3077
timestamp 1757982896
transform 1 0 113600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3078
timestamp 1757982896
transform 1 0 115100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3079
timestamp 1757982896
transform 1 0 116600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3080
timestamp 1757982896
transform 1 0 118100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3081
timestamp 1757982896
transform 1 0 119600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3082
timestamp 1757982896
transform 1 0 121100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3083
timestamp 1757982896
transform 1 0 122600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3084
timestamp 1757982896
transform 1 0 124100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3085
timestamp 1757982896
transform 1 0 125600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3086
timestamp 1757982896
transform 1 0 127100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3087
timestamp 1757982896
transform 1 0 128600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3088
timestamp 1757982896
transform 1 0 130100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3089
timestamp 1757982896
transform 1 0 131600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3090
timestamp 1757982896
transform 1 0 133100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3091
timestamp 1757982896
transform 1 0 134600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3092
timestamp 1757982896
transform 1 0 136100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3093
timestamp 1757982896
transform 1 0 137600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3094
timestamp 1757982896
transform 1 0 139100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3095
timestamp 1757982896
transform 1 0 140600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3096
timestamp 1757982896
transform 1 0 142100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3097
timestamp 1757982896
transform 1 0 143600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3098
timestamp 1757982896
transform 1 0 145100 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3099
timestamp 1757982896
transform 1 0 146600 0 1 -43650
box 1820 -1430 3480 230
use pixel  pixel_3100
timestamp 1757982896
transform 1 0 -1900 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3101
timestamp 1757982896
transform 1 0 -400 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3102
timestamp 1757982896
transform 1 0 1100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3103
timestamp 1757982896
transform 1 0 2600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3104
timestamp 1757982896
transform 1 0 4100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3105
timestamp 1757982896
transform 1 0 5600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3106
timestamp 1757982896
transform 1 0 7100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3107
timestamp 1757982896
transform 1 0 8600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3108
timestamp 1757982896
transform 1 0 10100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3109
timestamp 1757982896
transform 1 0 11600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3110
timestamp 1757982896
transform 1 0 13100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3111
timestamp 1757982896
transform 1 0 14600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3112
timestamp 1757982896
transform 1 0 16100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3113
timestamp 1757982896
transform 1 0 17600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3114
timestamp 1757982896
transform 1 0 19100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3115
timestamp 1757982896
transform 1 0 20600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3116
timestamp 1757982896
transform 1 0 22100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3117
timestamp 1757982896
transform 1 0 23600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3118
timestamp 1757982896
transform 1 0 25100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3119
timestamp 1757982896
transform 1 0 26600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3120
timestamp 1757982896
transform 1 0 28100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3121
timestamp 1757982896
transform 1 0 29600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3122
timestamp 1757982896
transform 1 0 31100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3123
timestamp 1757982896
transform 1 0 32600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3124
timestamp 1757982896
transform 1 0 34100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3125
timestamp 1757982896
transform 1 0 35600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3126
timestamp 1757982896
transform 1 0 37100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3127
timestamp 1757982896
transform 1 0 38600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3128
timestamp 1757982896
transform 1 0 40100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3129
timestamp 1757982896
transform 1 0 41600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3130
timestamp 1757982896
transform 1 0 43100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3131
timestamp 1757982896
transform 1 0 44600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3132
timestamp 1757982896
transform 1 0 46100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3133
timestamp 1757982896
transform 1 0 47600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3134
timestamp 1757982896
transform 1 0 49100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3135
timestamp 1757982896
transform 1 0 50600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3136
timestamp 1757982896
transform 1 0 52100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3137
timestamp 1757982896
transform 1 0 53600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3138
timestamp 1757982896
transform 1 0 55100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3139
timestamp 1757982896
transform 1 0 56600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3140
timestamp 1757982896
transform 1 0 58100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3141
timestamp 1757982896
transform 1 0 59600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3142
timestamp 1757982896
transform 1 0 61100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3143
timestamp 1757982896
transform 1 0 62600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3144
timestamp 1757982896
transform 1 0 64100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3145
timestamp 1757982896
transform 1 0 65600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3146
timestamp 1757982896
transform 1 0 67100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3147
timestamp 1757982896
transform 1 0 68600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3148
timestamp 1757982896
transform 1 0 70100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3149
timestamp 1757982896
transform 1 0 71600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3150
timestamp 1757982896
transform 1 0 73100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3151
timestamp 1757982896
transform 1 0 74600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3152
timestamp 1757982896
transform 1 0 76100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3153
timestamp 1757982896
transform 1 0 77600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3154
timestamp 1757982896
transform 1 0 79100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3155
timestamp 1757982896
transform 1 0 80600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3156
timestamp 1757982896
transform 1 0 82100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3157
timestamp 1757982896
transform 1 0 83600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3158
timestamp 1757982896
transform 1 0 85100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3159
timestamp 1757982896
transform 1 0 86600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3160
timestamp 1757982896
transform 1 0 88100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3161
timestamp 1757982896
transform 1 0 89600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3162
timestamp 1757982896
transform 1 0 91100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3163
timestamp 1757982896
transform 1 0 92600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3164
timestamp 1757982896
transform 1 0 94100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3165
timestamp 1757982896
transform 1 0 95600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3166
timestamp 1757982896
transform 1 0 97100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3167
timestamp 1757982896
transform 1 0 98600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3168
timestamp 1757982896
transform 1 0 100100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3169
timestamp 1757982896
transform 1 0 101600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3170
timestamp 1757982896
transform 1 0 103100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3171
timestamp 1757982896
transform 1 0 104600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3172
timestamp 1757982896
transform 1 0 106100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3173
timestamp 1757982896
transform 1 0 107600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3174
timestamp 1757982896
transform 1 0 109100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3175
timestamp 1757982896
transform 1 0 110600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3176
timestamp 1757982896
transform 1 0 112100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3177
timestamp 1757982896
transform 1 0 113600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3178
timestamp 1757982896
transform 1 0 115100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3179
timestamp 1757982896
transform 1 0 116600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3180
timestamp 1757982896
transform 1 0 118100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3181
timestamp 1757982896
transform 1 0 119600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3182
timestamp 1757982896
transform 1 0 121100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3183
timestamp 1757982896
transform 1 0 122600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3184
timestamp 1757982896
transform 1 0 124100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3185
timestamp 1757982896
transform 1 0 125600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3186
timestamp 1757982896
transform 1 0 127100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3187
timestamp 1757982896
transform 1 0 128600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3188
timestamp 1757982896
transform 1 0 130100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3189
timestamp 1757982896
transform 1 0 131600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3190
timestamp 1757982896
transform 1 0 133100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3191
timestamp 1757982896
transform 1 0 134600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3192
timestamp 1757982896
transform 1 0 136100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3193
timestamp 1757982896
transform 1 0 137600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3194
timestamp 1757982896
transform 1 0 139100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3195
timestamp 1757982896
transform 1 0 140600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3196
timestamp 1757982896
transform 1 0 142100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3197
timestamp 1757982896
transform 1 0 143600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3198
timestamp 1757982896
transform 1 0 145100 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3199
timestamp 1757982896
transform 1 0 146600 0 1 -45150
box 1820 -1430 3480 230
use pixel  pixel_3200
timestamp 1757982896
transform 1 0 -1900 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3201
timestamp 1757982896
transform 1 0 -400 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3202
timestamp 1757982896
transform 1 0 1100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3203
timestamp 1757982896
transform 1 0 2600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3204
timestamp 1757982896
transform 1 0 4100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3205
timestamp 1757982896
transform 1 0 5600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3206
timestamp 1757982896
transform 1 0 7100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3207
timestamp 1757982896
transform 1 0 8600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3208
timestamp 1757982896
transform 1 0 10100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3209
timestamp 1757982896
transform 1 0 11600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3210
timestamp 1757982896
transform 1 0 13100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3211
timestamp 1757982896
transform 1 0 14600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3212
timestamp 1757982896
transform 1 0 16100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3213
timestamp 1757982896
transform 1 0 17600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3214
timestamp 1757982896
transform 1 0 19100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3215
timestamp 1757982896
transform 1 0 20600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3216
timestamp 1757982896
transform 1 0 22100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3217
timestamp 1757982896
transform 1 0 23600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3218
timestamp 1757982896
transform 1 0 25100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3219
timestamp 1757982896
transform 1 0 26600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3220
timestamp 1757982896
transform 1 0 28100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3221
timestamp 1757982896
transform 1 0 29600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3222
timestamp 1757982896
transform 1 0 31100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3223
timestamp 1757982896
transform 1 0 32600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3224
timestamp 1757982896
transform 1 0 34100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3225
timestamp 1757982896
transform 1 0 35600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3226
timestamp 1757982896
transform 1 0 37100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3227
timestamp 1757982896
transform 1 0 38600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3228
timestamp 1757982896
transform 1 0 40100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3229
timestamp 1757982896
transform 1 0 41600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3230
timestamp 1757982896
transform 1 0 43100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3231
timestamp 1757982896
transform 1 0 44600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3232
timestamp 1757982896
transform 1 0 46100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3233
timestamp 1757982896
transform 1 0 47600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3234
timestamp 1757982896
transform 1 0 49100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3235
timestamp 1757982896
transform 1 0 50600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3236
timestamp 1757982896
transform 1 0 52100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3237
timestamp 1757982896
transform 1 0 53600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3238
timestamp 1757982896
transform 1 0 55100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3239
timestamp 1757982896
transform 1 0 56600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3240
timestamp 1757982896
transform 1 0 58100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3241
timestamp 1757982896
transform 1 0 59600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3242
timestamp 1757982896
transform 1 0 61100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3243
timestamp 1757982896
transform 1 0 62600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3244
timestamp 1757982896
transform 1 0 64100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3245
timestamp 1757982896
transform 1 0 65600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3246
timestamp 1757982896
transform 1 0 67100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3247
timestamp 1757982896
transform 1 0 68600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3248
timestamp 1757982896
transform 1 0 70100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3249
timestamp 1757982896
transform 1 0 71600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3250
timestamp 1757982896
transform 1 0 73100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3251
timestamp 1757982896
transform 1 0 74600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3252
timestamp 1757982896
transform 1 0 76100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3253
timestamp 1757982896
transform 1 0 77600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3254
timestamp 1757982896
transform 1 0 79100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3255
timestamp 1757982896
transform 1 0 80600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3256
timestamp 1757982896
transform 1 0 82100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3257
timestamp 1757982896
transform 1 0 83600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3258
timestamp 1757982896
transform 1 0 85100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3259
timestamp 1757982896
transform 1 0 86600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3260
timestamp 1757982896
transform 1 0 88100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3261
timestamp 1757982896
transform 1 0 89600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3262
timestamp 1757982896
transform 1 0 91100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3263
timestamp 1757982896
transform 1 0 92600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3264
timestamp 1757982896
transform 1 0 94100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3265
timestamp 1757982896
transform 1 0 95600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3266
timestamp 1757982896
transform 1 0 97100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3267
timestamp 1757982896
transform 1 0 98600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3268
timestamp 1757982896
transform 1 0 100100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3269
timestamp 1757982896
transform 1 0 101600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3270
timestamp 1757982896
transform 1 0 103100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3271
timestamp 1757982896
transform 1 0 104600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3272
timestamp 1757982896
transform 1 0 106100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3273
timestamp 1757982896
transform 1 0 107600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3274
timestamp 1757982896
transform 1 0 109100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3275
timestamp 1757982896
transform 1 0 110600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3276
timestamp 1757982896
transform 1 0 112100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3277
timestamp 1757982896
transform 1 0 113600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3278
timestamp 1757982896
transform 1 0 115100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3279
timestamp 1757982896
transform 1 0 116600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3280
timestamp 1757982896
transform 1 0 118100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3281
timestamp 1757982896
transform 1 0 119600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3282
timestamp 1757982896
transform 1 0 121100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3283
timestamp 1757982896
transform 1 0 122600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3284
timestamp 1757982896
transform 1 0 124100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3285
timestamp 1757982896
transform 1 0 125600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3286
timestamp 1757982896
transform 1 0 127100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3287
timestamp 1757982896
transform 1 0 128600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3288
timestamp 1757982896
transform 1 0 130100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3289
timestamp 1757982896
transform 1 0 131600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3290
timestamp 1757982896
transform 1 0 133100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3291
timestamp 1757982896
transform 1 0 134600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3292
timestamp 1757982896
transform 1 0 136100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3293
timestamp 1757982896
transform 1 0 137600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3294
timestamp 1757982896
transform 1 0 139100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3295
timestamp 1757982896
transform 1 0 140600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3296
timestamp 1757982896
transform 1 0 142100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3297
timestamp 1757982896
transform 1 0 143600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3298
timestamp 1757982896
transform 1 0 145100 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3299
timestamp 1757982896
transform 1 0 146600 0 1 -46650
box 1820 -1430 3480 230
use pixel  pixel_3300
timestamp 1757982896
transform 1 0 -1900 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3301
timestamp 1757982896
transform 1 0 -400 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3302
timestamp 1757982896
transform 1 0 1100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3303
timestamp 1757982896
transform 1 0 2600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3304
timestamp 1757982896
transform 1 0 4100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3305
timestamp 1757982896
transform 1 0 5600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3306
timestamp 1757982896
transform 1 0 7100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3307
timestamp 1757982896
transform 1 0 8600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3308
timestamp 1757982896
transform 1 0 10100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3309
timestamp 1757982896
transform 1 0 11600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3310
timestamp 1757982896
transform 1 0 13100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3311
timestamp 1757982896
transform 1 0 14600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3312
timestamp 1757982896
transform 1 0 16100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3313
timestamp 1757982896
transform 1 0 17600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3314
timestamp 1757982896
transform 1 0 19100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3315
timestamp 1757982896
transform 1 0 20600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3316
timestamp 1757982896
transform 1 0 22100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3317
timestamp 1757982896
transform 1 0 23600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3318
timestamp 1757982896
transform 1 0 25100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3319
timestamp 1757982896
transform 1 0 26600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3320
timestamp 1757982896
transform 1 0 28100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3321
timestamp 1757982896
transform 1 0 29600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3322
timestamp 1757982896
transform 1 0 31100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3323
timestamp 1757982896
transform 1 0 32600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3324
timestamp 1757982896
transform 1 0 34100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3325
timestamp 1757982896
transform 1 0 35600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3326
timestamp 1757982896
transform 1 0 37100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3327
timestamp 1757982896
transform 1 0 38600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3328
timestamp 1757982896
transform 1 0 40100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3329
timestamp 1757982896
transform 1 0 41600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3330
timestamp 1757982896
transform 1 0 43100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3331
timestamp 1757982896
transform 1 0 44600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3332
timestamp 1757982896
transform 1 0 46100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3333
timestamp 1757982896
transform 1 0 47600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3334
timestamp 1757982896
transform 1 0 49100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3335
timestamp 1757982896
transform 1 0 50600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3336
timestamp 1757982896
transform 1 0 52100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3337
timestamp 1757982896
transform 1 0 53600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3338
timestamp 1757982896
transform 1 0 55100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3339
timestamp 1757982896
transform 1 0 56600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3340
timestamp 1757982896
transform 1 0 58100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3341
timestamp 1757982896
transform 1 0 59600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3342
timestamp 1757982896
transform 1 0 61100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3343
timestamp 1757982896
transform 1 0 62600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3344
timestamp 1757982896
transform 1 0 64100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3345
timestamp 1757982896
transform 1 0 65600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3346
timestamp 1757982896
transform 1 0 67100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3347
timestamp 1757982896
transform 1 0 68600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3348
timestamp 1757982896
transform 1 0 70100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3349
timestamp 1757982896
transform 1 0 71600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3350
timestamp 1757982896
transform 1 0 73100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3351
timestamp 1757982896
transform 1 0 74600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3352
timestamp 1757982896
transform 1 0 76100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3353
timestamp 1757982896
transform 1 0 77600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3354
timestamp 1757982896
transform 1 0 79100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3355
timestamp 1757982896
transform 1 0 80600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3356
timestamp 1757982896
transform 1 0 82100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3357
timestamp 1757982896
transform 1 0 83600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3358
timestamp 1757982896
transform 1 0 85100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3359
timestamp 1757982896
transform 1 0 86600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3360
timestamp 1757982896
transform 1 0 88100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3361
timestamp 1757982896
transform 1 0 89600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3362
timestamp 1757982896
transform 1 0 91100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3363
timestamp 1757982896
transform 1 0 92600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3364
timestamp 1757982896
transform 1 0 94100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3365
timestamp 1757982896
transform 1 0 95600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3366
timestamp 1757982896
transform 1 0 97100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3367
timestamp 1757982896
transform 1 0 98600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3368
timestamp 1757982896
transform 1 0 100100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3369
timestamp 1757982896
transform 1 0 101600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3370
timestamp 1757982896
transform 1 0 103100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3371
timestamp 1757982896
transform 1 0 104600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3372
timestamp 1757982896
transform 1 0 106100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3373
timestamp 1757982896
transform 1 0 107600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3374
timestamp 1757982896
transform 1 0 109100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3375
timestamp 1757982896
transform 1 0 110600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3376
timestamp 1757982896
transform 1 0 112100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3377
timestamp 1757982896
transform 1 0 113600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3378
timestamp 1757982896
transform 1 0 115100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3379
timestamp 1757982896
transform 1 0 116600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3380
timestamp 1757982896
transform 1 0 118100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3381
timestamp 1757982896
transform 1 0 119600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3382
timestamp 1757982896
transform 1 0 121100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3383
timestamp 1757982896
transform 1 0 122600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3384
timestamp 1757982896
transform 1 0 124100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3385
timestamp 1757982896
transform 1 0 125600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3386
timestamp 1757982896
transform 1 0 127100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3387
timestamp 1757982896
transform 1 0 128600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3388
timestamp 1757982896
transform 1 0 130100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3389
timestamp 1757982896
transform 1 0 131600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3390
timestamp 1757982896
transform 1 0 133100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3391
timestamp 1757982896
transform 1 0 134600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3392
timestamp 1757982896
transform 1 0 136100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3393
timestamp 1757982896
transform 1 0 137600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3394
timestamp 1757982896
transform 1 0 139100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3395
timestamp 1757982896
transform 1 0 140600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3396
timestamp 1757982896
transform 1 0 142100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3397
timestamp 1757982896
transform 1 0 143600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3398
timestamp 1757982896
transform 1 0 145100 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3399
timestamp 1757982896
transform 1 0 146600 0 1 -48150
box 1820 -1430 3480 230
use pixel  pixel_3400
timestamp 1757982896
transform 1 0 -1900 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3401
timestamp 1757982896
transform 1 0 -400 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3402
timestamp 1757982896
transform 1 0 1100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3403
timestamp 1757982896
transform 1 0 2600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3404
timestamp 1757982896
transform 1 0 4100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3405
timestamp 1757982896
transform 1 0 5600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3406
timestamp 1757982896
transform 1 0 7100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3407
timestamp 1757982896
transform 1 0 8600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3408
timestamp 1757982896
transform 1 0 10100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3409
timestamp 1757982896
transform 1 0 11600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3410
timestamp 1757982896
transform 1 0 13100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3411
timestamp 1757982896
transform 1 0 14600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3412
timestamp 1757982896
transform 1 0 16100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3413
timestamp 1757982896
transform 1 0 17600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3414
timestamp 1757982896
transform 1 0 19100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3415
timestamp 1757982896
transform 1 0 20600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3416
timestamp 1757982896
transform 1 0 22100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3417
timestamp 1757982896
transform 1 0 23600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3418
timestamp 1757982896
transform 1 0 25100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3419
timestamp 1757982896
transform 1 0 26600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3420
timestamp 1757982896
transform 1 0 28100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3421
timestamp 1757982896
transform 1 0 29600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3422
timestamp 1757982896
transform 1 0 31100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3423
timestamp 1757982896
transform 1 0 32600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3424
timestamp 1757982896
transform 1 0 34100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3425
timestamp 1757982896
transform 1 0 35600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3426
timestamp 1757982896
transform 1 0 37100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3427
timestamp 1757982896
transform 1 0 38600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3428
timestamp 1757982896
transform 1 0 40100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3429
timestamp 1757982896
transform 1 0 41600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3430
timestamp 1757982896
transform 1 0 43100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3431
timestamp 1757982896
transform 1 0 44600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3432
timestamp 1757982896
transform 1 0 46100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3433
timestamp 1757982896
transform 1 0 47600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3434
timestamp 1757982896
transform 1 0 49100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3435
timestamp 1757982896
transform 1 0 50600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3436
timestamp 1757982896
transform 1 0 52100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3437
timestamp 1757982896
transform 1 0 53600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3438
timestamp 1757982896
transform 1 0 55100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3439
timestamp 1757982896
transform 1 0 56600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3440
timestamp 1757982896
transform 1 0 58100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3441
timestamp 1757982896
transform 1 0 59600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3442
timestamp 1757982896
transform 1 0 61100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3443
timestamp 1757982896
transform 1 0 62600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3444
timestamp 1757982896
transform 1 0 64100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3445
timestamp 1757982896
transform 1 0 65600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3446
timestamp 1757982896
transform 1 0 67100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3447
timestamp 1757982896
transform 1 0 68600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3448
timestamp 1757982896
transform 1 0 70100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3449
timestamp 1757982896
transform 1 0 71600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3450
timestamp 1757982896
transform 1 0 73100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3451
timestamp 1757982896
transform 1 0 74600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3452
timestamp 1757982896
transform 1 0 76100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3453
timestamp 1757982896
transform 1 0 77600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3454
timestamp 1757982896
transform 1 0 79100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3455
timestamp 1757982896
transform 1 0 80600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3456
timestamp 1757982896
transform 1 0 82100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3457
timestamp 1757982896
transform 1 0 83600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3458
timestamp 1757982896
transform 1 0 85100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3459
timestamp 1757982896
transform 1 0 86600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3460
timestamp 1757982896
transform 1 0 88100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3461
timestamp 1757982896
transform 1 0 89600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3462
timestamp 1757982896
transform 1 0 91100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3463
timestamp 1757982896
transform 1 0 92600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3464
timestamp 1757982896
transform 1 0 94100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3465
timestamp 1757982896
transform 1 0 95600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3466
timestamp 1757982896
transform 1 0 97100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3467
timestamp 1757982896
transform 1 0 98600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3468
timestamp 1757982896
transform 1 0 100100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3469
timestamp 1757982896
transform 1 0 101600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3470
timestamp 1757982896
transform 1 0 103100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3471
timestamp 1757982896
transform 1 0 104600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3472
timestamp 1757982896
transform 1 0 106100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3473
timestamp 1757982896
transform 1 0 107600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3474
timestamp 1757982896
transform 1 0 109100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3475
timestamp 1757982896
transform 1 0 110600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3476
timestamp 1757982896
transform 1 0 112100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3477
timestamp 1757982896
transform 1 0 113600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3478
timestamp 1757982896
transform 1 0 115100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3479
timestamp 1757982896
transform 1 0 116600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3480
timestamp 1757982896
transform 1 0 118100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3481
timestamp 1757982896
transform 1 0 119600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3482
timestamp 1757982896
transform 1 0 121100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3483
timestamp 1757982896
transform 1 0 122600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3484
timestamp 1757982896
transform 1 0 124100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3485
timestamp 1757982896
transform 1 0 125600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3486
timestamp 1757982896
transform 1 0 127100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3487
timestamp 1757982896
transform 1 0 128600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3488
timestamp 1757982896
transform 1 0 130100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3489
timestamp 1757982896
transform 1 0 131600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3490
timestamp 1757982896
transform 1 0 133100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3491
timestamp 1757982896
transform 1 0 134600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3492
timestamp 1757982896
transform 1 0 136100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3493
timestamp 1757982896
transform 1 0 137600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3494
timestamp 1757982896
transform 1 0 139100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3495
timestamp 1757982896
transform 1 0 140600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3496
timestamp 1757982896
transform 1 0 142100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3497
timestamp 1757982896
transform 1 0 143600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3498
timestamp 1757982896
transform 1 0 145100 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3499
timestamp 1757982896
transform 1 0 146600 0 1 -49650
box 1820 -1430 3480 230
use pixel  pixel_3500
timestamp 1757982896
transform 1 0 -1900 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3501
timestamp 1757982896
transform 1 0 -400 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3502
timestamp 1757982896
transform 1 0 1100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3503
timestamp 1757982896
transform 1 0 2600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3504
timestamp 1757982896
transform 1 0 4100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3505
timestamp 1757982896
transform 1 0 5600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3506
timestamp 1757982896
transform 1 0 7100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3507
timestamp 1757982896
transform 1 0 8600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3508
timestamp 1757982896
transform 1 0 10100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3509
timestamp 1757982896
transform 1 0 11600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3510
timestamp 1757982896
transform 1 0 13100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3511
timestamp 1757982896
transform 1 0 14600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3512
timestamp 1757982896
transform 1 0 16100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3513
timestamp 1757982896
transform 1 0 17600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3514
timestamp 1757982896
transform 1 0 19100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3515
timestamp 1757982896
transform 1 0 20600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3516
timestamp 1757982896
transform 1 0 22100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3517
timestamp 1757982896
transform 1 0 23600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3518
timestamp 1757982896
transform 1 0 25100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3519
timestamp 1757982896
transform 1 0 26600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3520
timestamp 1757982896
transform 1 0 28100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3521
timestamp 1757982896
transform 1 0 29600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3522
timestamp 1757982896
transform 1 0 31100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3523
timestamp 1757982896
transform 1 0 32600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3524
timestamp 1757982896
transform 1 0 34100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3525
timestamp 1757982896
transform 1 0 35600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3526
timestamp 1757982896
transform 1 0 37100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3527
timestamp 1757982896
transform 1 0 38600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3528
timestamp 1757982896
transform 1 0 40100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3529
timestamp 1757982896
transform 1 0 41600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3530
timestamp 1757982896
transform 1 0 43100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3531
timestamp 1757982896
transform 1 0 44600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3532
timestamp 1757982896
transform 1 0 46100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3533
timestamp 1757982896
transform 1 0 47600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3534
timestamp 1757982896
transform 1 0 49100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3535
timestamp 1757982896
transform 1 0 50600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3536
timestamp 1757982896
transform 1 0 52100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3537
timestamp 1757982896
transform 1 0 53600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3538
timestamp 1757982896
transform 1 0 55100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3539
timestamp 1757982896
transform 1 0 56600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3540
timestamp 1757982896
transform 1 0 58100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3541
timestamp 1757982896
transform 1 0 59600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3542
timestamp 1757982896
transform 1 0 61100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3543
timestamp 1757982896
transform 1 0 62600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3544
timestamp 1757982896
transform 1 0 64100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3545
timestamp 1757982896
transform 1 0 65600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3546
timestamp 1757982896
transform 1 0 67100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3547
timestamp 1757982896
transform 1 0 68600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3548
timestamp 1757982896
transform 1 0 70100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3549
timestamp 1757982896
transform 1 0 71600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3550
timestamp 1757982896
transform 1 0 73100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3551
timestamp 1757982896
transform 1 0 74600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3552
timestamp 1757982896
transform 1 0 76100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3553
timestamp 1757982896
transform 1 0 77600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3554
timestamp 1757982896
transform 1 0 79100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3555
timestamp 1757982896
transform 1 0 80600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3556
timestamp 1757982896
transform 1 0 82100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3557
timestamp 1757982896
transform 1 0 83600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3558
timestamp 1757982896
transform 1 0 85100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3559
timestamp 1757982896
transform 1 0 86600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3560
timestamp 1757982896
transform 1 0 88100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3561
timestamp 1757982896
transform 1 0 89600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3562
timestamp 1757982896
transform 1 0 91100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3563
timestamp 1757982896
transform 1 0 92600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3564
timestamp 1757982896
transform 1 0 94100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3565
timestamp 1757982896
transform 1 0 95600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3566
timestamp 1757982896
transform 1 0 97100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3567
timestamp 1757982896
transform 1 0 98600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3568
timestamp 1757982896
transform 1 0 100100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3569
timestamp 1757982896
transform 1 0 101600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3570
timestamp 1757982896
transform 1 0 103100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3571
timestamp 1757982896
transform 1 0 104600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3572
timestamp 1757982896
transform 1 0 106100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3573
timestamp 1757982896
transform 1 0 107600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3574
timestamp 1757982896
transform 1 0 109100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3575
timestamp 1757982896
transform 1 0 110600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3576
timestamp 1757982896
transform 1 0 112100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3577
timestamp 1757982896
transform 1 0 113600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3578
timestamp 1757982896
transform 1 0 115100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3579
timestamp 1757982896
transform 1 0 116600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3580
timestamp 1757982896
transform 1 0 118100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3581
timestamp 1757982896
transform 1 0 119600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3582
timestamp 1757982896
transform 1 0 121100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3583
timestamp 1757982896
transform 1 0 122600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3584
timestamp 1757982896
transform 1 0 124100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3585
timestamp 1757982896
transform 1 0 125600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3586
timestamp 1757982896
transform 1 0 127100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3587
timestamp 1757982896
transform 1 0 128600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3588
timestamp 1757982896
transform 1 0 130100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3589
timestamp 1757982896
transform 1 0 131600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3590
timestamp 1757982896
transform 1 0 133100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3591
timestamp 1757982896
transform 1 0 134600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3592
timestamp 1757982896
transform 1 0 136100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3593
timestamp 1757982896
transform 1 0 137600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3594
timestamp 1757982896
transform 1 0 139100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3595
timestamp 1757982896
transform 1 0 140600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3596
timestamp 1757982896
transform 1 0 142100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3597
timestamp 1757982896
transform 1 0 143600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3598
timestamp 1757982896
transform 1 0 145100 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3599
timestamp 1757982896
transform 1 0 146600 0 1 -51150
box 1820 -1430 3480 230
use pixel  pixel_3600
timestamp 1757982896
transform 1 0 -1900 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3601
timestamp 1757982896
transform 1 0 -400 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3602
timestamp 1757982896
transform 1 0 1100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3603
timestamp 1757982896
transform 1 0 2600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3604
timestamp 1757982896
transform 1 0 4100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3605
timestamp 1757982896
transform 1 0 5600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3606
timestamp 1757982896
transform 1 0 7100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3607
timestamp 1757982896
transform 1 0 8600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3608
timestamp 1757982896
transform 1 0 10100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3609
timestamp 1757982896
transform 1 0 11600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3610
timestamp 1757982896
transform 1 0 13100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3611
timestamp 1757982896
transform 1 0 14600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3612
timestamp 1757982896
transform 1 0 16100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3613
timestamp 1757982896
transform 1 0 17600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3614
timestamp 1757982896
transform 1 0 19100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3615
timestamp 1757982896
transform 1 0 20600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3616
timestamp 1757982896
transform 1 0 22100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3617
timestamp 1757982896
transform 1 0 23600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3618
timestamp 1757982896
transform 1 0 25100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3619
timestamp 1757982896
transform 1 0 26600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3620
timestamp 1757982896
transform 1 0 28100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3621
timestamp 1757982896
transform 1 0 29600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3622
timestamp 1757982896
transform 1 0 31100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3623
timestamp 1757982896
transform 1 0 32600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3624
timestamp 1757982896
transform 1 0 34100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3625
timestamp 1757982896
transform 1 0 35600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3626
timestamp 1757982896
transform 1 0 37100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3627
timestamp 1757982896
transform 1 0 38600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3628
timestamp 1757982896
transform 1 0 40100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3629
timestamp 1757982896
transform 1 0 41600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3630
timestamp 1757982896
transform 1 0 43100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3631
timestamp 1757982896
transform 1 0 44600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3632
timestamp 1757982896
transform 1 0 46100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3633
timestamp 1757982896
transform 1 0 47600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3634
timestamp 1757982896
transform 1 0 49100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3635
timestamp 1757982896
transform 1 0 50600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3636
timestamp 1757982896
transform 1 0 52100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3637
timestamp 1757982896
transform 1 0 53600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3638
timestamp 1757982896
transform 1 0 55100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3639
timestamp 1757982896
transform 1 0 56600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3640
timestamp 1757982896
transform 1 0 58100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3641
timestamp 1757982896
transform 1 0 59600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3642
timestamp 1757982896
transform 1 0 61100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3643
timestamp 1757982896
transform 1 0 62600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3644
timestamp 1757982896
transform 1 0 64100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3645
timestamp 1757982896
transform 1 0 65600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3646
timestamp 1757982896
transform 1 0 67100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3647
timestamp 1757982896
transform 1 0 68600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3648
timestamp 1757982896
transform 1 0 70100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3649
timestamp 1757982896
transform 1 0 71600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3650
timestamp 1757982896
transform 1 0 73100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3651
timestamp 1757982896
transform 1 0 74600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3652
timestamp 1757982896
transform 1 0 76100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3653
timestamp 1757982896
transform 1 0 77600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3654
timestamp 1757982896
transform 1 0 79100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3655
timestamp 1757982896
transform 1 0 80600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3656
timestamp 1757982896
transform 1 0 82100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3657
timestamp 1757982896
transform 1 0 83600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3658
timestamp 1757982896
transform 1 0 85100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3659
timestamp 1757982896
transform 1 0 86600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3660
timestamp 1757982896
transform 1 0 88100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3661
timestamp 1757982896
transform 1 0 89600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3662
timestamp 1757982896
transform 1 0 91100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3663
timestamp 1757982896
transform 1 0 92600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3664
timestamp 1757982896
transform 1 0 94100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3665
timestamp 1757982896
transform 1 0 95600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3666
timestamp 1757982896
transform 1 0 97100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3667
timestamp 1757982896
transform 1 0 98600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3668
timestamp 1757982896
transform 1 0 100100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3669
timestamp 1757982896
transform 1 0 101600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3670
timestamp 1757982896
transform 1 0 103100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3671
timestamp 1757982896
transform 1 0 104600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3672
timestamp 1757982896
transform 1 0 106100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3673
timestamp 1757982896
transform 1 0 107600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3674
timestamp 1757982896
transform 1 0 109100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3675
timestamp 1757982896
transform 1 0 110600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3676
timestamp 1757982896
transform 1 0 112100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3677
timestamp 1757982896
transform 1 0 113600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3678
timestamp 1757982896
transform 1 0 115100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3679
timestamp 1757982896
transform 1 0 116600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3680
timestamp 1757982896
transform 1 0 118100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3681
timestamp 1757982896
transform 1 0 119600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3682
timestamp 1757982896
transform 1 0 121100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3683
timestamp 1757982896
transform 1 0 122600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3684
timestamp 1757982896
transform 1 0 124100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3685
timestamp 1757982896
transform 1 0 125600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3686
timestamp 1757982896
transform 1 0 127100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3687
timestamp 1757982896
transform 1 0 128600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3688
timestamp 1757982896
transform 1 0 130100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3689
timestamp 1757982896
transform 1 0 131600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3690
timestamp 1757982896
transform 1 0 133100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3691
timestamp 1757982896
transform 1 0 134600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3692
timestamp 1757982896
transform 1 0 136100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3693
timestamp 1757982896
transform 1 0 137600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3694
timestamp 1757982896
transform 1 0 139100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3695
timestamp 1757982896
transform 1 0 140600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3696
timestamp 1757982896
transform 1 0 142100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3697
timestamp 1757982896
transform 1 0 143600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3698
timestamp 1757982896
transform 1 0 145100 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3699
timestamp 1757982896
transform 1 0 146600 0 1 -52650
box 1820 -1430 3480 230
use pixel  pixel_3700
timestamp 1757982896
transform 1 0 -1900 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3701
timestamp 1757982896
transform 1 0 -400 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3702
timestamp 1757982896
transform 1 0 1100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3703
timestamp 1757982896
transform 1 0 2600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3704
timestamp 1757982896
transform 1 0 4100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3705
timestamp 1757982896
transform 1 0 5600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3706
timestamp 1757982896
transform 1 0 7100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3707
timestamp 1757982896
transform 1 0 8600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3708
timestamp 1757982896
transform 1 0 10100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3709
timestamp 1757982896
transform 1 0 11600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3710
timestamp 1757982896
transform 1 0 13100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3711
timestamp 1757982896
transform 1 0 14600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3712
timestamp 1757982896
transform 1 0 16100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3713
timestamp 1757982896
transform 1 0 17600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3714
timestamp 1757982896
transform 1 0 19100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3715
timestamp 1757982896
transform 1 0 20600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3716
timestamp 1757982896
transform 1 0 22100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3717
timestamp 1757982896
transform 1 0 23600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3718
timestamp 1757982896
transform 1 0 25100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3719
timestamp 1757982896
transform 1 0 26600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3720
timestamp 1757982896
transform 1 0 28100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3721
timestamp 1757982896
transform 1 0 29600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3722
timestamp 1757982896
transform 1 0 31100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3723
timestamp 1757982896
transform 1 0 32600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3724
timestamp 1757982896
transform 1 0 34100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3725
timestamp 1757982896
transform 1 0 35600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3726
timestamp 1757982896
transform 1 0 37100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3727
timestamp 1757982896
transform 1 0 38600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3728
timestamp 1757982896
transform 1 0 40100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3729
timestamp 1757982896
transform 1 0 41600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3730
timestamp 1757982896
transform 1 0 43100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3731
timestamp 1757982896
transform 1 0 44600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3732
timestamp 1757982896
transform 1 0 46100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3733
timestamp 1757982896
transform 1 0 47600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3734
timestamp 1757982896
transform 1 0 49100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3735
timestamp 1757982896
transform 1 0 50600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3736
timestamp 1757982896
transform 1 0 52100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3737
timestamp 1757982896
transform 1 0 53600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3738
timestamp 1757982896
transform 1 0 55100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3739
timestamp 1757982896
transform 1 0 56600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3740
timestamp 1757982896
transform 1 0 58100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3741
timestamp 1757982896
transform 1 0 59600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3742
timestamp 1757982896
transform 1 0 61100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3743
timestamp 1757982896
transform 1 0 62600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3744
timestamp 1757982896
transform 1 0 64100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3745
timestamp 1757982896
transform 1 0 65600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3746
timestamp 1757982896
transform 1 0 67100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3747
timestamp 1757982896
transform 1 0 68600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3748
timestamp 1757982896
transform 1 0 70100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3749
timestamp 1757982896
transform 1 0 71600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3750
timestamp 1757982896
transform 1 0 73100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3751
timestamp 1757982896
transform 1 0 74600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3752
timestamp 1757982896
transform 1 0 76100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3753
timestamp 1757982896
transform 1 0 77600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3754
timestamp 1757982896
transform 1 0 79100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3755
timestamp 1757982896
transform 1 0 80600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3756
timestamp 1757982896
transform 1 0 82100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3757
timestamp 1757982896
transform 1 0 83600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3758
timestamp 1757982896
transform 1 0 85100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3759
timestamp 1757982896
transform 1 0 86600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3760
timestamp 1757982896
transform 1 0 88100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3761
timestamp 1757982896
transform 1 0 89600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3762
timestamp 1757982896
transform 1 0 91100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3763
timestamp 1757982896
transform 1 0 92600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3764
timestamp 1757982896
transform 1 0 94100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3765
timestamp 1757982896
transform 1 0 95600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3766
timestamp 1757982896
transform 1 0 97100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3767
timestamp 1757982896
transform 1 0 98600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3768
timestamp 1757982896
transform 1 0 100100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3769
timestamp 1757982896
transform 1 0 101600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3770
timestamp 1757982896
transform 1 0 103100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3771
timestamp 1757982896
transform 1 0 104600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3772
timestamp 1757982896
transform 1 0 106100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3773
timestamp 1757982896
transform 1 0 107600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3774
timestamp 1757982896
transform 1 0 109100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3775
timestamp 1757982896
transform 1 0 110600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3776
timestamp 1757982896
transform 1 0 112100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3777
timestamp 1757982896
transform 1 0 113600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3778
timestamp 1757982896
transform 1 0 115100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3779
timestamp 1757982896
transform 1 0 116600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3780
timestamp 1757982896
transform 1 0 118100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3781
timestamp 1757982896
transform 1 0 119600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3782
timestamp 1757982896
transform 1 0 121100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3783
timestamp 1757982896
transform 1 0 122600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3784
timestamp 1757982896
transform 1 0 124100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3785
timestamp 1757982896
transform 1 0 125600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3786
timestamp 1757982896
transform 1 0 127100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3787
timestamp 1757982896
transform 1 0 128600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3788
timestamp 1757982896
transform 1 0 130100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3789
timestamp 1757982896
transform 1 0 131600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3790
timestamp 1757982896
transform 1 0 133100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3791
timestamp 1757982896
transform 1 0 134600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3792
timestamp 1757982896
transform 1 0 136100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3793
timestamp 1757982896
transform 1 0 137600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3794
timestamp 1757982896
transform 1 0 139100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3795
timestamp 1757982896
transform 1 0 140600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3796
timestamp 1757982896
transform 1 0 142100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3797
timestamp 1757982896
transform 1 0 143600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3798
timestamp 1757982896
transform 1 0 145100 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3799
timestamp 1757982896
transform 1 0 146600 0 1 -54150
box 1820 -1430 3480 230
use pixel  pixel_3800
timestamp 1757982896
transform 1 0 -1900 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3801
timestamp 1757982896
transform 1 0 -400 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3802
timestamp 1757982896
transform 1 0 1100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3803
timestamp 1757982896
transform 1 0 2600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3804
timestamp 1757982896
transform 1 0 4100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3805
timestamp 1757982896
transform 1 0 5600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3806
timestamp 1757982896
transform 1 0 7100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3807
timestamp 1757982896
transform 1 0 8600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3808
timestamp 1757982896
transform 1 0 10100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3809
timestamp 1757982896
transform 1 0 11600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3810
timestamp 1757982896
transform 1 0 13100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3811
timestamp 1757982896
transform 1 0 14600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3812
timestamp 1757982896
transform 1 0 16100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3813
timestamp 1757982896
transform 1 0 17600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3814
timestamp 1757982896
transform 1 0 19100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3815
timestamp 1757982896
transform 1 0 20600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3816
timestamp 1757982896
transform 1 0 22100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3817
timestamp 1757982896
transform 1 0 23600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3818
timestamp 1757982896
transform 1 0 25100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3819
timestamp 1757982896
transform 1 0 26600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3820
timestamp 1757982896
transform 1 0 28100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3821
timestamp 1757982896
transform 1 0 29600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3822
timestamp 1757982896
transform 1 0 31100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3823
timestamp 1757982896
transform 1 0 32600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3824
timestamp 1757982896
transform 1 0 34100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3825
timestamp 1757982896
transform 1 0 35600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3826
timestamp 1757982896
transform 1 0 37100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3827
timestamp 1757982896
transform 1 0 38600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3828
timestamp 1757982896
transform 1 0 40100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3829
timestamp 1757982896
transform 1 0 41600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3830
timestamp 1757982896
transform 1 0 43100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3831
timestamp 1757982896
transform 1 0 44600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3832
timestamp 1757982896
transform 1 0 46100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3833
timestamp 1757982896
transform 1 0 47600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3834
timestamp 1757982896
transform 1 0 49100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3835
timestamp 1757982896
transform 1 0 50600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3836
timestamp 1757982896
transform 1 0 52100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3837
timestamp 1757982896
transform 1 0 53600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3838
timestamp 1757982896
transform 1 0 55100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3839
timestamp 1757982896
transform 1 0 56600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3840
timestamp 1757982896
transform 1 0 58100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3841
timestamp 1757982896
transform 1 0 59600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3842
timestamp 1757982896
transform 1 0 61100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3843
timestamp 1757982896
transform 1 0 62600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3844
timestamp 1757982896
transform 1 0 64100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3845
timestamp 1757982896
transform 1 0 65600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3846
timestamp 1757982896
transform 1 0 67100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3847
timestamp 1757982896
transform 1 0 68600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3848
timestamp 1757982896
transform 1 0 70100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3849
timestamp 1757982896
transform 1 0 71600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3850
timestamp 1757982896
transform 1 0 73100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3851
timestamp 1757982896
transform 1 0 74600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3852
timestamp 1757982896
transform 1 0 76100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3853
timestamp 1757982896
transform 1 0 77600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3854
timestamp 1757982896
transform 1 0 79100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3855
timestamp 1757982896
transform 1 0 80600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3856
timestamp 1757982896
transform 1 0 82100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3857
timestamp 1757982896
transform 1 0 83600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3858
timestamp 1757982896
transform 1 0 85100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3859
timestamp 1757982896
transform 1 0 86600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3860
timestamp 1757982896
transform 1 0 88100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3861
timestamp 1757982896
transform 1 0 89600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3862
timestamp 1757982896
transform 1 0 91100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3863
timestamp 1757982896
transform 1 0 92600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3864
timestamp 1757982896
transform 1 0 94100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3865
timestamp 1757982896
transform 1 0 95600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3866
timestamp 1757982896
transform 1 0 97100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3867
timestamp 1757982896
transform 1 0 98600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3868
timestamp 1757982896
transform 1 0 100100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3869
timestamp 1757982896
transform 1 0 101600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3870
timestamp 1757982896
transform 1 0 103100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3871
timestamp 1757982896
transform 1 0 104600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3872
timestamp 1757982896
transform 1 0 106100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3873
timestamp 1757982896
transform 1 0 107600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3874
timestamp 1757982896
transform 1 0 109100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3875
timestamp 1757982896
transform 1 0 110600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3876
timestamp 1757982896
transform 1 0 112100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3877
timestamp 1757982896
transform 1 0 113600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3878
timestamp 1757982896
transform 1 0 115100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3879
timestamp 1757982896
transform 1 0 116600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3880
timestamp 1757982896
transform 1 0 118100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3881
timestamp 1757982896
transform 1 0 119600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3882
timestamp 1757982896
transform 1 0 121100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3883
timestamp 1757982896
transform 1 0 122600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3884
timestamp 1757982896
transform 1 0 124100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3885
timestamp 1757982896
transform 1 0 125600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3886
timestamp 1757982896
transform 1 0 127100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3887
timestamp 1757982896
transform 1 0 128600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3888
timestamp 1757982896
transform 1 0 130100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3889
timestamp 1757982896
transform 1 0 131600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3890
timestamp 1757982896
transform 1 0 133100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3891
timestamp 1757982896
transform 1 0 134600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3892
timestamp 1757982896
transform 1 0 136100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3893
timestamp 1757982896
transform 1 0 137600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3894
timestamp 1757982896
transform 1 0 139100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3895
timestamp 1757982896
transform 1 0 140600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3896
timestamp 1757982896
transform 1 0 142100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3897
timestamp 1757982896
transform 1 0 143600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3898
timestamp 1757982896
transform 1 0 145100 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3899
timestamp 1757982896
transform 1 0 146600 0 1 -55650
box 1820 -1430 3480 230
use pixel  pixel_3900
timestamp 1757982896
transform 1 0 -1900 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3901
timestamp 1757982896
transform 1 0 -400 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3902
timestamp 1757982896
transform 1 0 1100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3903
timestamp 1757982896
transform 1 0 2600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3904
timestamp 1757982896
transform 1 0 4100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3905
timestamp 1757982896
transform 1 0 5600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3906
timestamp 1757982896
transform 1 0 7100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3907
timestamp 1757982896
transform 1 0 8600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3908
timestamp 1757982896
transform 1 0 10100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3909
timestamp 1757982896
transform 1 0 11600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3910
timestamp 1757982896
transform 1 0 13100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3911
timestamp 1757982896
transform 1 0 14600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3912
timestamp 1757982896
transform 1 0 16100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3913
timestamp 1757982896
transform 1 0 17600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3914
timestamp 1757982896
transform 1 0 19100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3915
timestamp 1757982896
transform 1 0 20600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3916
timestamp 1757982896
transform 1 0 22100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3917
timestamp 1757982896
transform 1 0 23600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3918
timestamp 1757982896
transform 1 0 25100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3919
timestamp 1757982896
transform 1 0 26600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3920
timestamp 1757982896
transform 1 0 28100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3921
timestamp 1757982896
transform 1 0 29600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3922
timestamp 1757982896
transform 1 0 31100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3923
timestamp 1757982896
transform 1 0 32600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3924
timestamp 1757982896
transform 1 0 34100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3925
timestamp 1757982896
transform 1 0 35600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3926
timestamp 1757982896
transform 1 0 37100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3927
timestamp 1757982896
transform 1 0 38600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3928
timestamp 1757982896
transform 1 0 40100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3929
timestamp 1757982896
transform 1 0 41600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3930
timestamp 1757982896
transform 1 0 43100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3931
timestamp 1757982896
transform 1 0 44600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3932
timestamp 1757982896
transform 1 0 46100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3933
timestamp 1757982896
transform 1 0 47600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3934
timestamp 1757982896
transform 1 0 49100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3935
timestamp 1757982896
transform 1 0 50600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3936
timestamp 1757982896
transform 1 0 52100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3937
timestamp 1757982896
transform 1 0 53600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3938
timestamp 1757982896
transform 1 0 55100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3939
timestamp 1757982896
transform 1 0 56600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3940
timestamp 1757982896
transform 1 0 58100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3941
timestamp 1757982896
transform 1 0 59600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3942
timestamp 1757982896
transform 1 0 61100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3943
timestamp 1757982896
transform 1 0 62600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3944
timestamp 1757982896
transform 1 0 64100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3945
timestamp 1757982896
transform 1 0 65600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3946
timestamp 1757982896
transform 1 0 67100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3947
timestamp 1757982896
transform 1 0 68600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3948
timestamp 1757982896
transform 1 0 70100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3949
timestamp 1757982896
transform 1 0 71600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3950
timestamp 1757982896
transform 1 0 73100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3951
timestamp 1757982896
transform 1 0 74600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3952
timestamp 1757982896
transform 1 0 76100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3953
timestamp 1757982896
transform 1 0 77600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3954
timestamp 1757982896
transform 1 0 79100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3955
timestamp 1757982896
transform 1 0 80600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3956
timestamp 1757982896
transform 1 0 82100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3957
timestamp 1757982896
transform 1 0 83600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3958
timestamp 1757982896
transform 1 0 85100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3959
timestamp 1757982896
transform 1 0 86600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3960
timestamp 1757982896
transform 1 0 88100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3961
timestamp 1757982896
transform 1 0 89600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3962
timestamp 1757982896
transform 1 0 91100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3963
timestamp 1757982896
transform 1 0 92600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3964
timestamp 1757982896
transform 1 0 94100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3965
timestamp 1757982896
transform 1 0 95600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3966
timestamp 1757982896
transform 1 0 97100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3967
timestamp 1757982896
transform 1 0 98600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3968
timestamp 1757982896
transform 1 0 100100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3969
timestamp 1757982896
transform 1 0 101600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3970
timestamp 1757982896
transform 1 0 103100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3971
timestamp 1757982896
transform 1 0 104600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3972
timestamp 1757982896
transform 1 0 106100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3973
timestamp 1757982896
transform 1 0 107600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3974
timestamp 1757982896
transform 1 0 109100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3975
timestamp 1757982896
transform 1 0 110600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3976
timestamp 1757982896
transform 1 0 112100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3977
timestamp 1757982896
transform 1 0 113600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3978
timestamp 1757982896
transform 1 0 115100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3979
timestamp 1757982896
transform 1 0 116600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3980
timestamp 1757982896
transform 1 0 118100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3981
timestamp 1757982896
transform 1 0 119600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3982
timestamp 1757982896
transform 1 0 121100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3983
timestamp 1757982896
transform 1 0 122600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3984
timestamp 1757982896
transform 1 0 124100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3985
timestamp 1757982896
transform 1 0 125600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3986
timestamp 1757982896
transform 1 0 127100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3987
timestamp 1757982896
transform 1 0 128600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3988
timestamp 1757982896
transform 1 0 130100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3989
timestamp 1757982896
transform 1 0 131600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3990
timestamp 1757982896
transform 1 0 133100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3991
timestamp 1757982896
transform 1 0 134600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3992
timestamp 1757982896
transform 1 0 136100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3993
timestamp 1757982896
transform 1 0 137600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3994
timestamp 1757982896
transform 1 0 139100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3995
timestamp 1757982896
transform 1 0 140600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3996
timestamp 1757982896
transform 1 0 142100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3997
timestamp 1757982896
transform 1 0 143600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3998
timestamp 1757982896
transform 1 0 145100 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_3999
timestamp 1757982896
transform 1 0 146600 0 1 -57150
box 1820 -1430 3480 230
use pixel  pixel_4000
timestamp 1757982896
transform 1 0 -1900 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4001
timestamp 1757982896
transform 1 0 -400 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4002
timestamp 1757982896
transform 1 0 1100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4003
timestamp 1757982896
transform 1 0 2600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4004
timestamp 1757982896
transform 1 0 4100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4005
timestamp 1757982896
transform 1 0 5600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4006
timestamp 1757982896
transform 1 0 7100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4007
timestamp 1757982896
transform 1 0 8600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4008
timestamp 1757982896
transform 1 0 10100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4009
timestamp 1757982896
transform 1 0 11600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4010
timestamp 1757982896
transform 1 0 13100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4011
timestamp 1757982896
transform 1 0 14600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4012
timestamp 1757982896
transform 1 0 16100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4013
timestamp 1757982896
transform 1 0 17600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4014
timestamp 1757982896
transform 1 0 19100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4015
timestamp 1757982896
transform 1 0 20600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4016
timestamp 1757982896
transform 1 0 22100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4017
timestamp 1757982896
transform 1 0 23600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4018
timestamp 1757982896
transform 1 0 25100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4019
timestamp 1757982896
transform 1 0 26600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4020
timestamp 1757982896
transform 1 0 28100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4021
timestamp 1757982896
transform 1 0 29600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4022
timestamp 1757982896
transform 1 0 31100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4023
timestamp 1757982896
transform 1 0 32600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4024
timestamp 1757982896
transform 1 0 34100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4025
timestamp 1757982896
transform 1 0 35600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4026
timestamp 1757982896
transform 1 0 37100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4027
timestamp 1757982896
transform 1 0 38600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4028
timestamp 1757982896
transform 1 0 40100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4029
timestamp 1757982896
transform 1 0 41600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4030
timestamp 1757982896
transform 1 0 43100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4031
timestamp 1757982896
transform 1 0 44600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4032
timestamp 1757982896
transform 1 0 46100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4033
timestamp 1757982896
transform 1 0 47600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4034
timestamp 1757982896
transform 1 0 49100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4035
timestamp 1757982896
transform 1 0 50600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4036
timestamp 1757982896
transform 1 0 52100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4037
timestamp 1757982896
transform 1 0 53600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4038
timestamp 1757982896
transform 1 0 55100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4039
timestamp 1757982896
transform 1 0 56600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4040
timestamp 1757982896
transform 1 0 58100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4041
timestamp 1757982896
transform 1 0 59600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4042
timestamp 1757982896
transform 1 0 61100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4043
timestamp 1757982896
transform 1 0 62600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4044
timestamp 1757982896
transform 1 0 64100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4045
timestamp 1757982896
transform 1 0 65600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4046
timestamp 1757982896
transform 1 0 67100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4047
timestamp 1757982896
transform 1 0 68600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4048
timestamp 1757982896
transform 1 0 70100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4049
timestamp 1757982896
transform 1 0 71600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4050
timestamp 1757982896
transform 1 0 73100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4051
timestamp 1757982896
transform 1 0 74600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4052
timestamp 1757982896
transform 1 0 76100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4053
timestamp 1757982896
transform 1 0 77600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4054
timestamp 1757982896
transform 1 0 79100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4055
timestamp 1757982896
transform 1 0 80600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4056
timestamp 1757982896
transform 1 0 82100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4057
timestamp 1757982896
transform 1 0 83600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4058
timestamp 1757982896
transform 1 0 85100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4059
timestamp 1757982896
transform 1 0 86600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4060
timestamp 1757982896
transform 1 0 88100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4061
timestamp 1757982896
transform 1 0 89600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4062
timestamp 1757982896
transform 1 0 91100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4063
timestamp 1757982896
transform 1 0 92600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4064
timestamp 1757982896
transform 1 0 94100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4065
timestamp 1757982896
transform 1 0 95600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4066
timestamp 1757982896
transform 1 0 97100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4067
timestamp 1757982896
transform 1 0 98600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4068
timestamp 1757982896
transform 1 0 100100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4069
timestamp 1757982896
transform 1 0 101600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4070
timestamp 1757982896
transform 1 0 103100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4071
timestamp 1757982896
transform 1 0 104600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4072
timestamp 1757982896
transform 1 0 106100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4073
timestamp 1757982896
transform 1 0 107600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4074
timestamp 1757982896
transform 1 0 109100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4075
timestamp 1757982896
transform 1 0 110600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4076
timestamp 1757982896
transform 1 0 112100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4077
timestamp 1757982896
transform 1 0 113600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4078
timestamp 1757982896
transform 1 0 115100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4079
timestamp 1757982896
transform 1 0 116600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4080
timestamp 1757982896
transform 1 0 118100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4081
timestamp 1757982896
transform 1 0 119600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4082
timestamp 1757982896
transform 1 0 121100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4083
timestamp 1757982896
transform 1 0 122600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4084
timestamp 1757982896
transform 1 0 124100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4085
timestamp 1757982896
transform 1 0 125600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4086
timestamp 1757982896
transform 1 0 127100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4087
timestamp 1757982896
transform 1 0 128600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4088
timestamp 1757982896
transform 1 0 130100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4089
timestamp 1757982896
transform 1 0 131600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4090
timestamp 1757982896
transform 1 0 133100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4091
timestamp 1757982896
transform 1 0 134600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4092
timestamp 1757982896
transform 1 0 136100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4093
timestamp 1757982896
transform 1 0 137600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4094
timestamp 1757982896
transform 1 0 139100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4095
timestamp 1757982896
transform 1 0 140600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4096
timestamp 1757982896
transform 1 0 142100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4097
timestamp 1757982896
transform 1 0 143600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4098
timestamp 1757982896
transform 1 0 145100 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4099
timestamp 1757982896
transform 1 0 146600 0 1 -58650
box 1820 -1430 3480 230
use pixel  pixel_4100
timestamp 1757982896
transform 1 0 -1900 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4101
timestamp 1757982896
transform 1 0 -400 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4102
timestamp 1757982896
transform 1 0 1100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4103
timestamp 1757982896
transform 1 0 2600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4104
timestamp 1757982896
transform 1 0 4100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4105
timestamp 1757982896
transform 1 0 5600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4106
timestamp 1757982896
transform 1 0 7100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4107
timestamp 1757982896
transform 1 0 8600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4108
timestamp 1757982896
transform 1 0 10100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4109
timestamp 1757982896
transform 1 0 11600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4110
timestamp 1757982896
transform 1 0 13100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4111
timestamp 1757982896
transform 1 0 14600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4112
timestamp 1757982896
transform 1 0 16100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4113
timestamp 1757982896
transform 1 0 17600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4114
timestamp 1757982896
transform 1 0 19100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4115
timestamp 1757982896
transform 1 0 20600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4116
timestamp 1757982896
transform 1 0 22100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4117
timestamp 1757982896
transform 1 0 23600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4118
timestamp 1757982896
transform 1 0 25100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4119
timestamp 1757982896
transform 1 0 26600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4120
timestamp 1757982896
transform 1 0 28100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4121
timestamp 1757982896
transform 1 0 29600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4122
timestamp 1757982896
transform 1 0 31100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4123
timestamp 1757982896
transform 1 0 32600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4124
timestamp 1757982896
transform 1 0 34100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4125
timestamp 1757982896
transform 1 0 35600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4126
timestamp 1757982896
transform 1 0 37100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4127
timestamp 1757982896
transform 1 0 38600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4128
timestamp 1757982896
transform 1 0 40100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4129
timestamp 1757982896
transform 1 0 41600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4130
timestamp 1757982896
transform 1 0 43100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4131
timestamp 1757982896
transform 1 0 44600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4132
timestamp 1757982896
transform 1 0 46100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4133
timestamp 1757982896
transform 1 0 47600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4134
timestamp 1757982896
transform 1 0 49100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4135
timestamp 1757982896
transform 1 0 50600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4136
timestamp 1757982896
transform 1 0 52100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4137
timestamp 1757982896
transform 1 0 53600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4138
timestamp 1757982896
transform 1 0 55100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4139
timestamp 1757982896
transform 1 0 56600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4140
timestamp 1757982896
transform 1 0 58100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4141
timestamp 1757982896
transform 1 0 59600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4142
timestamp 1757982896
transform 1 0 61100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4143
timestamp 1757982896
transform 1 0 62600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4144
timestamp 1757982896
transform 1 0 64100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4145
timestamp 1757982896
transform 1 0 65600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4146
timestamp 1757982896
transform 1 0 67100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4147
timestamp 1757982896
transform 1 0 68600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4148
timestamp 1757982896
transform 1 0 70100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4149
timestamp 1757982896
transform 1 0 71600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4150
timestamp 1757982896
transform 1 0 73100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4151
timestamp 1757982896
transform 1 0 74600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4152
timestamp 1757982896
transform 1 0 76100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4153
timestamp 1757982896
transform 1 0 77600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4154
timestamp 1757982896
transform 1 0 79100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4155
timestamp 1757982896
transform 1 0 80600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4156
timestamp 1757982896
transform 1 0 82100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4157
timestamp 1757982896
transform 1 0 83600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4158
timestamp 1757982896
transform 1 0 85100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4159
timestamp 1757982896
transform 1 0 86600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4160
timestamp 1757982896
transform 1 0 88100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4161
timestamp 1757982896
transform 1 0 89600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4162
timestamp 1757982896
transform 1 0 91100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4163
timestamp 1757982896
transform 1 0 92600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4164
timestamp 1757982896
transform 1 0 94100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4165
timestamp 1757982896
transform 1 0 95600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4166
timestamp 1757982896
transform 1 0 97100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4167
timestamp 1757982896
transform 1 0 98600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4168
timestamp 1757982896
transform 1 0 100100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4169
timestamp 1757982896
transform 1 0 101600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4170
timestamp 1757982896
transform 1 0 103100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4171
timestamp 1757982896
transform 1 0 104600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4172
timestamp 1757982896
transform 1 0 106100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4173
timestamp 1757982896
transform 1 0 107600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4174
timestamp 1757982896
transform 1 0 109100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4175
timestamp 1757982896
transform 1 0 110600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4176
timestamp 1757982896
transform 1 0 112100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4177
timestamp 1757982896
transform 1 0 113600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4178
timestamp 1757982896
transform 1 0 115100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4179
timestamp 1757982896
transform 1 0 116600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4180
timestamp 1757982896
transform 1 0 118100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4181
timestamp 1757982896
transform 1 0 119600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4182
timestamp 1757982896
transform 1 0 121100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4183
timestamp 1757982896
transform 1 0 122600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4184
timestamp 1757982896
transform 1 0 124100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4185
timestamp 1757982896
transform 1 0 125600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4186
timestamp 1757982896
transform 1 0 127100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4187
timestamp 1757982896
transform 1 0 128600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4188
timestamp 1757982896
transform 1 0 130100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4189
timestamp 1757982896
transform 1 0 131600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4190
timestamp 1757982896
transform 1 0 133100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4191
timestamp 1757982896
transform 1 0 134600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4192
timestamp 1757982896
transform 1 0 136100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4193
timestamp 1757982896
transform 1 0 137600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4194
timestamp 1757982896
transform 1 0 139100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4195
timestamp 1757982896
transform 1 0 140600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4196
timestamp 1757982896
transform 1 0 142100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4197
timestamp 1757982896
transform 1 0 143600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4198
timestamp 1757982896
transform 1 0 145100 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4199
timestamp 1757982896
transform 1 0 146600 0 1 -60150
box 1820 -1430 3480 230
use pixel  pixel_4200
timestamp 1757982896
transform 1 0 -1900 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4201
timestamp 1757982896
transform 1 0 -400 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4202
timestamp 1757982896
transform 1 0 1100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4203
timestamp 1757982896
transform 1 0 2600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4204
timestamp 1757982896
transform 1 0 4100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4205
timestamp 1757982896
transform 1 0 5600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4206
timestamp 1757982896
transform 1 0 7100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4207
timestamp 1757982896
transform 1 0 8600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4208
timestamp 1757982896
transform 1 0 10100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4209
timestamp 1757982896
transform 1 0 11600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4210
timestamp 1757982896
transform 1 0 13100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4211
timestamp 1757982896
transform 1 0 14600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4212
timestamp 1757982896
transform 1 0 16100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4213
timestamp 1757982896
transform 1 0 17600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4214
timestamp 1757982896
transform 1 0 19100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4215
timestamp 1757982896
transform 1 0 20600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4216
timestamp 1757982896
transform 1 0 22100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4217
timestamp 1757982896
transform 1 0 23600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4218
timestamp 1757982896
transform 1 0 25100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4219
timestamp 1757982896
transform 1 0 26600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4220
timestamp 1757982896
transform 1 0 28100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4221
timestamp 1757982896
transform 1 0 29600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4222
timestamp 1757982896
transform 1 0 31100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4223
timestamp 1757982896
transform 1 0 32600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4224
timestamp 1757982896
transform 1 0 34100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4225
timestamp 1757982896
transform 1 0 35600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4226
timestamp 1757982896
transform 1 0 37100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4227
timestamp 1757982896
transform 1 0 38600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4228
timestamp 1757982896
transform 1 0 40100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4229
timestamp 1757982896
transform 1 0 41600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4230
timestamp 1757982896
transform 1 0 43100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4231
timestamp 1757982896
transform 1 0 44600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4232
timestamp 1757982896
transform 1 0 46100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4233
timestamp 1757982896
transform 1 0 47600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4234
timestamp 1757982896
transform 1 0 49100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4235
timestamp 1757982896
transform 1 0 50600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4236
timestamp 1757982896
transform 1 0 52100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4237
timestamp 1757982896
transform 1 0 53600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4238
timestamp 1757982896
transform 1 0 55100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4239
timestamp 1757982896
transform 1 0 56600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4240
timestamp 1757982896
transform 1 0 58100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4241
timestamp 1757982896
transform 1 0 59600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4242
timestamp 1757982896
transform 1 0 61100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4243
timestamp 1757982896
transform 1 0 62600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4244
timestamp 1757982896
transform 1 0 64100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4245
timestamp 1757982896
transform 1 0 65600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4246
timestamp 1757982896
transform 1 0 67100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4247
timestamp 1757982896
transform 1 0 68600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4248
timestamp 1757982896
transform 1 0 70100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4249
timestamp 1757982896
transform 1 0 71600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4250
timestamp 1757982896
transform 1 0 73100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4251
timestamp 1757982896
transform 1 0 74600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4252
timestamp 1757982896
transform 1 0 76100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4253
timestamp 1757982896
transform 1 0 77600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4254
timestamp 1757982896
transform 1 0 79100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4255
timestamp 1757982896
transform 1 0 80600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4256
timestamp 1757982896
transform 1 0 82100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4257
timestamp 1757982896
transform 1 0 83600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4258
timestamp 1757982896
transform 1 0 85100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4259
timestamp 1757982896
transform 1 0 86600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4260
timestamp 1757982896
transform 1 0 88100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4261
timestamp 1757982896
transform 1 0 89600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4262
timestamp 1757982896
transform 1 0 91100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4263
timestamp 1757982896
transform 1 0 92600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4264
timestamp 1757982896
transform 1 0 94100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4265
timestamp 1757982896
transform 1 0 95600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4266
timestamp 1757982896
transform 1 0 97100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4267
timestamp 1757982896
transform 1 0 98600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4268
timestamp 1757982896
transform 1 0 100100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4269
timestamp 1757982896
transform 1 0 101600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4270
timestamp 1757982896
transform 1 0 103100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4271
timestamp 1757982896
transform 1 0 104600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4272
timestamp 1757982896
transform 1 0 106100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4273
timestamp 1757982896
transform 1 0 107600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4274
timestamp 1757982896
transform 1 0 109100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4275
timestamp 1757982896
transform 1 0 110600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4276
timestamp 1757982896
transform 1 0 112100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4277
timestamp 1757982896
transform 1 0 113600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4278
timestamp 1757982896
transform 1 0 115100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4279
timestamp 1757982896
transform 1 0 116600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4280
timestamp 1757982896
transform 1 0 118100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4281
timestamp 1757982896
transform 1 0 119600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4282
timestamp 1757982896
transform 1 0 121100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4283
timestamp 1757982896
transform 1 0 122600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4284
timestamp 1757982896
transform 1 0 124100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4285
timestamp 1757982896
transform 1 0 125600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4286
timestamp 1757982896
transform 1 0 127100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4287
timestamp 1757982896
transform 1 0 128600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4288
timestamp 1757982896
transform 1 0 130100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4289
timestamp 1757982896
transform 1 0 131600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4290
timestamp 1757982896
transform 1 0 133100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4291
timestamp 1757982896
transform 1 0 134600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4292
timestamp 1757982896
transform 1 0 136100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4293
timestamp 1757982896
transform 1 0 137600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4294
timestamp 1757982896
transform 1 0 139100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4295
timestamp 1757982896
transform 1 0 140600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4296
timestamp 1757982896
transform 1 0 142100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4297
timestamp 1757982896
transform 1 0 143600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4298
timestamp 1757982896
transform 1 0 145100 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4299
timestamp 1757982896
transform 1 0 146600 0 1 -61650
box 1820 -1430 3480 230
use pixel  pixel_4300
timestamp 1757982896
transform 1 0 -1900 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4301
timestamp 1757982896
transform 1 0 -400 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4302
timestamp 1757982896
transform 1 0 1100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4303
timestamp 1757982896
transform 1 0 2600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4304
timestamp 1757982896
transform 1 0 4100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4305
timestamp 1757982896
transform 1 0 5600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4306
timestamp 1757982896
transform 1 0 7100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4307
timestamp 1757982896
transform 1 0 8600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4308
timestamp 1757982896
transform 1 0 10100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4309
timestamp 1757982896
transform 1 0 11600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4310
timestamp 1757982896
transform 1 0 13100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4311
timestamp 1757982896
transform 1 0 14600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4312
timestamp 1757982896
transform 1 0 16100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4313
timestamp 1757982896
transform 1 0 17600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4314
timestamp 1757982896
transform 1 0 19100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4315
timestamp 1757982896
transform 1 0 20600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4316
timestamp 1757982896
transform 1 0 22100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4317
timestamp 1757982896
transform 1 0 23600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4318
timestamp 1757982896
transform 1 0 25100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4319
timestamp 1757982896
transform 1 0 26600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4320
timestamp 1757982896
transform 1 0 28100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4321
timestamp 1757982896
transform 1 0 29600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4322
timestamp 1757982896
transform 1 0 31100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4323
timestamp 1757982896
transform 1 0 32600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4324
timestamp 1757982896
transform 1 0 34100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4325
timestamp 1757982896
transform 1 0 35600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4326
timestamp 1757982896
transform 1 0 37100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4327
timestamp 1757982896
transform 1 0 38600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4328
timestamp 1757982896
transform 1 0 40100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4329
timestamp 1757982896
transform 1 0 41600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4330
timestamp 1757982896
transform 1 0 43100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4331
timestamp 1757982896
transform 1 0 44600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4332
timestamp 1757982896
transform 1 0 46100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4333
timestamp 1757982896
transform 1 0 47600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4334
timestamp 1757982896
transform 1 0 49100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4335
timestamp 1757982896
transform 1 0 50600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4336
timestamp 1757982896
transform 1 0 52100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4337
timestamp 1757982896
transform 1 0 53600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4338
timestamp 1757982896
transform 1 0 55100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4339
timestamp 1757982896
transform 1 0 56600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4340
timestamp 1757982896
transform 1 0 58100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4341
timestamp 1757982896
transform 1 0 59600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4342
timestamp 1757982896
transform 1 0 61100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4343
timestamp 1757982896
transform 1 0 62600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4344
timestamp 1757982896
transform 1 0 64100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4345
timestamp 1757982896
transform 1 0 65600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4346
timestamp 1757982896
transform 1 0 67100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4347
timestamp 1757982896
transform 1 0 68600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4348
timestamp 1757982896
transform 1 0 70100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4349
timestamp 1757982896
transform 1 0 71600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4350
timestamp 1757982896
transform 1 0 73100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4351
timestamp 1757982896
transform 1 0 74600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4352
timestamp 1757982896
transform 1 0 76100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4353
timestamp 1757982896
transform 1 0 77600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4354
timestamp 1757982896
transform 1 0 79100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4355
timestamp 1757982896
transform 1 0 80600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4356
timestamp 1757982896
transform 1 0 82100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4357
timestamp 1757982896
transform 1 0 83600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4358
timestamp 1757982896
transform 1 0 85100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4359
timestamp 1757982896
transform 1 0 86600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4360
timestamp 1757982896
transform 1 0 88100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4361
timestamp 1757982896
transform 1 0 89600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4362
timestamp 1757982896
transform 1 0 91100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4363
timestamp 1757982896
transform 1 0 92600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4364
timestamp 1757982896
transform 1 0 94100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4365
timestamp 1757982896
transform 1 0 95600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4366
timestamp 1757982896
transform 1 0 97100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4367
timestamp 1757982896
transform 1 0 98600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4368
timestamp 1757982896
transform 1 0 100100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4369
timestamp 1757982896
transform 1 0 101600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4370
timestamp 1757982896
transform 1 0 103100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4371
timestamp 1757982896
transform 1 0 104600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4372
timestamp 1757982896
transform 1 0 106100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4373
timestamp 1757982896
transform 1 0 107600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4374
timestamp 1757982896
transform 1 0 109100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4375
timestamp 1757982896
transform 1 0 110600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4376
timestamp 1757982896
transform 1 0 112100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4377
timestamp 1757982896
transform 1 0 113600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4378
timestamp 1757982896
transform 1 0 115100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4379
timestamp 1757982896
transform 1 0 116600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4380
timestamp 1757982896
transform 1 0 118100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4381
timestamp 1757982896
transform 1 0 119600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4382
timestamp 1757982896
transform 1 0 121100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4383
timestamp 1757982896
transform 1 0 122600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4384
timestamp 1757982896
transform 1 0 124100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4385
timestamp 1757982896
transform 1 0 125600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4386
timestamp 1757982896
transform 1 0 127100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4387
timestamp 1757982896
transform 1 0 128600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4388
timestamp 1757982896
transform 1 0 130100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4389
timestamp 1757982896
transform 1 0 131600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4390
timestamp 1757982896
transform 1 0 133100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4391
timestamp 1757982896
transform 1 0 134600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4392
timestamp 1757982896
transform 1 0 136100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4393
timestamp 1757982896
transform 1 0 137600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4394
timestamp 1757982896
transform 1 0 139100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4395
timestamp 1757982896
transform 1 0 140600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4396
timestamp 1757982896
transform 1 0 142100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4397
timestamp 1757982896
transform 1 0 143600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4398
timestamp 1757982896
transform 1 0 145100 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4399
timestamp 1757982896
transform 1 0 146600 0 1 -63150
box 1820 -1430 3480 230
use pixel  pixel_4400
timestamp 1757982896
transform 1 0 -1900 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4401
timestamp 1757982896
transform 1 0 -400 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4402
timestamp 1757982896
transform 1 0 1100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4403
timestamp 1757982896
transform 1 0 2600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4404
timestamp 1757982896
transform 1 0 4100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4405
timestamp 1757982896
transform 1 0 5600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4406
timestamp 1757982896
transform 1 0 7100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4407
timestamp 1757982896
transform 1 0 8600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4408
timestamp 1757982896
transform 1 0 10100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4409
timestamp 1757982896
transform 1 0 11600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4410
timestamp 1757982896
transform 1 0 13100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4411
timestamp 1757982896
transform 1 0 14600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4412
timestamp 1757982896
transform 1 0 16100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4413
timestamp 1757982896
transform 1 0 17600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4414
timestamp 1757982896
transform 1 0 19100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4415
timestamp 1757982896
transform 1 0 20600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4416
timestamp 1757982896
transform 1 0 22100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4417
timestamp 1757982896
transform 1 0 23600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4418
timestamp 1757982896
transform 1 0 25100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4419
timestamp 1757982896
transform 1 0 26600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4420
timestamp 1757982896
transform 1 0 28100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4421
timestamp 1757982896
transform 1 0 29600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4422
timestamp 1757982896
transform 1 0 31100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4423
timestamp 1757982896
transform 1 0 32600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4424
timestamp 1757982896
transform 1 0 34100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4425
timestamp 1757982896
transform 1 0 35600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4426
timestamp 1757982896
transform 1 0 37100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4427
timestamp 1757982896
transform 1 0 38600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4428
timestamp 1757982896
transform 1 0 40100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4429
timestamp 1757982896
transform 1 0 41600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4430
timestamp 1757982896
transform 1 0 43100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4431
timestamp 1757982896
transform 1 0 44600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4432
timestamp 1757982896
transform 1 0 46100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4433
timestamp 1757982896
transform 1 0 47600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4434
timestamp 1757982896
transform 1 0 49100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4435
timestamp 1757982896
transform 1 0 50600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4436
timestamp 1757982896
transform 1 0 52100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4437
timestamp 1757982896
transform 1 0 53600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4438
timestamp 1757982896
transform 1 0 55100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4439
timestamp 1757982896
transform 1 0 56600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4440
timestamp 1757982896
transform 1 0 58100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4441
timestamp 1757982896
transform 1 0 59600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4442
timestamp 1757982896
transform 1 0 61100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4443
timestamp 1757982896
transform 1 0 62600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4444
timestamp 1757982896
transform 1 0 64100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4445
timestamp 1757982896
transform 1 0 65600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4446
timestamp 1757982896
transform 1 0 67100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4447
timestamp 1757982896
transform 1 0 68600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4448
timestamp 1757982896
transform 1 0 70100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4449
timestamp 1757982896
transform 1 0 71600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4450
timestamp 1757982896
transform 1 0 73100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4451
timestamp 1757982896
transform 1 0 74600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4452
timestamp 1757982896
transform 1 0 76100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4453
timestamp 1757982896
transform 1 0 77600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4454
timestamp 1757982896
transform 1 0 79100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4455
timestamp 1757982896
transform 1 0 80600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4456
timestamp 1757982896
transform 1 0 82100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4457
timestamp 1757982896
transform 1 0 83600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4458
timestamp 1757982896
transform 1 0 85100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4459
timestamp 1757982896
transform 1 0 86600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4460
timestamp 1757982896
transform 1 0 88100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4461
timestamp 1757982896
transform 1 0 89600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4462
timestamp 1757982896
transform 1 0 91100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4463
timestamp 1757982896
transform 1 0 92600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4464
timestamp 1757982896
transform 1 0 94100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4465
timestamp 1757982896
transform 1 0 95600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4466
timestamp 1757982896
transform 1 0 97100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4467
timestamp 1757982896
transform 1 0 98600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4468
timestamp 1757982896
transform 1 0 100100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4469
timestamp 1757982896
transform 1 0 101600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4470
timestamp 1757982896
transform 1 0 103100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4471
timestamp 1757982896
transform 1 0 104600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4472
timestamp 1757982896
transform 1 0 106100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4473
timestamp 1757982896
transform 1 0 107600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4474
timestamp 1757982896
transform 1 0 109100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4475
timestamp 1757982896
transform 1 0 110600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4476
timestamp 1757982896
transform 1 0 112100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4477
timestamp 1757982896
transform 1 0 113600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4478
timestamp 1757982896
transform 1 0 115100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4479
timestamp 1757982896
transform 1 0 116600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4480
timestamp 1757982896
transform 1 0 118100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4481
timestamp 1757982896
transform 1 0 119600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4482
timestamp 1757982896
transform 1 0 121100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4483
timestamp 1757982896
transform 1 0 122600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4484
timestamp 1757982896
transform 1 0 124100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4485
timestamp 1757982896
transform 1 0 125600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4486
timestamp 1757982896
transform 1 0 127100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4487
timestamp 1757982896
transform 1 0 128600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4488
timestamp 1757982896
transform 1 0 130100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4489
timestamp 1757982896
transform 1 0 131600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4490
timestamp 1757982896
transform 1 0 133100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4491
timestamp 1757982896
transform 1 0 134600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4492
timestamp 1757982896
transform 1 0 136100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4493
timestamp 1757982896
transform 1 0 137600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4494
timestamp 1757982896
transform 1 0 139100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4495
timestamp 1757982896
transform 1 0 140600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4496
timestamp 1757982896
transform 1 0 142100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4497
timestamp 1757982896
transform 1 0 143600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4498
timestamp 1757982896
transform 1 0 145100 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4499
timestamp 1757982896
transform 1 0 146600 0 1 -64650
box 1820 -1430 3480 230
use pixel  pixel_4500
timestamp 1757982896
transform 1 0 -1900 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4501
timestamp 1757982896
transform 1 0 -400 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4502
timestamp 1757982896
transform 1 0 1100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4503
timestamp 1757982896
transform 1 0 2600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4504
timestamp 1757982896
transform 1 0 4100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4505
timestamp 1757982896
transform 1 0 5600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4506
timestamp 1757982896
transform 1 0 7100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4507
timestamp 1757982896
transform 1 0 8600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4508
timestamp 1757982896
transform 1 0 10100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4509
timestamp 1757982896
transform 1 0 11600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4510
timestamp 1757982896
transform 1 0 13100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4511
timestamp 1757982896
transform 1 0 14600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4512
timestamp 1757982896
transform 1 0 16100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4513
timestamp 1757982896
transform 1 0 17600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4514
timestamp 1757982896
transform 1 0 19100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4515
timestamp 1757982896
transform 1 0 20600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4516
timestamp 1757982896
transform 1 0 22100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4517
timestamp 1757982896
transform 1 0 23600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4518
timestamp 1757982896
transform 1 0 25100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4519
timestamp 1757982896
transform 1 0 26600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4520
timestamp 1757982896
transform 1 0 28100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4521
timestamp 1757982896
transform 1 0 29600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4522
timestamp 1757982896
transform 1 0 31100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4523
timestamp 1757982896
transform 1 0 32600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4524
timestamp 1757982896
transform 1 0 34100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4525
timestamp 1757982896
transform 1 0 35600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4526
timestamp 1757982896
transform 1 0 37100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4527
timestamp 1757982896
transform 1 0 38600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4528
timestamp 1757982896
transform 1 0 40100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4529
timestamp 1757982896
transform 1 0 41600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4530
timestamp 1757982896
transform 1 0 43100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4531
timestamp 1757982896
transform 1 0 44600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4532
timestamp 1757982896
transform 1 0 46100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4533
timestamp 1757982896
transform 1 0 47600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4534
timestamp 1757982896
transform 1 0 49100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4535
timestamp 1757982896
transform 1 0 50600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4536
timestamp 1757982896
transform 1 0 52100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4537
timestamp 1757982896
transform 1 0 53600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4538
timestamp 1757982896
transform 1 0 55100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4539
timestamp 1757982896
transform 1 0 56600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4540
timestamp 1757982896
transform 1 0 58100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4541
timestamp 1757982896
transform 1 0 59600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4542
timestamp 1757982896
transform 1 0 61100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4543
timestamp 1757982896
transform 1 0 62600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4544
timestamp 1757982896
transform 1 0 64100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4545
timestamp 1757982896
transform 1 0 65600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4546
timestamp 1757982896
transform 1 0 67100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4547
timestamp 1757982896
transform 1 0 68600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4548
timestamp 1757982896
transform 1 0 70100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4549
timestamp 1757982896
transform 1 0 71600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4550
timestamp 1757982896
transform 1 0 73100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4551
timestamp 1757982896
transform 1 0 74600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4552
timestamp 1757982896
transform 1 0 76100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4553
timestamp 1757982896
transform 1 0 77600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4554
timestamp 1757982896
transform 1 0 79100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4555
timestamp 1757982896
transform 1 0 80600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4556
timestamp 1757982896
transform 1 0 82100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4557
timestamp 1757982896
transform 1 0 83600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4558
timestamp 1757982896
transform 1 0 85100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4559
timestamp 1757982896
transform 1 0 86600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4560
timestamp 1757982896
transform 1 0 88100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4561
timestamp 1757982896
transform 1 0 89600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4562
timestamp 1757982896
transform 1 0 91100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4563
timestamp 1757982896
transform 1 0 92600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4564
timestamp 1757982896
transform 1 0 94100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4565
timestamp 1757982896
transform 1 0 95600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4566
timestamp 1757982896
transform 1 0 97100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4567
timestamp 1757982896
transform 1 0 98600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4568
timestamp 1757982896
transform 1 0 100100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4569
timestamp 1757982896
transform 1 0 101600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4570
timestamp 1757982896
transform 1 0 103100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4571
timestamp 1757982896
transform 1 0 104600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4572
timestamp 1757982896
transform 1 0 106100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4573
timestamp 1757982896
transform 1 0 107600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4574
timestamp 1757982896
transform 1 0 109100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4575
timestamp 1757982896
transform 1 0 110600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4576
timestamp 1757982896
transform 1 0 112100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4577
timestamp 1757982896
transform 1 0 113600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4578
timestamp 1757982896
transform 1 0 115100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4579
timestamp 1757982896
transform 1 0 116600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4580
timestamp 1757982896
transform 1 0 118100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4581
timestamp 1757982896
transform 1 0 119600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4582
timestamp 1757982896
transform 1 0 121100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4583
timestamp 1757982896
transform 1 0 122600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4584
timestamp 1757982896
transform 1 0 124100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4585
timestamp 1757982896
transform 1 0 125600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4586
timestamp 1757982896
transform 1 0 127100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4587
timestamp 1757982896
transform 1 0 128600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4588
timestamp 1757982896
transform 1 0 130100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4589
timestamp 1757982896
transform 1 0 131600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4590
timestamp 1757982896
transform 1 0 133100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4591
timestamp 1757982896
transform 1 0 134600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4592
timestamp 1757982896
transform 1 0 136100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4593
timestamp 1757982896
transform 1 0 137600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4594
timestamp 1757982896
transform 1 0 139100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4595
timestamp 1757982896
transform 1 0 140600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4596
timestamp 1757982896
transform 1 0 142100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4597
timestamp 1757982896
transform 1 0 143600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4598
timestamp 1757982896
transform 1 0 145100 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4599
timestamp 1757982896
transform 1 0 146600 0 1 -66150
box 1820 -1430 3480 230
use pixel  pixel_4600
timestamp 1757982896
transform 1 0 -1900 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4601
timestamp 1757982896
transform 1 0 -400 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4602
timestamp 1757982896
transform 1 0 1100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4603
timestamp 1757982896
transform 1 0 2600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4604
timestamp 1757982896
transform 1 0 4100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4605
timestamp 1757982896
transform 1 0 5600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4606
timestamp 1757982896
transform 1 0 7100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4607
timestamp 1757982896
transform 1 0 8600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4608
timestamp 1757982896
transform 1 0 10100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4609
timestamp 1757982896
transform 1 0 11600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4610
timestamp 1757982896
transform 1 0 13100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4611
timestamp 1757982896
transform 1 0 14600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4612
timestamp 1757982896
transform 1 0 16100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4613
timestamp 1757982896
transform 1 0 17600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4614
timestamp 1757982896
transform 1 0 19100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4615
timestamp 1757982896
transform 1 0 20600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4616
timestamp 1757982896
transform 1 0 22100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4617
timestamp 1757982896
transform 1 0 23600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4618
timestamp 1757982896
transform 1 0 25100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4619
timestamp 1757982896
transform 1 0 26600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4620
timestamp 1757982896
transform 1 0 28100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4621
timestamp 1757982896
transform 1 0 29600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4622
timestamp 1757982896
transform 1 0 31100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4623
timestamp 1757982896
transform 1 0 32600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4624
timestamp 1757982896
transform 1 0 34100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4625
timestamp 1757982896
transform 1 0 35600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4626
timestamp 1757982896
transform 1 0 37100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4627
timestamp 1757982896
transform 1 0 38600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4628
timestamp 1757982896
transform 1 0 40100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4629
timestamp 1757982896
transform 1 0 41600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4630
timestamp 1757982896
transform 1 0 43100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4631
timestamp 1757982896
transform 1 0 44600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4632
timestamp 1757982896
transform 1 0 46100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4633
timestamp 1757982896
transform 1 0 47600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4634
timestamp 1757982896
transform 1 0 49100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4635
timestamp 1757982896
transform 1 0 50600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4636
timestamp 1757982896
transform 1 0 52100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4637
timestamp 1757982896
transform 1 0 53600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4638
timestamp 1757982896
transform 1 0 55100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4639
timestamp 1757982896
transform 1 0 56600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4640
timestamp 1757982896
transform 1 0 58100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4641
timestamp 1757982896
transform 1 0 59600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4642
timestamp 1757982896
transform 1 0 61100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4643
timestamp 1757982896
transform 1 0 62600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4644
timestamp 1757982896
transform 1 0 64100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4645
timestamp 1757982896
transform 1 0 65600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4646
timestamp 1757982896
transform 1 0 67100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4647
timestamp 1757982896
transform 1 0 68600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4648
timestamp 1757982896
transform 1 0 70100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4649
timestamp 1757982896
transform 1 0 71600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4650
timestamp 1757982896
transform 1 0 73100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4651
timestamp 1757982896
transform 1 0 74600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4652
timestamp 1757982896
transform 1 0 76100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4653
timestamp 1757982896
transform 1 0 77600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4654
timestamp 1757982896
transform 1 0 79100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4655
timestamp 1757982896
transform 1 0 80600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4656
timestamp 1757982896
transform 1 0 82100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4657
timestamp 1757982896
transform 1 0 83600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4658
timestamp 1757982896
transform 1 0 85100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4659
timestamp 1757982896
transform 1 0 86600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4660
timestamp 1757982896
transform 1 0 88100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4661
timestamp 1757982896
transform 1 0 89600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4662
timestamp 1757982896
transform 1 0 91100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4663
timestamp 1757982896
transform 1 0 92600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4664
timestamp 1757982896
transform 1 0 94100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4665
timestamp 1757982896
transform 1 0 95600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4666
timestamp 1757982896
transform 1 0 97100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4667
timestamp 1757982896
transform 1 0 98600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4668
timestamp 1757982896
transform 1 0 100100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4669
timestamp 1757982896
transform 1 0 101600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4670
timestamp 1757982896
transform 1 0 103100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4671
timestamp 1757982896
transform 1 0 104600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4672
timestamp 1757982896
transform 1 0 106100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4673
timestamp 1757982896
transform 1 0 107600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4674
timestamp 1757982896
transform 1 0 109100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4675
timestamp 1757982896
transform 1 0 110600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4676
timestamp 1757982896
transform 1 0 112100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4677
timestamp 1757982896
transform 1 0 113600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4678
timestamp 1757982896
transform 1 0 115100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4679
timestamp 1757982896
transform 1 0 116600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4680
timestamp 1757982896
transform 1 0 118100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4681
timestamp 1757982896
transform 1 0 119600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4682
timestamp 1757982896
transform 1 0 121100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4683
timestamp 1757982896
transform 1 0 122600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4684
timestamp 1757982896
transform 1 0 124100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4685
timestamp 1757982896
transform 1 0 125600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4686
timestamp 1757982896
transform 1 0 127100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4687
timestamp 1757982896
transform 1 0 128600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4688
timestamp 1757982896
transform 1 0 130100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4689
timestamp 1757982896
transform 1 0 131600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4690
timestamp 1757982896
transform 1 0 133100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4691
timestamp 1757982896
transform 1 0 134600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4692
timestamp 1757982896
transform 1 0 136100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4693
timestamp 1757982896
transform 1 0 137600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4694
timestamp 1757982896
transform 1 0 139100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4695
timestamp 1757982896
transform 1 0 140600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4696
timestamp 1757982896
transform 1 0 142100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4697
timestamp 1757982896
transform 1 0 143600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4698
timestamp 1757982896
transform 1 0 145100 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4699
timestamp 1757982896
transform 1 0 146600 0 1 -67650
box 1820 -1430 3480 230
use pixel  pixel_4700
timestamp 1757982896
transform 1 0 -1900 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4701
timestamp 1757982896
transform 1 0 -400 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4702
timestamp 1757982896
transform 1 0 1100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4703
timestamp 1757982896
transform 1 0 2600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4704
timestamp 1757982896
transform 1 0 4100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4705
timestamp 1757982896
transform 1 0 5600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4706
timestamp 1757982896
transform 1 0 7100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4707
timestamp 1757982896
transform 1 0 8600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4708
timestamp 1757982896
transform 1 0 10100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4709
timestamp 1757982896
transform 1 0 11600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4710
timestamp 1757982896
transform 1 0 13100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4711
timestamp 1757982896
transform 1 0 14600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4712
timestamp 1757982896
transform 1 0 16100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4713
timestamp 1757982896
transform 1 0 17600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4714
timestamp 1757982896
transform 1 0 19100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4715
timestamp 1757982896
transform 1 0 20600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4716
timestamp 1757982896
transform 1 0 22100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4717
timestamp 1757982896
transform 1 0 23600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4718
timestamp 1757982896
transform 1 0 25100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4719
timestamp 1757982896
transform 1 0 26600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4720
timestamp 1757982896
transform 1 0 28100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4721
timestamp 1757982896
transform 1 0 29600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4722
timestamp 1757982896
transform 1 0 31100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4723
timestamp 1757982896
transform 1 0 32600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4724
timestamp 1757982896
transform 1 0 34100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4725
timestamp 1757982896
transform 1 0 35600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4726
timestamp 1757982896
transform 1 0 37100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4727
timestamp 1757982896
transform 1 0 38600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4728
timestamp 1757982896
transform 1 0 40100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4729
timestamp 1757982896
transform 1 0 41600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4730
timestamp 1757982896
transform 1 0 43100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4731
timestamp 1757982896
transform 1 0 44600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4732
timestamp 1757982896
transform 1 0 46100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4733
timestamp 1757982896
transform 1 0 47600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4734
timestamp 1757982896
transform 1 0 49100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4735
timestamp 1757982896
transform 1 0 50600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4736
timestamp 1757982896
transform 1 0 52100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4737
timestamp 1757982896
transform 1 0 53600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4738
timestamp 1757982896
transform 1 0 55100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4739
timestamp 1757982896
transform 1 0 56600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4740
timestamp 1757982896
transform 1 0 58100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4741
timestamp 1757982896
transform 1 0 59600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4742
timestamp 1757982896
transform 1 0 61100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4743
timestamp 1757982896
transform 1 0 62600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4744
timestamp 1757982896
transform 1 0 64100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4745
timestamp 1757982896
transform 1 0 65600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4746
timestamp 1757982896
transform 1 0 67100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4747
timestamp 1757982896
transform 1 0 68600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4748
timestamp 1757982896
transform 1 0 70100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4749
timestamp 1757982896
transform 1 0 71600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4750
timestamp 1757982896
transform 1 0 73100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4751
timestamp 1757982896
transform 1 0 74600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4752
timestamp 1757982896
transform 1 0 76100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4753
timestamp 1757982896
transform 1 0 77600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4754
timestamp 1757982896
transform 1 0 79100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4755
timestamp 1757982896
transform 1 0 80600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4756
timestamp 1757982896
transform 1 0 82100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4757
timestamp 1757982896
transform 1 0 83600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4758
timestamp 1757982896
transform 1 0 85100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4759
timestamp 1757982896
transform 1 0 86600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4760
timestamp 1757982896
transform 1 0 88100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4761
timestamp 1757982896
transform 1 0 89600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4762
timestamp 1757982896
transform 1 0 91100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4763
timestamp 1757982896
transform 1 0 92600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4764
timestamp 1757982896
transform 1 0 94100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4765
timestamp 1757982896
transform 1 0 95600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4766
timestamp 1757982896
transform 1 0 97100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4767
timestamp 1757982896
transform 1 0 98600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4768
timestamp 1757982896
transform 1 0 100100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4769
timestamp 1757982896
transform 1 0 101600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4770
timestamp 1757982896
transform 1 0 103100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4771
timestamp 1757982896
transform 1 0 104600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4772
timestamp 1757982896
transform 1 0 106100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4773
timestamp 1757982896
transform 1 0 107600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4774
timestamp 1757982896
transform 1 0 109100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4775
timestamp 1757982896
transform 1 0 110600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4776
timestamp 1757982896
transform 1 0 112100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4777
timestamp 1757982896
transform 1 0 113600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4778
timestamp 1757982896
transform 1 0 115100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4779
timestamp 1757982896
transform 1 0 116600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4780
timestamp 1757982896
transform 1 0 118100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4781
timestamp 1757982896
transform 1 0 119600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4782
timestamp 1757982896
transform 1 0 121100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4783
timestamp 1757982896
transform 1 0 122600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4784
timestamp 1757982896
transform 1 0 124100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4785
timestamp 1757982896
transform 1 0 125600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4786
timestamp 1757982896
transform 1 0 127100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4787
timestamp 1757982896
transform 1 0 128600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4788
timestamp 1757982896
transform 1 0 130100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4789
timestamp 1757982896
transform 1 0 131600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4790
timestamp 1757982896
transform 1 0 133100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4791
timestamp 1757982896
transform 1 0 134600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4792
timestamp 1757982896
transform 1 0 136100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4793
timestamp 1757982896
transform 1 0 137600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4794
timestamp 1757982896
transform 1 0 139100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4795
timestamp 1757982896
transform 1 0 140600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4796
timestamp 1757982896
transform 1 0 142100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4797
timestamp 1757982896
transform 1 0 143600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4798
timestamp 1757982896
transform 1 0 145100 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4799
timestamp 1757982896
transform 1 0 146600 0 1 -69150
box 1820 -1430 3480 230
use pixel  pixel_4800
timestamp 1757982896
transform 1 0 -1900 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4801
timestamp 1757982896
transform 1 0 -400 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4802
timestamp 1757982896
transform 1 0 1100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4803
timestamp 1757982896
transform 1 0 2600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4804
timestamp 1757982896
transform 1 0 4100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4805
timestamp 1757982896
transform 1 0 5600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4806
timestamp 1757982896
transform 1 0 7100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4807
timestamp 1757982896
transform 1 0 8600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4808
timestamp 1757982896
transform 1 0 10100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4809
timestamp 1757982896
transform 1 0 11600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4810
timestamp 1757982896
transform 1 0 13100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4811
timestamp 1757982896
transform 1 0 14600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4812
timestamp 1757982896
transform 1 0 16100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4813
timestamp 1757982896
transform 1 0 17600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4814
timestamp 1757982896
transform 1 0 19100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4815
timestamp 1757982896
transform 1 0 20600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4816
timestamp 1757982896
transform 1 0 22100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4817
timestamp 1757982896
transform 1 0 23600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4818
timestamp 1757982896
transform 1 0 25100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4819
timestamp 1757982896
transform 1 0 26600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4820
timestamp 1757982896
transform 1 0 28100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4821
timestamp 1757982896
transform 1 0 29600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4822
timestamp 1757982896
transform 1 0 31100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4823
timestamp 1757982896
transform 1 0 32600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4824
timestamp 1757982896
transform 1 0 34100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4825
timestamp 1757982896
transform 1 0 35600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4826
timestamp 1757982896
transform 1 0 37100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4827
timestamp 1757982896
transform 1 0 38600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4828
timestamp 1757982896
transform 1 0 40100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4829
timestamp 1757982896
transform 1 0 41600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4830
timestamp 1757982896
transform 1 0 43100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4831
timestamp 1757982896
transform 1 0 44600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4832
timestamp 1757982896
transform 1 0 46100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4833
timestamp 1757982896
transform 1 0 47600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4834
timestamp 1757982896
transform 1 0 49100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4835
timestamp 1757982896
transform 1 0 50600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4836
timestamp 1757982896
transform 1 0 52100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4837
timestamp 1757982896
transform 1 0 53600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4838
timestamp 1757982896
transform 1 0 55100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4839
timestamp 1757982896
transform 1 0 56600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4840
timestamp 1757982896
transform 1 0 58100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4841
timestamp 1757982896
transform 1 0 59600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4842
timestamp 1757982896
transform 1 0 61100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4843
timestamp 1757982896
transform 1 0 62600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4844
timestamp 1757982896
transform 1 0 64100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4845
timestamp 1757982896
transform 1 0 65600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4846
timestamp 1757982896
transform 1 0 67100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4847
timestamp 1757982896
transform 1 0 68600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4848
timestamp 1757982896
transform 1 0 70100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4849
timestamp 1757982896
transform 1 0 71600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4850
timestamp 1757982896
transform 1 0 73100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4851
timestamp 1757982896
transform 1 0 74600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4852
timestamp 1757982896
transform 1 0 76100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4853
timestamp 1757982896
transform 1 0 77600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4854
timestamp 1757982896
transform 1 0 79100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4855
timestamp 1757982896
transform 1 0 80600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4856
timestamp 1757982896
transform 1 0 82100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4857
timestamp 1757982896
transform 1 0 83600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4858
timestamp 1757982896
transform 1 0 85100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4859
timestamp 1757982896
transform 1 0 86600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4860
timestamp 1757982896
transform 1 0 88100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4861
timestamp 1757982896
transform 1 0 89600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4862
timestamp 1757982896
transform 1 0 91100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4863
timestamp 1757982896
transform 1 0 92600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4864
timestamp 1757982896
transform 1 0 94100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4865
timestamp 1757982896
transform 1 0 95600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4866
timestamp 1757982896
transform 1 0 97100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4867
timestamp 1757982896
transform 1 0 98600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4868
timestamp 1757982896
transform 1 0 100100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4869
timestamp 1757982896
transform 1 0 101600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4870
timestamp 1757982896
transform 1 0 103100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4871
timestamp 1757982896
transform 1 0 104600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4872
timestamp 1757982896
transform 1 0 106100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4873
timestamp 1757982896
transform 1 0 107600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4874
timestamp 1757982896
transform 1 0 109100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4875
timestamp 1757982896
transform 1 0 110600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4876
timestamp 1757982896
transform 1 0 112100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4877
timestamp 1757982896
transform 1 0 113600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4878
timestamp 1757982896
transform 1 0 115100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4879
timestamp 1757982896
transform 1 0 116600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4880
timestamp 1757982896
transform 1 0 118100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4881
timestamp 1757982896
transform 1 0 119600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4882
timestamp 1757982896
transform 1 0 121100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4883
timestamp 1757982896
transform 1 0 122600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4884
timestamp 1757982896
transform 1 0 124100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4885
timestamp 1757982896
transform 1 0 125600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4886
timestamp 1757982896
transform 1 0 127100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4887
timestamp 1757982896
transform 1 0 128600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4888
timestamp 1757982896
transform 1 0 130100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4889
timestamp 1757982896
transform 1 0 131600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4890
timestamp 1757982896
transform 1 0 133100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4891
timestamp 1757982896
transform 1 0 134600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4892
timestamp 1757982896
transform 1 0 136100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4893
timestamp 1757982896
transform 1 0 137600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4894
timestamp 1757982896
transform 1 0 139100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4895
timestamp 1757982896
transform 1 0 140600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4896
timestamp 1757982896
transform 1 0 142100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4897
timestamp 1757982896
transform 1 0 143600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4898
timestamp 1757982896
transform 1 0 145100 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4899
timestamp 1757982896
transform 1 0 146600 0 1 -70650
box 1820 -1430 3480 230
use pixel  pixel_4900
timestamp 1757982896
transform 1 0 -1900 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4901
timestamp 1757982896
transform 1 0 -400 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4902
timestamp 1757982896
transform 1 0 1100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4903
timestamp 1757982896
transform 1 0 2600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4904
timestamp 1757982896
transform 1 0 4100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4905
timestamp 1757982896
transform 1 0 5600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4906
timestamp 1757982896
transform 1 0 7100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4907
timestamp 1757982896
transform 1 0 8600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4908
timestamp 1757982896
transform 1 0 10100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4909
timestamp 1757982896
transform 1 0 11600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4910
timestamp 1757982896
transform 1 0 13100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4911
timestamp 1757982896
transform 1 0 14600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4912
timestamp 1757982896
transform 1 0 16100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4913
timestamp 1757982896
transform 1 0 17600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4914
timestamp 1757982896
transform 1 0 19100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4915
timestamp 1757982896
transform 1 0 20600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4916
timestamp 1757982896
transform 1 0 22100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4917
timestamp 1757982896
transform 1 0 23600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4918
timestamp 1757982896
transform 1 0 25100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4919
timestamp 1757982896
transform 1 0 26600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4920
timestamp 1757982896
transform 1 0 28100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4921
timestamp 1757982896
transform 1 0 29600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4922
timestamp 1757982896
transform 1 0 31100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4923
timestamp 1757982896
transform 1 0 32600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4924
timestamp 1757982896
transform 1 0 34100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4925
timestamp 1757982896
transform 1 0 35600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4926
timestamp 1757982896
transform 1 0 37100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4927
timestamp 1757982896
transform 1 0 38600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4928
timestamp 1757982896
transform 1 0 40100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4929
timestamp 1757982896
transform 1 0 41600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4930
timestamp 1757982896
transform 1 0 43100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4931
timestamp 1757982896
transform 1 0 44600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4932
timestamp 1757982896
transform 1 0 46100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4933
timestamp 1757982896
transform 1 0 47600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4934
timestamp 1757982896
transform 1 0 49100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4935
timestamp 1757982896
transform 1 0 50600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4936
timestamp 1757982896
transform 1 0 52100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4937
timestamp 1757982896
transform 1 0 53600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4938
timestamp 1757982896
transform 1 0 55100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4939
timestamp 1757982896
transform 1 0 56600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4940
timestamp 1757982896
transform 1 0 58100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4941
timestamp 1757982896
transform 1 0 59600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4942
timestamp 1757982896
transform 1 0 61100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4943
timestamp 1757982896
transform 1 0 62600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4944
timestamp 1757982896
transform 1 0 64100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4945
timestamp 1757982896
transform 1 0 65600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4946
timestamp 1757982896
transform 1 0 67100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4947
timestamp 1757982896
transform 1 0 68600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4948
timestamp 1757982896
transform 1 0 70100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4949
timestamp 1757982896
transform 1 0 71600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4950
timestamp 1757982896
transform 1 0 73100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4951
timestamp 1757982896
transform 1 0 74600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4952
timestamp 1757982896
transform 1 0 76100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4953
timestamp 1757982896
transform 1 0 77600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4954
timestamp 1757982896
transform 1 0 79100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4955
timestamp 1757982896
transform 1 0 80600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4956
timestamp 1757982896
transform 1 0 82100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4957
timestamp 1757982896
transform 1 0 83600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4958
timestamp 1757982896
transform 1 0 85100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4959
timestamp 1757982896
transform 1 0 86600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4960
timestamp 1757982896
transform 1 0 88100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4961
timestamp 1757982896
transform 1 0 89600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4962
timestamp 1757982896
transform 1 0 91100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4963
timestamp 1757982896
transform 1 0 92600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4964
timestamp 1757982896
transform 1 0 94100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4965
timestamp 1757982896
transform 1 0 95600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4966
timestamp 1757982896
transform 1 0 97100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4967
timestamp 1757982896
transform 1 0 98600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4968
timestamp 1757982896
transform 1 0 100100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4969
timestamp 1757982896
transform 1 0 101600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4970
timestamp 1757982896
transform 1 0 103100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4971
timestamp 1757982896
transform 1 0 104600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4972
timestamp 1757982896
transform 1 0 106100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4973
timestamp 1757982896
transform 1 0 107600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4974
timestamp 1757982896
transform 1 0 109100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4975
timestamp 1757982896
transform 1 0 110600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4976
timestamp 1757982896
transform 1 0 112100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4977
timestamp 1757982896
transform 1 0 113600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4978
timestamp 1757982896
transform 1 0 115100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4979
timestamp 1757982896
transform 1 0 116600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4980
timestamp 1757982896
transform 1 0 118100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4981
timestamp 1757982896
transform 1 0 119600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4982
timestamp 1757982896
transform 1 0 121100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4983
timestamp 1757982896
transform 1 0 122600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4984
timestamp 1757982896
transform 1 0 124100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4985
timestamp 1757982896
transform 1 0 125600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4986
timestamp 1757982896
transform 1 0 127100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4987
timestamp 1757982896
transform 1 0 128600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4988
timestamp 1757982896
transform 1 0 130100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4989
timestamp 1757982896
transform 1 0 131600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4990
timestamp 1757982896
transform 1 0 133100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4991
timestamp 1757982896
transform 1 0 134600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4992
timestamp 1757982896
transform 1 0 136100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4993
timestamp 1757982896
transform 1 0 137600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4994
timestamp 1757982896
transform 1 0 139100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4995
timestamp 1757982896
transform 1 0 140600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4996
timestamp 1757982896
transform 1 0 142100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4997
timestamp 1757982896
transform 1 0 143600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4998
timestamp 1757982896
transform 1 0 145100 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_4999
timestamp 1757982896
transform 1 0 146600 0 1 -72150
box 1820 -1430 3480 230
use pixel  pixel_5000
timestamp 1757982896
transform 1 0 -1900 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5001
timestamp 1757982896
transform 1 0 -400 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5002
timestamp 1757982896
transform 1 0 1100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5003
timestamp 1757982896
transform 1 0 2600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5004
timestamp 1757982896
transform 1 0 4100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5005
timestamp 1757982896
transform 1 0 5600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5006
timestamp 1757982896
transform 1 0 7100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5007
timestamp 1757982896
transform 1 0 8600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5008
timestamp 1757982896
transform 1 0 10100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5009
timestamp 1757982896
transform 1 0 11600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5010
timestamp 1757982896
transform 1 0 13100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5011
timestamp 1757982896
transform 1 0 14600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5012
timestamp 1757982896
transform 1 0 16100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5013
timestamp 1757982896
transform 1 0 17600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5014
timestamp 1757982896
transform 1 0 19100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5015
timestamp 1757982896
transform 1 0 20600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5016
timestamp 1757982896
transform 1 0 22100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5017
timestamp 1757982896
transform 1 0 23600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5018
timestamp 1757982896
transform 1 0 25100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5019
timestamp 1757982896
transform 1 0 26600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5020
timestamp 1757982896
transform 1 0 28100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5021
timestamp 1757982896
transform 1 0 29600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5022
timestamp 1757982896
transform 1 0 31100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5023
timestamp 1757982896
transform 1 0 32600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5024
timestamp 1757982896
transform 1 0 34100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5025
timestamp 1757982896
transform 1 0 35600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5026
timestamp 1757982896
transform 1 0 37100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5027
timestamp 1757982896
transform 1 0 38600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5028
timestamp 1757982896
transform 1 0 40100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5029
timestamp 1757982896
transform 1 0 41600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5030
timestamp 1757982896
transform 1 0 43100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5031
timestamp 1757982896
transform 1 0 44600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5032
timestamp 1757982896
transform 1 0 46100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5033
timestamp 1757982896
transform 1 0 47600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5034
timestamp 1757982896
transform 1 0 49100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5035
timestamp 1757982896
transform 1 0 50600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5036
timestamp 1757982896
transform 1 0 52100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5037
timestamp 1757982896
transform 1 0 53600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5038
timestamp 1757982896
transform 1 0 55100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5039
timestamp 1757982896
transform 1 0 56600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5040
timestamp 1757982896
transform 1 0 58100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5041
timestamp 1757982896
transform 1 0 59600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5042
timestamp 1757982896
transform 1 0 61100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5043
timestamp 1757982896
transform 1 0 62600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5044
timestamp 1757982896
transform 1 0 64100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5045
timestamp 1757982896
transform 1 0 65600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5046
timestamp 1757982896
transform 1 0 67100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5047
timestamp 1757982896
transform 1 0 68600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5048
timestamp 1757982896
transform 1 0 70100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5049
timestamp 1757982896
transform 1 0 71600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5050
timestamp 1757982896
transform 1 0 73100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5051
timestamp 1757982896
transform 1 0 74600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5052
timestamp 1757982896
transform 1 0 76100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5053
timestamp 1757982896
transform 1 0 77600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5054
timestamp 1757982896
transform 1 0 79100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5055
timestamp 1757982896
transform 1 0 80600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5056
timestamp 1757982896
transform 1 0 82100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5057
timestamp 1757982896
transform 1 0 83600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5058
timestamp 1757982896
transform 1 0 85100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5059
timestamp 1757982896
transform 1 0 86600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5060
timestamp 1757982896
transform 1 0 88100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5061
timestamp 1757982896
transform 1 0 89600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5062
timestamp 1757982896
transform 1 0 91100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5063
timestamp 1757982896
transform 1 0 92600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5064
timestamp 1757982896
transform 1 0 94100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5065
timestamp 1757982896
transform 1 0 95600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5066
timestamp 1757982896
transform 1 0 97100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5067
timestamp 1757982896
transform 1 0 98600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5068
timestamp 1757982896
transform 1 0 100100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5069
timestamp 1757982896
transform 1 0 101600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5070
timestamp 1757982896
transform 1 0 103100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5071
timestamp 1757982896
transform 1 0 104600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5072
timestamp 1757982896
transform 1 0 106100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5073
timestamp 1757982896
transform 1 0 107600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5074
timestamp 1757982896
transform 1 0 109100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5075
timestamp 1757982896
transform 1 0 110600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5076
timestamp 1757982896
transform 1 0 112100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5077
timestamp 1757982896
transform 1 0 113600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5078
timestamp 1757982896
transform 1 0 115100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5079
timestamp 1757982896
transform 1 0 116600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5080
timestamp 1757982896
transform 1 0 118100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5081
timestamp 1757982896
transform 1 0 119600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5082
timestamp 1757982896
transform 1 0 121100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5083
timestamp 1757982896
transform 1 0 122600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5084
timestamp 1757982896
transform 1 0 124100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5085
timestamp 1757982896
transform 1 0 125600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5086
timestamp 1757982896
transform 1 0 127100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5087
timestamp 1757982896
transform 1 0 128600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5088
timestamp 1757982896
transform 1 0 130100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5089
timestamp 1757982896
transform 1 0 131600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5090
timestamp 1757982896
transform 1 0 133100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5091
timestamp 1757982896
transform 1 0 134600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5092
timestamp 1757982896
transform 1 0 136100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5093
timestamp 1757982896
transform 1 0 137600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5094
timestamp 1757982896
transform 1 0 139100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5095
timestamp 1757982896
transform 1 0 140600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5096
timestamp 1757982896
transform 1 0 142100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5097
timestamp 1757982896
transform 1 0 143600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5098
timestamp 1757982896
transform 1 0 145100 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5099
timestamp 1757982896
transform 1 0 146600 0 1 -73650
box 1820 -1430 3480 230
use pixel  pixel_5100
timestamp 1757982896
transform 1 0 -1900 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5101
timestamp 1757982896
transform 1 0 -400 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5102
timestamp 1757982896
transform 1 0 1100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5103
timestamp 1757982896
transform 1 0 2600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5104
timestamp 1757982896
transform 1 0 4100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5105
timestamp 1757982896
transform 1 0 5600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5106
timestamp 1757982896
transform 1 0 7100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5107
timestamp 1757982896
transform 1 0 8600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5108
timestamp 1757982896
transform 1 0 10100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5109
timestamp 1757982896
transform 1 0 11600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5110
timestamp 1757982896
transform 1 0 13100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5111
timestamp 1757982896
transform 1 0 14600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5112
timestamp 1757982896
transform 1 0 16100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5113
timestamp 1757982896
transform 1 0 17600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5114
timestamp 1757982896
transform 1 0 19100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5115
timestamp 1757982896
transform 1 0 20600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5116
timestamp 1757982896
transform 1 0 22100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5117
timestamp 1757982896
transform 1 0 23600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5118
timestamp 1757982896
transform 1 0 25100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5119
timestamp 1757982896
transform 1 0 26600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5120
timestamp 1757982896
transform 1 0 28100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5121
timestamp 1757982896
transform 1 0 29600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5122
timestamp 1757982896
transform 1 0 31100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5123
timestamp 1757982896
transform 1 0 32600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5124
timestamp 1757982896
transform 1 0 34100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5125
timestamp 1757982896
transform 1 0 35600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5126
timestamp 1757982896
transform 1 0 37100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5127
timestamp 1757982896
transform 1 0 38600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5128
timestamp 1757982896
transform 1 0 40100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5129
timestamp 1757982896
transform 1 0 41600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5130
timestamp 1757982896
transform 1 0 43100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5131
timestamp 1757982896
transform 1 0 44600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5132
timestamp 1757982896
transform 1 0 46100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5133
timestamp 1757982896
transform 1 0 47600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5134
timestamp 1757982896
transform 1 0 49100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5135
timestamp 1757982896
transform 1 0 50600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5136
timestamp 1757982896
transform 1 0 52100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5137
timestamp 1757982896
transform 1 0 53600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5138
timestamp 1757982896
transform 1 0 55100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5139
timestamp 1757982896
transform 1 0 56600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5140
timestamp 1757982896
transform 1 0 58100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5141
timestamp 1757982896
transform 1 0 59600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5142
timestamp 1757982896
transform 1 0 61100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5143
timestamp 1757982896
transform 1 0 62600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5144
timestamp 1757982896
transform 1 0 64100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5145
timestamp 1757982896
transform 1 0 65600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5146
timestamp 1757982896
transform 1 0 67100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5147
timestamp 1757982896
transform 1 0 68600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5148
timestamp 1757982896
transform 1 0 70100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5149
timestamp 1757982896
transform 1 0 71600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5150
timestamp 1757982896
transform 1 0 73100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5151
timestamp 1757982896
transform 1 0 74600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5152
timestamp 1757982896
transform 1 0 76100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5153
timestamp 1757982896
transform 1 0 77600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5154
timestamp 1757982896
transform 1 0 79100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5155
timestamp 1757982896
transform 1 0 80600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5156
timestamp 1757982896
transform 1 0 82100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5157
timestamp 1757982896
transform 1 0 83600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5158
timestamp 1757982896
transform 1 0 85100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5159
timestamp 1757982896
transform 1 0 86600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5160
timestamp 1757982896
transform 1 0 88100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5161
timestamp 1757982896
transform 1 0 89600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5162
timestamp 1757982896
transform 1 0 91100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5163
timestamp 1757982896
transform 1 0 92600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5164
timestamp 1757982896
transform 1 0 94100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5165
timestamp 1757982896
transform 1 0 95600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5166
timestamp 1757982896
transform 1 0 97100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5167
timestamp 1757982896
transform 1 0 98600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5168
timestamp 1757982896
transform 1 0 100100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5169
timestamp 1757982896
transform 1 0 101600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5170
timestamp 1757982896
transform 1 0 103100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5171
timestamp 1757982896
transform 1 0 104600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5172
timestamp 1757982896
transform 1 0 106100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5173
timestamp 1757982896
transform 1 0 107600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5174
timestamp 1757982896
transform 1 0 109100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5175
timestamp 1757982896
transform 1 0 110600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5176
timestamp 1757982896
transform 1 0 112100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5177
timestamp 1757982896
transform 1 0 113600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5178
timestamp 1757982896
transform 1 0 115100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5179
timestamp 1757982896
transform 1 0 116600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5180
timestamp 1757982896
transform 1 0 118100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5181
timestamp 1757982896
transform 1 0 119600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5182
timestamp 1757982896
transform 1 0 121100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5183
timestamp 1757982896
transform 1 0 122600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5184
timestamp 1757982896
transform 1 0 124100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5185
timestamp 1757982896
transform 1 0 125600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5186
timestamp 1757982896
transform 1 0 127100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5187
timestamp 1757982896
transform 1 0 128600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5188
timestamp 1757982896
transform 1 0 130100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5189
timestamp 1757982896
transform 1 0 131600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5190
timestamp 1757982896
transform 1 0 133100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5191
timestamp 1757982896
transform 1 0 134600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5192
timestamp 1757982896
transform 1 0 136100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5193
timestamp 1757982896
transform 1 0 137600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5194
timestamp 1757982896
transform 1 0 139100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5195
timestamp 1757982896
transform 1 0 140600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5196
timestamp 1757982896
transform 1 0 142100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5197
timestamp 1757982896
transform 1 0 143600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5198
timestamp 1757982896
transform 1 0 145100 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5199
timestamp 1757982896
transform 1 0 146600 0 1 -75150
box 1820 -1430 3480 230
use pixel  pixel_5200
timestamp 1757982896
transform 1 0 -1900 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5201
timestamp 1757982896
transform 1 0 -400 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5202
timestamp 1757982896
transform 1 0 1100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5203
timestamp 1757982896
transform 1 0 2600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5204
timestamp 1757982896
transform 1 0 4100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5205
timestamp 1757982896
transform 1 0 5600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5206
timestamp 1757982896
transform 1 0 7100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5207
timestamp 1757982896
transform 1 0 8600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5208
timestamp 1757982896
transform 1 0 10100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5209
timestamp 1757982896
transform 1 0 11600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5210
timestamp 1757982896
transform 1 0 13100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5211
timestamp 1757982896
transform 1 0 14600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5212
timestamp 1757982896
transform 1 0 16100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5213
timestamp 1757982896
transform 1 0 17600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5214
timestamp 1757982896
transform 1 0 19100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5215
timestamp 1757982896
transform 1 0 20600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5216
timestamp 1757982896
transform 1 0 22100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5217
timestamp 1757982896
transform 1 0 23600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5218
timestamp 1757982896
transform 1 0 25100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5219
timestamp 1757982896
transform 1 0 26600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5220
timestamp 1757982896
transform 1 0 28100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5221
timestamp 1757982896
transform 1 0 29600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5222
timestamp 1757982896
transform 1 0 31100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5223
timestamp 1757982896
transform 1 0 32600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5224
timestamp 1757982896
transform 1 0 34100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5225
timestamp 1757982896
transform 1 0 35600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5226
timestamp 1757982896
transform 1 0 37100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5227
timestamp 1757982896
transform 1 0 38600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5228
timestamp 1757982896
transform 1 0 40100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5229
timestamp 1757982896
transform 1 0 41600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5230
timestamp 1757982896
transform 1 0 43100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5231
timestamp 1757982896
transform 1 0 44600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5232
timestamp 1757982896
transform 1 0 46100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5233
timestamp 1757982896
transform 1 0 47600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5234
timestamp 1757982896
transform 1 0 49100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5235
timestamp 1757982896
transform 1 0 50600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5236
timestamp 1757982896
transform 1 0 52100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5237
timestamp 1757982896
transform 1 0 53600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5238
timestamp 1757982896
transform 1 0 55100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5239
timestamp 1757982896
transform 1 0 56600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5240
timestamp 1757982896
transform 1 0 58100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5241
timestamp 1757982896
transform 1 0 59600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5242
timestamp 1757982896
transform 1 0 61100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5243
timestamp 1757982896
transform 1 0 62600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5244
timestamp 1757982896
transform 1 0 64100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5245
timestamp 1757982896
transform 1 0 65600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5246
timestamp 1757982896
transform 1 0 67100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5247
timestamp 1757982896
transform 1 0 68600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5248
timestamp 1757982896
transform 1 0 70100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5249
timestamp 1757982896
transform 1 0 71600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5250
timestamp 1757982896
transform 1 0 73100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5251
timestamp 1757982896
transform 1 0 74600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5252
timestamp 1757982896
transform 1 0 76100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5253
timestamp 1757982896
transform 1 0 77600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5254
timestamp 1757982896
transform 1 0 79100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5255
timestamp 1757982896
transform 1 0 80600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5256
timestamp 1757982896
transform 1 0 82100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5257
timestamp 1757982896
transform 1 0 83600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5258
timestamp 1757982896
transform 1 0 85100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5259
timestamp 1757982896
transform 1 0 86600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5260
timestamp 1757982896
transform 1 0 88100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5261
timestamp 1757982896
transform 1 0 89600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5262
timestamp 1757982896
transform 1 0 91100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5263
timestamp 1757982896
transform 1 0 92600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5264
timestamp 1757982896
transform 1 0 94100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5265
timestamp 1757982896
transform 1 0 95600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5266
timestamp 1757982896
transform 1 0 97100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5267
timestamp 1757982896
transform 1 0 98600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5268
timestamp 1757982896
transform 1 0 100100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5269
timestamp 1757982896
transform 1 0 101600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5270
timestamp 1757982896
transform 1 0 103100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5271
timestamp 1757982896
transform 1 0 104600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5272
timestamp 1757982896
transform 1 0 106100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5273
timestamp 1757982896
transform 1 0 107600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5274
timestamp 1757982896
transform 1 0 109100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5275
timestamp 1757982896
transform 1 0 110600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5276
timestamp 1757982896
transform 1 0 112100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5277
timestamp 1757982896
transform 1 0 113600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5278
timestamp 1757982896
transform 1 0 115100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5279
timestamp 1757982896
transform 1 0 116600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5280
timestamp 1757982896
transform 1 0 118100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5281
timestamp 1757982896
transform 1 0 119600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5282
timestamp 1757982896
transform 1 0 121100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5283
timestamp 1757982896
transform 1 0 122600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5284
timestamp 1757982896
transform 1 0 124100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5285
timestamp 1757982896
transform 1 0 125600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5286
timestamp 1757982896
transform 1 0 127100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5287
timestamp 1757982896
transform 1 0 128600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5288
timestamp 1757982896
transform 1 0 130100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5289
timestamp 1757982896
transform 1 0 131600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5290
timestamp 1757982896
transform 1 0 133100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5291
timestamp 1757982896
transform 1 0 134600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5292
timestamp 1757982896
transform 1 0 136100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5293
timestamp 1757982896
transform 1 0 137600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5294
timestamp 1757982896
transform 1 0 139100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5295
timestamp 1757982896
transform 1 0 140600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5296
timestamp 1757982896
transform 1 0 142100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5297
timestamp 1757982896
transform 1 0 143600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5298
timestamp 1757982896
transform 1 0 145100 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5299
timestamp 1757982896
transform 1 0 146600 0 1 -76650
box 1820 -1430 3480 230
use pixel  pixel_5300
timestamp 1757982896
transform 1 0 -1900 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5301
timestamp 1757982896
transform 1 0 -400 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5302
timestamp 1757982896
transform 1 0 1100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5303
timestamp 1757982896
transform 1 0 2600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5304
timestamp 1757982896
transform 1 0 4100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5305
timestamp 1757982896
transform 1 0 5600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5306
timestamp 1757982896
transform 1 0 7100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5307
timestamp 1757982896
transform 1 0 8600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5308
timestamp 1757982896
transform 1 0 10100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5309
timestamp 1757982896
transform 1 0 11600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5310
timestamp 1757982896
transform 1 0 13100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5311
timestamp 1757982896
transform 1 0 14600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5312
timestamp 1757982896
transform 1 0 16100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5313
timestamp 1757982896
transform 1 0 17600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5314
timestamp 1757982896
transform 1 0 19100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5315
timestamp 1757982896
transform 1 0 20600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5316
timestamp 1757982896
transform 1 0 22100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5317
timestamp 1757982896
transform 1 0 23600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5318
timestamp 1757982896
transform 1 0 25100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5319
timestamp 1757982896
transform 1 0 26600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5320
timestamp 1757982896
transform 1 0 28100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5321
timestamp 1757982896
transform 1 0 29600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5322
timestamp 1757982896
transform 1 0 31100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5323
timestamp 1757982896
transform 1 0 32600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5324
timestamp 1757982896
transform 1 0 34100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5325
timestamp 1757982896
transform 1 0 35600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5326
timestamp 1757982896
transform 1 0 37100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5327
timestamp 1757982896
transform 1 0 38600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5328
timestamp 1757982896
transform 1 0 40100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5329
timestamp 1757982896
transform 1 0 41600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5330
timestamp 1757982896
transform 1 0 43100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5331
timestamp 1757982896
transform 1 0 44600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5332
timestamp 1757982896
transform 1 0 46100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5333
timestamp 1757982896
transform 1 0 47600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5334
timestamp 1757982896
transform 1 0 49100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5335
timestamp 1757982896
transform 1 0 50600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5336
timestamp 1757982896
transform 1 0 52100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5337
timestamp 1757982896
transform 1 0 53600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5338
timestamp 1757982896
transform 1 0 55100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5339
timestamp 1757982896
transform 1 0 56600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5340
timestamp 1757982896
transform 1 0 58100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5341
timestamp 1757982896
transform 1 0 59600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5342
timestamp 1757982896
transform 1 0 61100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5343
timestamp 1757982896
transform 1 0 62600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5344
timestamp 1757982896
transform 1 0 64100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5345
timestamp 1757982896
transform 1 0 65600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5346
timestamp 1757982896
transform 1 0 67100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5347
timestamp 1757982896
transform 1 0 68600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5348
timestamp 1757982896
transform 1 0 70100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5349
timestamp 1757982896
transform 1 0 71600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5350
timestamp 1757982896
transform 1 0 73100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5351
timestamp 1757982896
transform 1 0 74600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5352
timestamp 1757982896
transform 1 0 76100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5353
timestamp 1757982896
transform 1 0 77600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5354
timestamp 1757982896
transform 1 0 79100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5355
timestamp 1757982896
transform 1 0 80600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5356
timestamp 1757982896
transform 1 0 82100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5357
timestamp 1757982896
transform 1 0 83600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5358
timestamp 1757982896
transform 1 0 85100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5359
timestamp 1757982896
transform 1 0 86600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5360
timestamp 1757982896
transform 1 0 88100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5361
timestamp 1757982896
transform 1 0 89600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5362
timestamp 1757982896
transform 1 0 91100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5363
timestamp 1757982896
transform 1 0 92600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5364
timestamp 1757982896
transform 1 0 94100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5365
timestamp 1757982896
transform 1 0 95600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5366
timestamp 1757982896
transform 1 0 97100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5367
timestamp 1757982896
transform 1 0 98600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5368
timestamp 1757982896
transform 1 0 100100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5369
timestamp 1757982896
transform 1 0 101600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5370
timestamp 1757982896
transform 1 0 103100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5371
timestamp 1757982896
transform 1 0 104600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5372
timestamp 1757982896
transform 1 0 106100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5373
timestamp 1757982896
transform 1 0 107600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5374
timestamp 1757982896
transform 1 0 109100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5375
timestamp 1757982896
transform 1 0 110600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5376
timestamp 1757982896
transform 1 0 112100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5377
timestamp 1757982896
transform 1 0 113600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5378
timestamp 1757982896
transform 1 0 115100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5379
timestamp 1757982896
transform 1 0 116600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5380
timestamp 1757982896
transform 1 0 118100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5381
timestamp 1757982896
transform 1 0 119600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5382
timestamp 1757982896
transform 1 0 121100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5383
timestamp 1757982896
transform 1 0 122600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5384
timestamp 1757982896
transform 1 0 124100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5385
timestamp 1757982896
transform 1 0 125600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5386
timestamp 1757982896
transform 1 0 127100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5387
timestamp 1757982896
transform 1 0 128600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5388
timestamp 1757982896
transform 1 0 130100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5389
timestamp 1757982896
transform 1 0 131600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5390
timestamp 1757982896
transform 1 0 133100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5391
timestamp 1757982896
transform 1 0 134600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5392
timestamp 1757982896
transform 1 0 136100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5393
timestamp 1757982896
transform 1 0 137600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5394
timestamp 1757982896
transform 1 0 139100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5395
timestamp 1757982896
transform 1 0 140600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5396
timestamp 1757982896
transform 1 0 142100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5397
timestamp 1757982896
transform 1 0 143600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5398
timestamp 1757982896
transform 1 0 145100 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5399
timestamp 1757982896
transform 1 0 146600 0 1 -78150
box 1820 -1430 3480 230
use pixel  pixel_5400
timestamp 1757982896
transform 1 0 -1900 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5401
timestamp 1757982896
transform 1 0 -400 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5402
timestamp 1757982896
transform 1 0 1100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5403
timestamp 1757982896
transform 1 0 2600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5404
timestamp 1757982896
transform 1 0 4100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5405
timestamp 1757982896
transform 1 0 5600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5406
timestamp 1757982896
transform 1 0 7100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5407
timestamp 1757982896
transform 1 0 8600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5408
timestamp 1757982896
transform 1 0 10100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5409
timestamp 1757982896
transform 1 0 11600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5410
timestamp 1757982896
transform 1 0 13100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5411
timestamp 1757982896
transform 1 0 14600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5412
timestamp 1757982896
transform 1 0 16100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5413
timestamp 1757982896
transform 1 0 17600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5414
timestamp 1757982896
transform 1 0 19100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5415
timestamp 1757982896
transform 1 0 20600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5416
timestamp 1757982896
transform 1 0 22100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5417
timestamp 1757982896
transform 1 0 23600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5418
timestamp 1757982896
transform 1 0 25100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5419
timestamp 1757982896
transform 1 0 26600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5420
timestamp 1757982896
transform 1 0 28100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5421
timestamp 1757982896
transform 1 0 29600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5422
timestamp 1757982896
transform 1 0 31100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5423
timestamp 1757982896
transform 1 0 32600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5424
timestamp 1757982896
transform 1 0 34100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5425
timestamp 1757982896
transform 1 0 35600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5426
timestamp 1757982896
transform 1 0 37100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5427
timestamp 1757982896
transform 1 0 38600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5428
timestamp 1757982896
transform 1 0 40100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5429
timestamp 1757982896
transform 1 0 41600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5430
timestamp 1757982896
transform 1 0 43100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5431
timestamp 1757982896
transform 1 0 44600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5432
timestamp 1757982896
transform 1 0 46100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5433
timestamp 1757982896
transform 1 0 47600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5434
timestamp 1757982896
transform 1 0 49100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5435
timestamp 1757982896
transform 1 0 50600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5436
timestamp 1757982896
transform 1 0 52100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5437
timestamp 1757982896
transform 1 0 53600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5438
timestamp 1757982896
transform 1 0 55100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5439
timestamp 1757982896
transform 1 0 56600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5440
timestamp 1757982896
transform 1 0 58100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5441
timestamp 1757982896
transform 1 0 59600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5442
timestamp 1757982896
transform 1 0 61100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5443
timestamp 1757982896
transform 1 0 62600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5444
timestamp 1757982896
transform 1 0 64100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5445
timestamp 1757982896
transform 1 0 65600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5446
timestamp 1757982896
transform 1 0 67100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5447
timestamp 1757982896
transform 1 0 68600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5448
timestamp 1757982896
transform 1 0 70100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5449
timestamp 1757982896
transform 1 0 71600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5450
timestamp 1757982896
transform 1 0 73100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5451
timestamp 1757982896
transform 1 0 74600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5452
timestamp 1757982896
transform 1 0 76100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5453
timestamp 1757982896
transform 1 0 77600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5454
timestamp 1757982896
transform 1 0 79100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5455
timestamp 1757982896
transform 1 0 80600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5456
timestamp 1757982896
transform 1 0 82100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5457
timestamp 1757982896
transform 1 0 83600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5458
timestamp 1757982896
transform 1 0 85100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5459
timestamp 1757982896
transform 1 0 86600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5460
timestamp 1757982896
transform 1 0 88100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5461
timestamp 1757982896
transform 1 0 89600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5462
timestamp 1757982896
transform 1 0 91100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5463
timestamp 1757982896
transform 1 0 92600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5464
timestamp 1757982896
transform 1 0 94100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5465
timestamp 1757982896
transform 1 0 95600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5466
timestamp 1757982896
transform 1 0 97100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5467
timestamp 1757982896
transform 1 0 98600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5468
timestamp 1757982896
transform 1 0 100100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5469
timestamp 1757982896
transform 1 0 101600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5470
timestamp 1757982896
transform 1 0 103100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5471
timestamp 1757982896
transform 1 0 104600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5472
timestamp 1757982896
transform 1 0 106100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5473
timestamp 1757982896
transform 1 0 107600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5474
timestamp 1757982896
transform 1 0 109100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5475
timestamp 1757982896
transform 1 0 110600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5476
timestamp 1757982896
transform 1 0 112100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5477
timestamp 1757982896
transform 1 0 113600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5478
timestamp 1757982896
transform 1 0 115100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5479
timestamp 1757982896
transform 1 0 116600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5480
timestamp 1757982896
transform 1 0 118100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5481
timestamp 1757982896
transform 1 0 119600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5482
timestamp 1757982896
transform 1 0 121100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5483
timestamp 1757982896
transform 1 0 122600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5484
timestamp 1757982896
transform 1 0 124100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5485
timestamp 1757982896
transform 1 0 125600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5486
timestamp 1757982896
transform 1 0 127100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5487
timestamp 1757982896
transform 1 0 128600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5488
timestamp 1757982896
transform 1 0 130100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5489
timestamp 1757982896
transform 1 0 131600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5490
timestamp 1757982896
transform 1 0 133100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5491
timestamp 1757982896
transform 1 0 134600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5492
timestamp 1757982896
transform 1 0 136100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5493
timestamp 1757982896
transform 1 0 137600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5494
timestamp 1757982896
transform 1 0 139100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5495
timestamp 1757982896
transform 1 0 140600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5496
timestamp 1757982896
transform 1 0 142100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5497
timestamp 1757982896
transform 1 0 143600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5498
timestamp 1757982896
transform 1 0 145100 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5499
timestamp 1757982896
transform 1 0 146600 0 1 -79650
box 1820 -1430 3480 230
use pixel  pixel_5500
timestamp 1757982896
transform 1 0 -1900 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5501
timestamp 1757982896
transform 1 0 -400 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5502
timestamp 1757982896
transform 1 0 1100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5503
timestamp 1757982896
transform 1 0 2600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5504
timestamp 1757982896
transform 1 0 4100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5505
timestamp 1757982896
transform 1 0 5600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5506
timestamp 1757982896
transform 1 0 7100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5507
timestamp 1757982896
transform 1 0 8600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5508
timestamp 1757982896
transform 1 0 10100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5509
timestamp 1757982896
transform 1 0 11600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5510
timestamp 1757982896
transform 1 0 13100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5511
timestamp 1757982896
transform 1 0 14600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5512
timestamp 1757982896
transform 1 0 16100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5513
timestamp 1757982896
transform 1 0 17600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5514
timestamp 1757982896
transform 1 0 19100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5515
timestamp 1757982896
transform 1 0 20600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5516
timestamp 1757982896
transform 1 0 22100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5517
timestamp 1757982896
transform 1 0 23600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5518
timestamp 1757982896
transform 1 0 25100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5519
timestamp 1757982896
transform 1 0 26600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5520
timestamp 1757982896
transform 1 0 28100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5521
timestamp 1757982896
transform 1 0 29600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5522
timestamp 1757982896
transform 1 0 31100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5523
timestamp 1757982896
transform 1 0 32600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5524
timestamp 1757982896
transform 1 0 34100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5525
timestamp 1757982896
transform 1 0 35600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5526
timestamp 1757982896
transform 1 0 37100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5527
timestamp 1757982896
transform 1 0 38600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5528
timestamp 1757982896
transform 1 0 40100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5529
timestamp 1757982896
transform 1 0 41600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5530
timestamp 1757982896
transform 1 0 43100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5531
timestamp 1757982896
transform 1 0 44600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5532
timestamp 1757982896
transform 1 0 46100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5533
timestamp 1757982896
transform 1 0 47600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5534
timestamp 1757982896
transform 1 0 49100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5535
timestamp 1757982896
transform 1 0 50600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5536
timestamp 1757982896
transform 1 0 52100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5537
timestamp 1757982896
transform 1 0 53600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5538
timestamp 1757982896
transform 1 0 55100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5539
timestamp 1757982896
transform 1 0 56600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5540
timestamp 1757982896
transform 1 0 58100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5541
timestamp 1757982896
transform 1 0 59600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5542
timestamp 1757982896
transform 1 0 61100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5543
timestamp 1757982896
transform 1 0 62600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5544
timestamp 1757982896
transform 1 0 64100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5545
timestamp 1757982896
transform 1 0 65600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5546
timestamp 1757982896
transform 1 0 67100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5547
timestamp 1757982896
transform 1 0 68600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5548
timestamp 1757982896
transform 1 0 70100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5549
timestamp 1757982896
transform 1 0 71600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5550
timestamp 1757982896
transform 1 0 73100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5551
timestamp 1757982896
transform 1 0 74600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5552
timestamp 1757982896
transform 1 0 76100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5553
timestamp 1757982896
transform 1 0 77600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5554
timestamp 1757982896
transform 1 0 79100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5555
timestamp 1757982896
transform 1 0 80600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5556
timestamp 1757982896
transform 1 0 82100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5557
timestamp 1757982896
transform 1 0 83600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5558
timestamp 1757982896
transform 1 0 85100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5559
timestamp 1757982896
transform 1 0 86600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5560
timestamp 1757982896
transform 1 0 88100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5561
timestamp 1757982896
transform 1 0 89600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5562
timestamp 1757982896
transform 1 0 91100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5563
timestamp 1757982896
transform 1 0 92600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5564
timestamp 1757982896
transform 1 0 94100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5565
timestamp 1757982896
transform 1 0 95600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5566
timestamp 1757982896
transform 1 0 97100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5567
timestamp 1757982896
transform 1 0 98600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5568
timestamp 1757982896
transform 1 0 100100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5569
timestamp 1757982896
transform 1 0 101600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5570
timestamp 1757982896
transform 1 0 103100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5571
timestamp 1757982896
transform 1 0 104600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5572
timestamp 1757982896
transform 1 0 106100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5573
timestamp 1757982896
transform 1 0 107600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5574
timestamp 1757982896
transform 1 0 109100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5575
timestamp 1757982896
transform 1 0 110600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5576
timestamp 1757982896
transform 1 0 112100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5577
timestamp 1757982896
transform 1 0 113600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5578
timestamp 1757982896
transform 1 0 115100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5579
timestamp 1757982896
transform 1 0 116600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5580
timestamp 1757982896
transform 1 0 118100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5581
timestamp 1757982896
transform 1 0 119600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5582
timestamp 1757982896
transform 1 0 121100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5583
timestamp 1757982896
transform 1 0 122600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5584
timestamp 1757982896
transform 1 0 124100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5585
timestamp 1757982896
transform 1 0 125600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5586
timestamp 1757982896
transform 1 0 127100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5587
timestamp 1757982896
transform 1 0 128600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5588
timestamp 1757982896
transform 1 0 130100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5589
timestamp 1757982896
transform 1 0 131600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5590
timestamp 1757982896
transform 1 0 133100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5591
timestamp 1757982896
transform 1 0 134600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5592
timestamp 1757982896
transform 1 0 136100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5593
timestamp 1757982896
transform 1 0 137600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5594
timestamp 1757982896
transform 1 0 139100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5595
timestamp 1757982896
transform 1 0 140600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5596
timestamp 1757982896
transform 1 0 142100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5597
timestamp 1757982896
transform 1 0 143600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5598
timestamp 1757982896
transform 1 0 145100 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5599
timestamp 1757982896
transform 1 0 146600 0 1 -81150
box 1820 -1430 3480 230
use pixel  pixel_5600
timestamp 1757982896
transform 1 0 -1900 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5601
timestamp 1757982896
transform 1 0 -400 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5602
timestamp 1757982896
transform 1 0 1100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5603
timestamp 1757982896
transform 1 0 2600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5604
timestamp 1757982896
transform 1 0 4100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5605
timestamp 1757982896
transform 1 0 5600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5606
timestamp 1757982896
transform 1 0 7100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5607
timestamp 1757982896
transform 1 0 8600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5608
timestamp 1757982896
transform 1 0 10100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5609
timestamp 1757982896
transform 1 0 11600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5610
timestamp 1757982896
transform 1 0 13100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5611
timestamp 1757982896
transform 1 0 14600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5612
timestamp 1757982896
transform 1 0 16100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5613
timestamp 1757982896
transform 1 0 17600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5614
timestamp 1757982896
transform 1 0 19100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5615
timestamp 1757982896
transform 1 0 20600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5616
timestamp 1757982896
transform 1 0 22100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5617
timestamp 1757982896
transform 1 0 23600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5618
timestamp 1757982896
transform 1 0 25100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5619
timestamp 1757982896
transform 1 0 26600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5620
timestamp 1757982896
transform 1 0 28100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5621
timestamp 1757982896
transform 1 0 29600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5622
timestamp 1757982896
transform 1 0 31100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5623
timestamp 1757982896
transform 1 0 32600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5624
timestamp 1757982896
transform 1 0 34100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5625
timestamp 1757982896
transform 1 0 35600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5626
timestamp 1757982896
transform 1 0 37100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5627
timestamp 1757982896
transform 1 0 38600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5628
timestamp 1757982896
transform 1 0 40100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5629
timestamp 1757982896
transform 1 0 41600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5630
timestamp 1757982896
transform 1 0 43100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5631
timestamp 1757982896
transform 1 0 44600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5632
timestamp 1757982896
transform 1 0 46100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5633
timestamp 1757982896
transform 1 0 47600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5634
timestamp 1757982896
transform 1 0 49100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5635
timestamp 1757982896
transform 1 0 50600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5636
timestamp 1757982896
transform 1 0 52100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5637
timestamp 1757982896
transform 1 0 53600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5638
timestamp 1757982896
transform 1 0 55100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5639
timestamp 1757982896
transform 1 0 56600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5640
timestamp 1757982896
transform 1 0 58100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5641
timestamp 1757982896
transform 1 0 59600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5642
timestamp 1757982896
transform 1 0 61100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5643
timestamp 1757982896
transform 1 0 62600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5644
timestamp 1757982896
transform 1 0 64100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5645
timestamp 1757982896
transform 1 0 65600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5646
timestamp 1757982896
transform 1 0 67100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5647
timestamp 1757982896
transform 1 0 68600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5648
timestamp 1757982896
transform 1 0 70100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5649
timestamp 1757982896
transform 1 0 71600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5650
timestamp 1757982896
transform 1 0 73100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5651
timestamp 1757982896
transform 1 0 74600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5652
timestamp 1757982896
transform 1 0 76100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5653
timestamp 1757982896
transform 1 0 77600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5654
timestamp 1757982896
transform 1 0 79100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5655
timestamp 1757982896
transform 1 0 80600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5656
timestamp 1757982896
transform 1 0 82100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5657
timestamp 1757982896
transform 1 0 83600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5658
timestamp 1757982896
transform 1 0 85100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5659
timestamp 1757982896
transform 1 0 86600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5660
timestamp 1757982896
transform 1 0 88100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5661
timestamp 1757982896
transform 1 0 89600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5662
timestamp 1757982896
transform 1 0 91100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5663
timestamp 1757982896
transform 1 0 92600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5664
timestamp 1757982896
transform 1 0 94100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5665
timestamp 1757982896
transform 1 0 95600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5666
timestamp 1757982896
transform 1 0 97100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5667
timestamp 1757982896
transform 1 0 98600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5668
timestamp 1757982896
transform 1 0 100100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5669
timestamp 1757982896
transform 1 0 101600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5670
timestamp 1757982896
transform 1 0 103100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5671
timestamp 1757982896
transform 1 0 104600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5672
timestamp 1757982896
transform 1 0 106100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5673
timestamp 1757982896
transform 1 0 107600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5674
timestamp 1757982896
transform 1 0 109100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5675
timestamp 1757982896
transform 1 0 110600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5676
timestamp 1757982896
transform 1 0 112100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5677
timestamp 1757982896
transform 1 0 113600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5678
timestamp 1757982896
transform 1 0 115100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5679
timestamp 1757982896
transform 1 0 116600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5680
timestamp 1757982896
transform 1 0 118100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5681
timestamp 1757982896
transform 1 0 119600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5682
timestamp 1757982896
transform 1 0 121100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5683
timestamp 1757982896
transform 1 0 122600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5684
timestamp 1757982896
transform 1 0 124100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5685
timestamp 1757982896
transform 1 0 125600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5686
timestamp 1757982896
transform 1 0 127100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5687
timestamp 1757982896
transform 1 0 128600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5688
timestamp 1757982896
transform 1 0 130100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5689
timestamp 1757982896
transform 1 0 131600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5690
timestamp 1757982896
transform 1 0 133100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5691
timestamp 1757982896
transform 1 0 134600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5692
timestamp 1757982896
transform 1 0 136100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5693
timestamp 1757982896
transform 1 0 137600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5694
timestamp 1757982896
transform 1 0 139100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5695
timestamp 1757982896
transform 1 0 140600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5696
timestamp 1757982896
transform 1 0 142100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5697
timestamp 1757982896
transform 1 0 143600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5698
timestamp 1757982896
transform 1 0 145100 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5699
timestamp 1757982896
transform 1 0 146600 0 1 -82650
box 1820 -1430 3480 230
use pixel  pixel_5700
timestamp 1757982896
transform 1 0 -1900 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5701
timestamp 1757982896
transform 1 0 -400 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5702
timestamp 1757982896
transform 1 0 1100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5703
timestamp 1757982896
transform 1 0 2600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5704
timestamp 1757982896
transform 1 0 4100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5705
timestamp 1757982896
transform 1 0 5600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5706
timestamp 1757982896
transform 1 0 7100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5707
timestamp 1757982896
transform 1 0 8600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5708
timestamp 1757982896
transform 1 0 10100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5709
timestamp 1757982896
transform 1 0 11600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5710
timestamp 1757982896
transform 1 0 13100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5711
timestamp 1757982896
transform 1 0 14600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5712
timestamp 1757982896
transform 1 0 16100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5713
timestamp 1757982896
transform 1 0 17600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5714
timestamp 1757982896
transform 1 0 19100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5715
timestamp 1757982896
transform 1 0 20600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5716
timestamp 1757982896
transform 1 0 22100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5717
timestamp 1757982896
transform 1 0 23600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5718
timestamp 1757982896
transform 1 0 25100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5719
timestamp 1757982896
transform 1 0 26600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5720
timestamp 1757982896
transform 1 0 28100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5721
timestamp 1757982896
transform 1 0 29600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5722
timestamp 1757982896
transform 1 0 31100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5723
timestamp 1757982896
transform 1 0 32600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5724
timestamp 1757982896
transform 1 0 34100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5725
timestamp 1757982896
transform 1 0 35600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5726
timestamp 1757982896
transform 1 0 37100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5727
timestamp 1757982896
transform 1 0 38600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5728
timestamp 1757982896
transform 1 0 40100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5729
timestamp 1757982896
transform 1 0 41600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5730
timestamp 1757982896
transform 1 0 43100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5731
timestamp 1757982896
transform 1 0 44600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5732
timestamp 1757982896
transform 1 0 46100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5733
timestamp 1757982896
transform 1 0 47600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5734
timestamp 1757982896
transform 1 0 49100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5735
timestamp 1757982896
transform 1 0 50600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5736
timestamp 1757982896
transform 1 0 52100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5737
timestamp 1757982896
transform 1 0 53600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5738
timestamp 1757982896
transform 1 0 55100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5739
timestamp 1757982896
transform 1 0 56600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5740
timestamp 1757982896
transform 1 0 58100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5741
timestamp 1757982896
transform 1 0 59600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5742
timestamp 1757982896
transform 1 0 61100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5743
timestamp 1757982896
transform 1 0 62600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5744
timestamp 1757982896
transform 1 0 64100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5745
timestamp 1757982896
transform 1 0 65600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5746
timestamp 1757982896
transform 1 0 67100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5747
timestamp 1757982896
transform 1 0 68600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5748
timestamp 1757982896
transform 1 0 70100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5749
timestamp 1757982896
transform 1 0 71600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5750
timestamp 1757982896
transform 1 0 73100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5751
timestamp 1757982896
transform 1 0 74600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5752
timestamp 1757982896
transform 1 0 76100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5753
timestamp 1757982896
transform 1 0 77600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5754
timestamp 1757982896
transform 1 0 79100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5755
timestamp 1757982896
transform 1 0 80600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5756
timestamp 1757982896
transform 1 0 82100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5757
timestamp 1757982896
transform 1 0 83600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5758
timestamp 1757982896
transform 1 0 85100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5759
timestamp 1757982896
transform 1 0 86600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5760
timestamp 1757982896
transform 1 0 88100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5761
timestamp 1757982896
transform 1 0 89600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5762
timestamp 1757982896
transform 1 0 91100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5763
timestamp 1757982896
transform 1 0 92600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5764
timestamp 1757982896
transform 1 0 94100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5765
timestamp 1757982896
transform 1 0 95600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5766
timestamp 1757982896
transform 1 0 97100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5767
timestamp 1757982896
transform 1 0 98600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5768
timestamp 1757982896
transform 1 0 100100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5769
timestamp 1757982896
transform 1 0 101600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5770
timestamp 1757982896
transform 1 0 103100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5771
timestamp 1757982896
transform 1 0 104600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5772
timestamp 1757982896
transform 1 0 106100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5773
timestamp 1757982896
transform 1 0 107600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5774
timestamp 1757982896
transform 1 0 109100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5775
timestamp 1757982896
transform 1 0 110600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5776
timestamp 1757982896
transform 1 0 112100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5777
timestamp 1757982896
transform 1 0 113600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5778
timestamp 1757982896
transform 1 0 115100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5779
timestamp 1757982896
transform 1 0 116600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5780
timestamp 1757982896
transform 1 0 118100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5781
timestamp 1757982896
transform 1 0 119600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5782
timestamp 1757982896
transform 1 0 121100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5783
timestamp 1757982896
transform 1 0 122600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5784
timestamp 1757982896
transform 1 0 124100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5785
timestamp 1757982896
transform 1 0 125600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5786
timestamp 1757982896
transform 1 0 127100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5787
timestamp 1757982896
transform 1 0 128600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5788
timestamp 1757982896
transform 1 0 130100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5789
timestamp 1757982896
transform 1 0 131600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5790
timestamp 1757982896
transform 1 0 133100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5791
timestamp 1757982896
transform 1 0 134600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5792
timestamp 1757982896
transform 1 0 136100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5793
timestamp 1757982896
transform 1 0 137600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5794
timestamp 1757982896
transform 1 0 139100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5795
timestamp 1757982896
transform 1 0 140600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5796
timestamp 1757982896
transform 1 0 142100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5797
timestamp 1757982896
transform 1 0 143600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5798
timestamp 1757982896
transform 1 0 145100 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5799
timestamp 1757982896
transform 1 0 146600 0 1 -84150
box 1820 -1430 3480 230
use pixel  pixel_5800
timestamp 1757982896
transform 1 0 -1900 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5801
timestamp 1757982896
transform 1 0 -400 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5802
timestamp 1757982896
transform 1 0 1100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5803
timestamp 1757982896
transform 1 0 2600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5804
timestamp 1757982896
transform 1 0 4100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5805
timestamp 1757982896
transform 1 0 5600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5806
timestamp 1757982896
transform 1 0 7100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5807
timestamp 1757982896
transform 1 0 8600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5808
timestamp 1757982896
transform 1 0 10100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5809
timestamp 1757982896
transform 1 0 11600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5810
timestamp 1757982896
transform 1 0 13100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5811
timestamp 1757982896
transform 1 0 14600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5812
timestamp 1757982896
transform 1 0 16100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5813
timestamp 1757982896
transform 1 0 17600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5814
timestamp 1757982896
transform 1 0 19100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5815
timestamp 1757982896
transform 1 0 20600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5816
timestamp 1757982896
transform 1 0 22100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5817
timestamp 1757982896
transform 1 0 23600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5818
timestamp 1757982896
transform 1 0 25100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5819
timestamp 1757982896
transform 1 0 26600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5820
timestamp 1757982896
transform 1 0 28100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5821
timestamp 1757982896
transform 1 0 29600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5822
timestamp 1757982896
transform 1 0 31100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5823
timestamp 1757982896
transform 1 0 32600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5824
timestamp 1757982896
transform 1 0 34100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5825
timestamp 1757982896
transform 1 0 35600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5826
timestamp 1757982896
transform 1 0 37100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5827
timestamp 1757982896
transform 1 0 38600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5828
timestamp 1757982896
transform 1 0 40100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5829
timestamp 1757982896
transform 1 0 41600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5830
timestamp 1757982896
transform 1 0 43100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5831
timestamp 1757982896
transform 1 0 44600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5832
timestamp 1757982896
transform 1 0 46100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5833
timestamp 1757982896
transform 1 0 47600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5834
timestamp 1757982896
transform 1 0 49100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5835
timestamp 1757982896
transform 1 0 50600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5836
timestamp 1757982896
transform 1 0 52100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5837
timestamp 1757982896
transform 1 0 53600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5838
timestamp 1757982896
transform 1 0 55100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5839
timestamp 1757982896
transform 1 0 56600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5840
timestamp 1757982896
transform 1 0 58100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5841
timestamp 1757982896
transform 1 0 59600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5842
timestamp 1757982896
transform 1 0 61100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5843
timestamp 1757982896
transform 1 0 62600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5844
timestamp 1757982896
transform 1 0 64100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5845
timestamp 1757982896
transform 1 0 65600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5846
timestamp 1757982896
transform 1 0 67100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5847
timestamp 1757982896
transform 1 0 68600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5848
timestamp 1757982896
transform 1 0 70100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5849
timestamp 1757982896
transform 1 0 71600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5850
timestamp 1757982896
transform 1 0 73100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5851
timestamp 1757982896
transform 1 0 74600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5852
timestamp 1757982896
transform 1 0 76100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5853
timestamp 1757982896
transform 1 0 77600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5854
timestamp 1757982896
transform 1 0 79100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5855
timestamp 1757982896
transform 1 0 80600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5856
timestamp 1757982896
transform 1 0 82100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5857
timestamp 1757982896
transform 1 0 83600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5858
timestamp 1757982896
transform 1 0 85100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5859
timestamp 1757982896
transform 1 0 86600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5860
timestamp 1757982896
transform 1 0 88100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5861
timestamp 1757982896
transform 1 0 89600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5862
timestamp 1757982896
transform 1 0 91100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5863
timestamp 1757982896
transform 1 0 92600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5864
timestamp 1757982896
transform 1 0 94100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5865
timestamp 1757982896
transform 1 0 95600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5866
timestamp 1757982896
transform 1 0 97100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5867
timestamp 1757982896
transform 1 0 98600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5868
timestamp 1757982896
transform 1 0 100100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5869
timestamp 1757982896
transform 1 0 101600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5870
timestamp 1757982896
transform 1 0 103100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5871
timestamp 1757982896
transform 1 0 104600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5872
timestamp 1757982896
transform 1 0 106100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5873
timestamp 1757982896
transform 1 0 107600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5874
timestamp 1757982896
transform 1 0 109100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5875
timestamp 1757982896
transform 1 0 110600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5876
timestamp 1757982896
transform 1 0 112100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5877
timestamp 1757982896
transform 1 0 113600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5878
timestamp 1757982896
transform 1 0 115100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5879
timestamp 1757982896
transform 1 0 116600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5880
timestamp 1757982896
transform 1 0 118100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5881
timestamp 1757982896
transform 1 0 119600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5882
timestamp 1757982896
transform 1 0 121100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5883
timestamp 1757982896
transform 1 0 122600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5884
timestamp 1757982896
transform 1 0 124100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5885
timestamp 1757982896
transform 1 0 125600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5886
timestamp 1757982896
transform 1 0 127100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5887
timestamp 1757982896
transform 1 0 128600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5888
timestamp 1757982896
transform 1 0 130100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5889
timestamp 1757982896
transform 1 0 131600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5890
timestamp 1757982896
transform 1 0 133100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5891
timestamp 1757982896
transform 1 0 134600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5892
timestamp 1757982896
transform 1 0 136100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5893
timestamp 1757982896
transform 1 0 137600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5894
timestamp 1757982896
transform 1 0 139100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5895
timestamp 1757982896
transform 1 0 140600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5896
timestamp 1757982896
transform 1 0 142100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5897
timestamp 1757982896
transform 1 0 143600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5898
timestamp 1757982896
transform 1 0 145100 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5899
timestamp 1757982896
transform 1 0 146600 0 1 -85650
box 1820 -1430 3480 230
use pixel  pixel_5900
timestamp 1757982896
transform 1 0 -1900 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5901
timestamp 1757982896
transform 1 0 -400 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5902
timestamp 1757982896
transform 1 0 1100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5903
timestamp 1757982896
transform 1 0 2600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5904
timestamp 1757982896
transform 1 0 4100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5905
timestamp 1757982896
transform 1 0 5600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5906
timestamp 1757982896
transform 1 0 7100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5907
timestamp 1757982896
transform 1 0 8600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5908
timestamp 1757982896
transform 1 0 10100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5909
timestamp 1757982896
transform 1 0 11600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5910
timestamp 1757982896
transform 1 0 13100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5911
timestamp 1757982896
transform 1 0 14600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5912
timestamp 1757982896
transform 1 0 16100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5913
timestamp 1757982896
transform 1 0 17600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5914
timestamp 1757982896
transform 1 0 19100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5915
timestamp 1757982896
transform 1 0 20600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5916
timestamp 1757982896
transform 1 0 22100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5917
timestamp 1757982896
transform 1 0 23600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5918
timestamp 1757982896
transform 1 0 25100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5919
timestamp 1757982896
transform 1 0 26600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5920
timestamp 1757982896
transform 1 0 28100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5921
timestamp 1757982896
transform 1 0 29600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5922
timestamp 1757982896
transform 1 0 31100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5923
timestamp 1757982896
transform 1 0 32600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5924
timestamp 1757982896
transform 1 0 34100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5925
timestamp 1757982896
transform 1 0 35600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5926
timestamp 1757982896
transform 1 0 37100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5927
timestamp 1757982896
transform 1 0 38600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5928
timestamp 1757982896
transform 1 0 40100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5929
timestamp 1757982896
transform 1 0 41600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5930
timestamp 1757982896
transform 1 0 43100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5931
timestamp 1757982896
transform 1 0 44600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5932
timestamp 1757982896
transform 1 0 46100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5933
timestamp 1757982896
transform 1 0 47600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5934
timestamp 1757982896
transform 1 0 49100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5935
timestamp 1757982896
transform 1 0 50600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5936
timestamp 1757982896
transform 1 0 52100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5937
timestamp 1757982896
transform 1 0 53600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5938
timestamp 1757982896
transform 1 0 55100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5939
timestamp 1757982896
transform 1 0 56600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5940
timestamp 1757982896
transform 1 0 58100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5941
timestamp 1757982896
transform 1 0 59600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5942
timestamp 1757982896
transform 1 0 61100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5943
timestamp 1757982896
transform 1 0 62600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5944
timestamp 1757982896
transform 1 0 64100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5945
timestamp 1757982896
transform 1 0 65600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5946
timestamp 1757982896
transform 1 0 67100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5947
timestamp 1757982896
transform 1 0 68600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5948
timestamp 1757982896
transform 1 0 70100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5949
timestamp 1757982896
transform 1 0 71600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5950
timestamp 1757982896
transform 1 0 73100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5951
timestamp 1757982896
transform 1 0 74600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5952
timestamp 1757982896
transform 1 0 76100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5953
timestamp 1757982896
transform 1 0 77600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5954
timestamp 1757982896
transform 1 0 79100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5955
timestamp 1757982896
transform 1 0 80600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5956
timestamp 1757982896
transform 1 0 82100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5957
timestamp 1757982896
transform 1 0 83600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5958
timestamp 1757982896
transform 1 0 85100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5959
timestamp 1757982896
transform 1 0 86600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5960
timestamp 1757982896
transform 1 0 88100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5961
timestamp 1757982896
transform 1 0 89600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5962
timestamp 1757982896
transform 1 0 91100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5963
timestamp 1757982896
transform 1 0 92600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5964
timestamp 1757982896
transform 1 0 94100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5965
timestamp 1757982896
transform 1 0 95600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5966
timestamp 1757982896
transform 1 0 97100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5967
timestamp 1757982896
transform 1 0 98600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5968
timestamp 1757982896
transform 1 0 100100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5969
timestamp 1757982896
transform 1 0 101600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5970
timestamp 1757982896
transform 1 0 103100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5971
timestamp 1757982896
transform 1 0 104600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5972
timestamp 1757982896
transform 1 0 106100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5973
timestamp 1757982896
transform 1 0 107600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5974
timestamp 1757982896
transform 1 0 109100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5975
timestamp 1757982896
transform 1 0 110600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5976
timestamp 1757982896
transform 1 0 112100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5977
timestamp 1757982896
transform 1 0 113600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5978
timestamp 1757982896
transform 1 0 115100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5979
timestamp 1757982896
transform 1 0 116600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5980
timestamp 1757982896
transform 1 0 118100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5981
timestamp 1757982896
transform 1 0 119600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5982
timestamp 1757982896
transform 1 0 121100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5983
timestamp 1757982896
transform 1 0 122600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5984
timestamp 1757982896
transform 1 0 124100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5985
timestamp 1757982896
transform 1 0 125600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5986
timestamp 1757982896
transform 1 0 127100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5987
timestamp 1757982896
transform 1 0 128600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5988
timestamp 1757982896
transform 1 0 130100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5989
timestamp 1757982896
transform 1 0 131600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5990
timestamp 1757982896
transform 1 0 133100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5991
timestamp 1757982896
transform 1 0 134600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5992
timestamp 1757982896
transform 1 0 136100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5993
timestamp 1757982896
transform 1 0 137600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5994
timestamp 1757982896
transform 1 0 139100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5995
timestamp 1757982896
transform 1 0 140600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5996
timestamp 1757982896
transform 1 0 142100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5997
timestamp 1757982896
transform 1 0 143600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5998
timestamp 1757982896
transform 1 0 145100 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_5999
timestamp 1757982896
transform 1 0 146600 0 1 -87150
box 1820 -1430 3480 230
use pixel  pixel_6000
timestamp 1757982896
transform 1 0 -1900 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6001
timestamp 1757982896
transform 1 0 -400 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6002
timestamp 1757982896
transform 1 0 1100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6003
timestamp 1757982896
transform 1 0 2600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6004
timestamp 1757982896
transform 1 0 4100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6005
timestamp 1757982896
transform 1 0 5600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6006
timestamp 1757982896
transform 1 0 7100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6007
timestamp 1757982896
transform 1 0 8600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6008
timestamp 1757982896
transform 1 0 10100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6009
timestamp 1757982896
transform 1 0 11600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6010
timestamp 1757982896
transform 1 0 13100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6011
timestamp 1757982896
transform 1 0 14600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6012
timestamp 1757982896
transform 1 0 16100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6013
timestamp 1757982896
transform 1 0 17600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6014
timestamp 1757982896
transform 1 0 19100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6015
timestamp 1757982896
transform 1 0 20600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6016
timestamp 1757982896
transform 1 0 22100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6017
timestamp 1757982896
transform 1 0 23600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6018
timestamp 1757982896
transform 1 0 25100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6019
timestamp 1757982896
transform 1 0 26600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6020
timestamp 1757982896
transform 1 0 28100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6021
timestamp 1757982896
transform 1 0 29600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6022
timestamp 1757982896
transform 1 0 31100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6023
timestamp 1757982896
transform 1 0 32600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6024
timestamp 1757982896
transform 1 0 34100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6025
timestamp 1757982896
transform 1 0 35600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6026
timestamp 1757982896
transform 1 0 37100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6027
timestamp 1757982896
transform 1 0 38600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6028
timestamp 1757982896
transform 1 0 40100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6029
timestamp 1757982896
transform 1 0 41600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6030
timestamp 1757982896
transform 1 0 43100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6031
timestamp 1757982896
transform 1 0 44600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6032
timestamp 1757982896
transform 1 0 46100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6033
timestamp 1757982896
transform 1 0 47600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6034
timestamp 1757982896
transform 1 0 49100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6035
timestamp 1757982896
transform 1 0 50600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6036
timestamp 1757982896
transform 1 0 52100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6037
timestamp 1757982896
transform 1 0 53600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6038
timestamp 1757982896
transform 1 0 55100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6039
timestamp 1757982896
transform 1 0 56600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6040
timestamp 1757982896
transform 1 0 58100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6041
timestamp 1757982896
transform 1 0 59600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6042
timestamp 1757982896
transform 1 0 61100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6043
timestamp 1757982896
transform 1 0 62600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6044
timestamp 1757982896
transform 1 0 64100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6045
timestamp 1757982896
transform 1 0 65600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6046
timestamp 1757982896
transform 1 0 67100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6047
timestamp 1757982896
transform 1 0 68600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6048
timestamp 1757982896
transform 1 0 70100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6049
timestamp 1757982896
transform 1 0 71600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6050
timestamp 1757982896
transform 1 0 73100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6051
timestamp 1757982896
transform 1 0 74600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6052
timestamp 1757982896
transform 1 0 76100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6053
timestamp 1757982896
transform 1 0 77600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6054
timestamp 1757982896
transform 1 0 79100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6055
timestamp 1757982896
transform 1 0 80600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6056
timestamp 1757982896
transform 1 0 82100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6057
timestamp 1757982896
transform 1 0 83600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6058
timestamp 1757982896
transform 1 0 85100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6059
timestamp 1757982896
transform 1 0 86600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6060
timestamp 1757982896
transform 1 0 88100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6061
timestamp 1757982896
transform 1 0 89600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6062
timestamp 1757982896
transform 1 0 91100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6063
timestamp 1757982896
transform 1 0 92600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6064
timestamp 1757982896
transform 1 0 94100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6065
timestamp 1757982896
transform 1 0 95600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6066
timestamp 1757982896
transform 1 0 97100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6067
timestamp 1757982896
transform 1 0 98600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6068
timestamp 1757982896
transform 1 0 100100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6069
timestamp 1757982896
transform 1 0 101600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6070
timestamp 1757982896
transform 1 0 103100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6071
timestamp 1757982896
transform 1 0 104600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6072
timestamp 1757982896
transform 1 0 106100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6073
timestamp 1757982896
transform 1 0 107600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6074
timestamp 1757982896
transform 1 0 109100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6075
timestamp 1757982896
transform 1 0 110600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6076
timestamp 1757982896
transform 1 0 112100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6077
timestamp 1757982896
transform 1 0 113600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6078
timestamp 1757982896
transform 1 0 115100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6079
timestamp 1757982896
transform 1 0 116600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6080
timestamp 1757982896
transform 1 0 118100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6081
timestamp 1757982896
transform 1 0 119600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6082
timestamp 1757982896
transform 1 0 121100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6083
timestamp 1757982896
transform 1 0 122600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6084
timestamp 1757982896
transform 1 0 124100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6085
timestamp 1757982896
transform 1 0 125600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6086
timestamp 1757982896
transform 1 0 127100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6087
timestamp 1757982896
transform 1 0 128600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6088
timestamp 1757982896
transform 1 0 130100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6089
timestamp 1757982896
transform 1 0 131600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6090
timestamp 1757982896
transform 1 0 133100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6091
timestamp 1757982896
transform 1 0 134600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6092
timestamp 1757982896
transform 1 0 136100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6093
timestamp 1757982896
transform 1 0 137600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6094
timestamp 1757982896
transform 1 0 139100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6095
timestamp 1757982896
transform 1 0 140600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6096
timestamp 1757982896
transform 1 0 142100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6097
timestamp 1757982896
transform 1 0 143600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6098
timestamp 1757982896
transform 1 0 145100 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6099
timestamp 1757982896
transform 1 0 146600 0 1 -88650
box 1820 -1430 3480 230
use pixel  pixel_6100
timestamp 1757982896
transform 1 0 -1900 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6101
timestamp 1757982896
transform 1 0 -400 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6102
timestamp 1757982896
transform 1 0 1100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6103
timestamp 1757982896
transform 1 0 2600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6104
timestamp 1757982896
transform 1 0 4100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6105
timestamp 1757982896
transform 1 0 5600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6106
timestamp 1757982896
transform 1 0 7100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6107
timestamp 1757982896
transform 1 0 8600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6108
timestamp 1757982896
transform 1 0 10100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6109
timestamp 1757982896
transform 1 0 11600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6110
timestamp 1757982896
transform 1 0 13100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6111
timestamp 1757982896
transform 1 0 14600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6112
timestamp 1757982896
transform 1 0 16100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6113
timestamp 1757982896
transform 1 0 17600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6114
timestamp 1757982896
transform 1 0 19100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6115
timestamp 1757982896
transform 1 0 20600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6116
timestamp 1757982896
transform 1 0 22100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6117
timestamp 1757982896
transform 1 0 23600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6118
timestamp 1757982896
transform 1 0 25100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6119
timestamp 1757982896
transform 1 0 26600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6120
timestamp 1757982896
transform 1 0 28100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6121
timestamp 1757982896
transform 1 0 29600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6122
timestamp 1757982896
transform 1 0 31100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6123
timestamp 1757982896
transform 1 0 32600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6124
timestamp 1757982896
transform 1 0 34100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6125
timestamp 1757982896
transform 1 0 35600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6126
timestamp 1757982896
transform 1 0 37100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6127
timestamp 1757982896
transform 1 0 38600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6128
timestamp 1757982896
transform 1 0 40100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6129
timestamp 1757982896
transform 1 0 41600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6130
timestamp 1757982896
transform 1 0 43100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6131
timestamp 1757982896
transform 1 0 44600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6132
timestamp 1757982896
transform 1 0 46100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6133
timestamp 1757982896
transform 1 0 47600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6134
timestamp 1757982896
transform 1 0 49100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6135
timestamp 1757982896
transform 1 0 50600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6136
timestamp 1757982896
transform 1 0 52100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6137
timestamp 1757982896
transform 1 0 53600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6138
timestamp 1757982896
transform 1 0 55100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6139
timestamp 1757982896
transform 1 0 56600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6140
timestamp 1757982896
transform 1 0 58100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6141
timestamp 1757982896
transform 1 0 59600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6142
timestamp 1757982896
transform 1 0 61100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6143
timestamp 1757982896
transform 1 0 62600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6144
timestamp 1757982896
transform 1 0 64100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6145
timestamp 1757982896
transform 1 0 65600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6146
timestamp 1757982896
transform 1 0 67100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6147
timestamp 1757982896
transform 1 0 68600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6148
timestamp 1757982896
transform 1 0 70100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6149
timestamp 1757982896
transform 1 0 71600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6150
timestamp 1757982896
transform 1 0 73100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6151
timestamp 1757982896
transform 1 0 74600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6152
timestamp 1757982896
transform 1 0 76100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6153
timestamp 1757982896
transform 1 0 77600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6154
timestamp 1757982896
transform 1 0 79100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6155
timestamp 1757982896
transform 1 0 80600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6156
timestamp 1757982896
transform 1 0 82100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6157
timestamp 1757982896
transform 1 0 83600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6158
timestamp 1757982896
transform 1 0 85100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6159
timestamp 1757982896
transform 1 0 86600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6160
timestamp 1757982896
transform 1 0 88100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6161
timestamp 1757982896
transform 1 0 89600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6162
timestamp 1757982896
transform 1 0 91100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6163
timestamp 1757982896
transform 1 0 92600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6164
timestamp 1757982896
transform 1 0 94100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6165
timestamp 1757982896
transform 1 0 95600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6166
timestamp 1757982896
transform 1 0 97100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6167
timestamp 1757982896
transform 1 0 98600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6168
timestamp 1757982896
transform 1 0 100100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6169
timestamp 1757982896
transform 1 0 101600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6170
timestamp 1757982896
transform 1 0 103100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6171
timestamp 1757982896
transform 1 0 104600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6172
timestamp 1757982896
transform 1 0 106100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6173
timestamp 1757982896
transform 1 0 107600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6174
timestamp 1757982896
transform 1 0 109100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6175
timestamp 1757982896
transform 1 0 110600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6176
timestamp 1757982896
transform 1 0 112100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6177
timestamp 1757982896
transform 1 0 113600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6178
timestamp 1757982896
transform 1 0 115100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6179
timestamp 1757982896
transform 1 0 116600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6180
timestamp 1757982896
transform 1 0 118100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6181
timestamp 1757982896
transform 1 0 119600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6182
timestamp 1757982896
transform 1 0 121100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6183
timestamp 1757982896
transform 1 0 122600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6184
timestamp 1757982896
transform 1 0 124100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6185
timestamp 1757982896
transform 1 0 125600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6186
timestamp 1757982896
transform 1 0 127100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6187
timestamp 1757982896
transform 1 0 128600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6188
timestamp 1757982896
transform 1 0 130100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6189
timestamp 1757982896
transform 1 0 131600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6190
timestamp 1757982896
transform 1 0 133100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6191
timestamp 1757982896
transform 1 0 134600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6192
timestamp 1757982896
transform 1 0 136100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6193
timestamp 1757982896
transform 1 0 137600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6194
timestamp 1757982896
transform 1 0 139100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6195
timestamp 1757982896
transform 1 0 140600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6196
timestamp 1757982896
transform 1 0 142100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6197
timestamp 1757982896
transform 1 0 143600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6198
timestamp 1757982896
transform 1 0 145100 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6199
timestamp 1757982896
transform 1 0 146600 0 1 -90150
box 1820 -1430 3480 230
use pixel  pixel_6200
timestamp 1757982896
transform 1 0 -1900 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6201
timestamp 1757982896
transform 1 0 -400 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6202
timestamp 1757982896
transform 1 0 1100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6203
timestamp 1757982896
transform 1 0 2600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6204
timestamp 1757982896
transform 1 0 4100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6205
timestamp 1757982896
transform 1 0 5600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6206
timestamp 1757982896
transform 1 0 7100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6207
timestamp 1757982896
transform 1 0 8600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6208
timestamp 1757982896
transform 1 0 10100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6209
timestamp 1757982896
transform 1 0 11600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6210
timestamp 1757982896
transform 1 0 13100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6211
timestamp 1757982896
transform 1 0 14600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6212
timestamp 1757982896
transform 1 0 16100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6213
timestamp 1757982896
transform 1 0 17600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6214
timestamp 1757982896
transform 1 0 19100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6215
timestamp 1757982896
transform 1 0 20600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6216
timestamp 1757982896
transform 1 0 22100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6217
timestamp 1757982896
transform 1 0 23600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6218
timestamp 1757982896
transform 1 0 25100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6219
timestamp 1757982896
transform 1 0 26600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6220
timestamp 1757982896
transform 1 0 28100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6221
timestamp 1757982896
transform 1 0 29600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6222
timestamp 1757982896
transform 1 0 31100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6223
timestamp 1757982896
transform 1 0 32600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6224
timestamp 1757982896
transform 1 0 34100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6225
timestamp 1757982896
transform 1 0 35600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6226
timestamp 1757982896
transform 1 0 37100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6227
timestamp 1757982896
transform 1 0 38600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6228
timestamp 1757982896
transform 1 0 40100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6229
timestamp 1757982896
transform 1 0 41600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6230
timestamp 1757982896
transform 1 0 43100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6231
timestamp 1757982896
transform 1 0 44600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6232
timestamp 1757982896
transform 1 0 46100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6233
timestamp 1757982896
transform 1 0 47600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6234
timestamp 1757982896
transform 1 0 49100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6235
timestamp 1757982896
transform 1 0 50600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6236
timestamp 1757982896
transform 1 0 52100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6237
timestamp 1757982896
transform 1 0 53600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6238
timestamp 1757982896
transform 1 0 55100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6239
timestamp 1757982896
transform 1 0 56600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6240
timestamp 1757982896
transform 1 0 58100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6241
timestamp 1757982896
transform 1 0 59600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6242
timestamp 1757982896
transform 1 0 61100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6243
timestamp 1757982896
transform 1 0 62600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6244
timestamp 1757982896
transform 1 0 64100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6245
timestamp 1757982896
transform 1 0 65600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6246
timestamp 1757982896
transform 1 0 67100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6247
timestamp 1757982896
transform 1 0 68600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6248
timestamp 1757982896
transform 1 0 70100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6249
timestamp 1757982896
transform 1 0 71600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6250
timestamp 1757982896
transform 1 0 73100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6251
timestamp 1757982896
transform 1 0 74600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6252
timestamp 1757982896
transform 1 0 76100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6253
timestamp 1757982896
transform 1 0 77600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6254
timestamp 1757982896
transform 1 0 79100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6255
timestamp 1757982896
transform 1 0 80600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6256
timestamp 1757982896
transform 1 0 82100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6257
timestamp 1757982896
transform 1 0 83600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6258
timestamp 1757982896
transform 1 0 85100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6259
timestamp 1757982896
transform 1 0 86600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6260
timestamp 1757982896
transform 1 0 88100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6261
timestamp 1757982896
transform 1 0 89600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6262
timestamp 1757982896
transform 1 0 91100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6263
timestamp 1757982896
transform 1 0 92600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6264
timestamp 1757982896
transform 1 0 94100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6265
timestamp 1757982896
transform 1 0 95600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6266
timestamp 1757982896
transform 1 0 97100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6267
timestamp 1757982896
transform 1 0 98600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6268
timestamp 1757982896
transform 1 0 100100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6269
timestamp 1757982896
transform 1 0 101600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6270
timestamp 1757982896
transform 1 0 103100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6271
timestamp 1757982896
transform 1 0 104600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6272
timestamp 1757982896
transform 1 0 106100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6273
timestamp 1757982896
transform 1 0 107600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6274
timestamp 1757982896
transform 1 0 109100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6275
timestamp 1757982896
transform 1 0 110600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6276
timestamp 1757982896
transform 1 0 112100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6277
timestamp 1757982896
transform 1 0 113600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6278
timestamp 1757982896
transform 1 0 115100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6279
timestamp 1757982896
transform 1 0 116600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6280
timestamp 1757982896
transform 1 0 118100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6281
timestamp 1757982896
transform 1 0 119600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6282
timestamp 1757982896
transform 1 0 121100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6283
timestamp 1757982896
transform 1 0 122600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6284
timestamp 1757982896
transform 1 0 124100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6285
timestamp 1757982896
transform 1 0 125600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6286
timestamp 1757982896
transform 1 0 127100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6287
timestamp 1757982896
transform 1 0 128600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6288
timestamp 1757982896
transform 1 0 130100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6289
timestamp 1757982896
transform 1 0 131600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6290
timestamp 1757982896
transform 1 0 133100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6291
timestamp 1757982896
transform 1 0 134600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6292
timestamp 1757982896
transform 1 0 136100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6293
timestamp 1757982896
transform 1 0 137600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6294
timestamp 1757982896
transform 1 0 139100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6295
timestamp 1757982896
transform 1 0 140600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6296
timestamp 1757982896
transform 1 0 142100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6297
timestamp 1757982896
transform 1 0 143600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6298
timestamp 1757982896
transform 1 0 145100 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6299
timestamp 1757982896
transform 1 0 146600 0 1 -91650
box 1820 -1430 3480 230
use pixel  pixel_6300
timestamp 1757982896
transform 1 0 -1900 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6301
timestamp 1757982896
transform 1 0 -400 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6302
timestamp 1757982896
transform 1 0 1100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6303
timestamp 1757982896
transform 1 0 2600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6304
timestamp 1757982896
transform 1 0 4100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6305
timestamp 1757982896
transform 1 0 5600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6306
timestamp 1757982896
transform 1 0 7100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6307
timestamp 1757982896
transform 1 0 8600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6308
timestamp 1757982896
transform 1 0 10100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6309
timestamp 1757982896
transform 1 0 11600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6310
timestamp 1757982896
transform 1 0 13100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6311
timestamp 1757982896
transform 1 0 14600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6312
timestamp 1757982896
transform 1 0 16100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6313
timestamp 1757982896
transform 1 0 17600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6314
timestamp 1757982896
transform 1 0 19100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6315
timestamp 1757982896
transform 1 0 20600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6316
timestamp 1757982896
transform 1 0 22100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6317
timestamp 1757982896
transform 1 0 23600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6318
timestamp 1757982896
transform 1 0 25100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6319
timestamp 1757982896
transform 1 0 26600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6320
timestamp 1757982896
transform 1 0 28100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6321
timestamp 1757982896
transform 1 0 29600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6322
timestamp 1757982896
transform 1 0 31100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6323
timestamp 1757982896
transform 1 0 32600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6324
timestamp 1757982896
transform 1 0 34100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6325
timestamp 1757982896
transform 1 0 35600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6326
timestamp 1757982896
transform 1 0 37100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6327
timestamp 1757982896
transform 1 0 38600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6328
timestamp 1757982896
transform 1 0 40100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6329
timestamp 1757982896
transform 1 0 41600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6330
timestamp 1757982896
transform 1 0 43100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6331
timestamp 1757982896
transform 1 0 44600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6332
timestamp 1757982896
transform 1 0 46100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6333
timestamp 1757982896
transform 1 0 47600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6334
timestamp 1757982896
transform 1 0 49100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6335
timestamp 1757982896
transform 1 0 50600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6336
timestamp 1757982896
transform 1 0 52100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6337
timestamp 1757982896
transform 1 0 53600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6338
timestamp 1757982896
transform 1 0 55100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6339
timestamp 1757982896
transform 1 0 56600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6340
timestamp 1757982896
transform 1 0 58100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6341
timestamp 1757982896
transform 1 0 59600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6342
timestamp 1757982896
transform 1 0 61100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6343
timestamp 1757982896
transform 1 0 62600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6344
timestamp 1757982896
transform 1 0 64100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6345
timestamp 1757982896
transform 1 0 65600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6346
timestamp 1757982896
transform 1 0 67100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6347
timestamp 1757982896
transform 1 0 68600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6348
timestamp 1757982896
transform 1 0 70100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6349
timestamp 1757982896
transform 1 0 71600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6350
timestamp 1757982896
transform 1 0 73100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6351
timestamp 1757982896
transform 1 0 74600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6352
timestamp 1757982896
transform 1 0 76100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6353
timestamp 1757982896
transform 1 0 77600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6354
timestamp 1757982896
transform 1 0 79100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6355
timestamp 1757982896
transform 1 0 80600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6356
timestamp 1757982896
transform 1 0 82100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6357
timestamp 1757982896
transform 1 0 83600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6358
timestamp 1757982896
transform 1 0 85100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6359
timestamp 1757982896
transform 1 0 86600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6360
timestamp 1757982896
transform 1 0 88100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6361
timestamp 1757982896
transform 1 0 89600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6362
timestamp 1757982896
transform 1 0 91100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6363
timestamp 1757982896
transform 1 0 92600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6364
timestamp 1757982896
transform 1 0 94100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6365
timestamp 1757982896
transform 1 0 95600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6366
timestamp 1757982896
transform 1 0 97100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6367
timestamp 1757982896
transform 1 0 98600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6368
timestamp 1757982896
transform 1 0 100100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6369
timestamp 1757982896
transform 1 0 101600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6370
timestamp 1757982896
transform 1 0 103100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6371
timestamp 1757982896
transform 1 0 104600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6372
timestamp 1757982896
transform 1 0 106100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6373
timestamp 1757982896
transform 1 0 107600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6374
timestamp 1757982896
transform 1 0 109100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6375
timestamp 1757982896
transform 1 0 110600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6376
timestamp 1757982896
transform 1 0 112100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6377
timestamp 1757982896
transform 1 0 113600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6378
timestamp 1757982896
transform 1 0 115100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6379
timestamp 1757982896
transform 1 0 116600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6380
timestamp 1757982896
transform 1 0 118100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6381
timestamp 1757982896
transform 1 0 119600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6382
timestamp 1757982896
transform 1 0 121100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6383
timestamp 1757982896
transform 1 0 122600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6384
timestamp 1757982896
transform 1 0 124100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6385
timestamp 1757982896
transform 1 0 125600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6386
timestamp 1757982896
transform 1 0 127100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6387
timestamp 1757982896
transform 1 0 128600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6388
timestamp 1757982896
transform 1 0 130100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6389
timestamp 1757982896
transform 1 0 131600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6390
timestamp 1757982896
transform 1 0 133100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6391
timestamp 1757982896
transform 1 0 134600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6392
timestamp 1757982896
transform 1 0 136100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6393
timestamp 1757982896
transform 1 0 137600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6394
timestamp 1757982896
transform 1 0 139100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6395
timestamp 1757982896
transform 1 0 140600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6396
timestamp 1757982896
transform 1 0 142100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6397
timestamp 1757982896
transform 1 0 143600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6398
timestamp 1757982896
transform 1 0 145100 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6399
timestamp 1757982896
transform 1 0 146600 0 1 -93150
box 1820 -1430 3480 230
use pixel  pixel_6400
timestamp 1757982896
transform 1 0 -1900 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6401
timestamp 1757982896
transform 1 0 -400 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6402
timestamp 1757982896
transform 1 0 1100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6403
timestamp 1757982896
transform 1 0 2600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6404
timestamp 1757982896
transform 1 0 4100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6405
timestamp 1757982896
transform 1 0 5600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6406
timestamp 1757982896
transform 1 0 7100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6407
timestamp 1757982896
transform 1 0 8600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6408
timestamp 1757982896
transform 1 0 10100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6409
timestamp 1757982896
transform 1 0 11600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6410
timestamp 1757982896
transform 1 0 13100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6411
timestamp 1757982896
transform 1 0 14600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6412
timestamp 1757982896
transform 1 0 16100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6413
timestamp 1757982896
transform 1 0 17600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6414
timestamp 1757982896
transform 1 0 19100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6415
timestamp 1757982896
transform 1 0 20600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6416
timestamp 1757982896
transform 1 0 22100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6417
timestamp 1757982896
transform 1 0 23600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6418
timestamp 1757982896
transform 1 0 25100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6419
timestamp 1757982896
transform 1 0 26600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6420
timestamp 1757982896
transform 1 0 28100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6421
timestamp 1757982896
transform 1 0 29600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6422
timestamp 1757982896
transform 1 0 31100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6423
timestamp 1757982896
transform 1 0 32600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6424
timestamp 1757982896
transform 1 0 34100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6425
timestamp 1757982896
transform 1 0 35600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6426
timestamp 1757982896
transform 1 0 37100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6427
timestamp 1757982896
transform 1 0 38600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6428
timestamp 1757982896
transform 1 0 40100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6429
timestamp 1757982896
transform 1 0 41600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6430
timestamp 1757982896
transform 1 0 43100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6431
timestamp 1757982896
transform 1 0 44600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6432
timestamp 1757982896
transform 1 0 46100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6433
timestamp 1757982896
transform 1 0 47600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6434
timestamp 1757982896
transform 1 0 49100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6435
timestamp 1757982896
transform 1 0 50600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6436
timestamp 1757982896
transform 1 0 52100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6437
timestamp 1757982896
transform 1 0 53600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6438
timestamp 1757982896
transform 1 0 55100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6439
timestamp 1757982896
transform 1 0 56600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6440
timestamp 1757982896
transform 1 0 58100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6441
timestamp 1757982896
transform 1 0 59600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6442
timestamp 1757982896
transform 1 0 61100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6443
timestamp 1757982896
transform 1 0 62600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6444
timestamp 1757982896
transform 1 0 64100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6445
timestamp 1757982896
transform 1 0 65600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6446
timestamp 1757982896
transform 1 0 67100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6447
timestamp 1757982896
transform 1 0 68600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6448
timestamp 1757982896
transform 1 0 70100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6449
timestamp 1757982896
transform 1 0 71600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6450
timestamp 1757982896
transform 1 0 73100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6451
timestamp 1757982896
transform 1 0 74600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6452
timestamp 1757982896
transform 1 0 76100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6453
timestamp 1757982896
transform 1 0 77600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6454
timestamp 1757982896
transform 1 0 79100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6455
timestamp 1757982896
transform 1 0 80600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6456
timestamp 1757982896
transform 1 0 82100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6457
timestamp 1757982896
transform 1 0 83600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6458
timestamp 1757982896
transform 1 0 85100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6459
timestamp 1757982896
transform 1 0 86600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6460
timestamp 1757982896
transform 1 0 88100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6461
timestamp 1757982896
transform 1 0 89600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6462
timestamp 1757982896
transform 1 0 91100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6463
timestamp 1757982896
transform 1 0 92600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6464
timestamp 1757982896
transform 1 0 94100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6465
timestamp 1757982896
transform 1 0 95600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6466
timestamp 1757982896
transform 1 0 97100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6467
timestamp 1757982896
transform 1 0 98600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6468
timestamp 1757982896
transform 1 0 100100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6469
timestamp 1757982896
transform 1 0 101600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6470
timestamp 1757982896
transform 1 0 103100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6471
timestamp 1757982896
transform 1 0 104600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6472
timestamp 1757982896
transform 1 0 106100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6473
timestamp 1757982896
transform 1 0 107600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6474
timestamp 1757982896
transform 1 0 109100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6475
timestamp 1757982896
transform 1 0 110600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6476
timestamp 1757982896
transform 1 0 112100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6477
timestamp 1757982896
transform 1 0 113600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6478
timestamp 1757982896
transform 1 0 115100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6479
timestamp 1757982896
transform 1 0 116600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6480
timestamp 1757982896
transform 1 0 118100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6481
timestamp 1757982896
transform 1 0 119600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6482
timestamp 1757982896
transform 1 0 121100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6483
timestamp 1757982896
transform 1 0 122600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6484
timestamp 1757982896
transform 1 0 124100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6485
timestamp 1757982896
transform 1 0 125600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6486
timestamp 1757982896
transform 1 0 127100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6487
timestamp 1757982896
transform 1 0 128600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6488
timestamp 1757982896
transform 1 0 130100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6489
timestamp 1757982896
transform 1 0 131600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6490
timestamp 1757982896
transform 1 0 133100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6491
timestamp 1757982896
transform 1 0 134600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6492
timestamp 1757982896
transform 1 0 136100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6493
timestamp 1757982896
transform 1 0 137600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6494
timestamp 1757982896
transform 1 0 139100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6495
timestamp 1757982896
transform 1 0 140600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6496
timestamp 1757982896
transform 1 0 142100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6497
timestamp 1757982896
transform 1 0 143600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6498
timestamp 1757982896
transform 1 0 145100 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6499
timestamp 1757982896
transform 1 0 146600 0 1 -94650
box 1820 -1430 3480 230
use pixel  pixel_6500
timestamp 1757982896
transform 1 0 -1900 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6501
timestamp 1757982896
transform 1 0 -400 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6502
timestamp 1757982896
transform 1 0 1100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6503
timestamp 1757982896
transform 1 0 2600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6504
timestamp 1757982896
transform 1 0 4100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6505
timestamp 1757982896
transform 1 0 5600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6506
timestamp 1757982896
transform 1 0 7100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6507
timestamp 1757982896
transform 1 0 8600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6508
timestamp 1757982896
transform 1 0 10100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6509
timestamp 1757982896
transform 1 0 11600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6510
timestamp 1757982896
transform 1 0 13100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6511
timestamp 1757982896
transform 1 0 14600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6512
timestamp 1757982896
transform 1 0 16100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6513
timestamp 1757982896
transform 1 0 17600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6514
timestamp 1757982896
transform 1 0 19100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6515
timestamp 1757982896
transform 1 0 20600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6516
timestamp 1757982896
transform 1 0 22100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6517
timestamp 1757982896
transform 1 0 23600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6518
timestamp 1757982896
transform 1 0 25100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6519
timestamp 1757982896
transform 1 0 26600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6520
timestamp 1757982896
transform 1 0 28100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6521
timestamp 1757982896
transform 1 0 29600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6522
timestamp 1757982896
transform 1 0 31100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6523
timestamp 1757982896
transform 1 0 32600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6524
timestamp 1757982896
transform 1 0 34100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6525
timestamp 1757982896
transform 1 0 35600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6526
timestamp 1757982896
transform 1 0 37100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6527
timestamp 1757982896
transform 1 0 38600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6528
timestamp 1757982896
transform 1 0 40100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6529
timestamp 1757982896
transform 1 0 41600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6530
timestamp 1757982896
transform 1 0 43100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6531
timestamp 1757982896
transform 1 0 44600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6532
timestamp 1757982896
transform 1 0 46100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6533
timestamp 1757982896
transform 1 0 47600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6534
timestamp 1757982896
transform 1 0 49100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6535
timestamp 1757982896
transform 1 0 50600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6536
timestamp 1757982896
transform 1 0 52100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6537
timestamp 1757982896
transform 1 0 53600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6538
timestamp 1757982896
transform 1 0 55100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6539
timestamp 1757982896
transform 1 0 56600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6540
timestamp 1757982896
transform 1 0 58100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6541
timestamp 1757982896
transform 1 0 59600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6542
timestamp 1757982896
transform 1 0 61100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6543
timestamp 1757982896
transform 1 0 62600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6544
timestamp 1757982896
transform 1 0 64100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6545
timestamp 1757982896
transform 1 0 65600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6546
timestamp 1757982896
transform 1 0 67100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6547
timestamp 1757982896
transform 1 0 68600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6548
timestamp 1757982896
transform 1 0 70100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6549
timestamp 1757982896
transform 1 0 71600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6550
timestamp 1757982896
transform 1 0 73100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6551
timestamp 1757982896
transform 1 0 74600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6552
timestamp 1757982896
transform 1 0 76100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6553
timestamp 1757982896
transform 1 0 77600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6554
timestamp 1757982896
transform 1 0 79100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6555
timestamp 1757982896
transform 1 0 80600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6556
timestamp 1757982896
transform 1 0 82100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6557
timestamp 1757982896
transform 1 0 83600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6558
timestamp 1757982896
transform 1 0 85100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6559
timestamp 1757982896
transform 1 0 86600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6560
timestamp 1757982896
transform 1 0 88100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6561
timestamp 1757982896
transform 1 0 89600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6562
timestamp 1757982896
transform 1 0 91100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6563
timestamp 1757982896
transform 1 0 92600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6564
timestamp 1757982896
transform 1 0 94100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6565
timestamp 1757982896
transform 1 0 95600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6566
timestamp 1757982896
transform 1 0 97100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6567
timestamp 1757982896
transform 1 0 98600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6568
timestamp 1757982896
transform 1 0 100100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6569
timestamp 1757982896
transform 1 0 101600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6570
timestamp 1757982896
transform 1 0 103100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6571
timestamp 1757982896
transform 1 0 104600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6572
timestamp 1757982896
transform 1 0 106100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6573
timestamp 1757982896
transform 1 0 107600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6574
timestamp 1757982896
transform 1 0 109100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6575
timestamp 1757982896
transform 1 0 110600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6576
timestamp 1757982896
transform 1 0 112100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6577
timestamp 1757982896
transform 1 0 113600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6578
timestamp 1757982896
transform 1 0 115100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6579
timestamp 1757982896
transform 1 0 116600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6580
timestamp 1757982896
transform 1 0 118100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6581
timestamp 1757982896
transform 1 0 119600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6582
timestamp 1757982896
transform 1 0 121100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6583
timestamp 1757982896
transform 1 0 122600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6584
timestamp 1757982896
transform 1 0 124100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6585
timestamp 1757982896
transform 1 0 125600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6586
timestamp 1757982896
transform 1 0 127100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6587
timestamp 1757982896
transform 1 0 128600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6588
timestamp 1757982896
transform 1 0 130100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6589
timestamp 1757982896
transform 1 0 131600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6590
timestamp 1757982896
transform 1 0 133100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6591
timestamp 1757982896
transform 1 0 134600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6592
timestamp 1757982896
transform 1 0 136100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6593
timestamp 1757982896
transform 1 0 137600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6594
timestamp 1757982896
transform 1 0 139100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6595
timestamp 1757982896
transform 1 0 140600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6596
timestamp 1757982896
transform 1 0 142100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6597
timestamp 1757982896
transform 1 0 143600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6598
timestamp 1757982896
transform 1 0 145100 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6599
timestamp 1757982896
transform 1 0 146600 0 1 -96150
box 1820 -1430 3480 230
use pixel  pixel_6600
timestamp 1757982896
transform 1 0 -1900 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6601
timestamp 1757982896
transform 1 0 -400 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6602
timestamp 1757982896
transform 1 0 1100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6603
timestamp 1757982896
transform 1 0 2600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6604
timestamp 1757982896
transform 1 0 4100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6605
timestamp 1757982896
transform 1 0 5600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6606
timestamp 1757982896
transform 1 0 7100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6607
timestamp 1757982896
transform 1 0 8600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6608
timestamp 1757982896
transform 1 0 10100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6609
timestamp 1757982896
transform 1 0 11600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6610
timestamp 1757982896
transform 1 0 13100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6611
timestamp 1757982896
transform 1 0 14600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6612
timestamp 1757982896
transform 1 0 16100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6613
timestamp 1757982896
transform 1 0 17600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6614
timestamp 1757982896
transform 1 0 19100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6615
timestamp 1757982896
transform 1 0 20600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6616
timestamp 1757982896
transform 1 0 22100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6617
timestamp 1757982896
transform 1 0 23600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6618
timestamp 1757982896
transform 1 0 25100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6619
timestamp 1757982896
transform 1 0 26600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6620
timestamp 1757982896
transform 1 0 28100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6621
timestamp 1757982896
transform 1 0 29600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6622
timestamp 1757982896
transform 1 0 31100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6623
timestamp 1757982896
transform 1 0 32600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6624
timestamp 1757982896
transform 1 0 34100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6625
timestamp 1757982896
transform 1 0 35600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6626
timestamp 1757982896
transform 1 0 37100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6627
timestamp 1757982896
transform 1 0 38600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6628
timestamp 1757982896
transform 1 0 40100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6629
timestamp 1757982896
transform 1 0 41600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6630
timestamp 1757982896
transform 1 0 43100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6631
timestamp 1757982896
transform 1 0 44600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6632
timestamp 1757982896
transform 1 0 46100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6633
timestamp 1757982896
transform 1 0 47600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6634
timestamp 1757982896
transform 1 0 49100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6635
timestamp 1757982896
transform 1 0 50600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6636
timestamp 1757982896
transform 1 0 52100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6637
timestamp 1757982896
transform 1 0 53600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6638
timestamp 1757982896
transform 1 0 55100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6639
timestamp 1757982896
transform 1 0 56600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6640
timestamp 1757982896
transform 1 0 58100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6641
timestamp 1757982896
transform 1 0 59600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6642
timestamp 1757982896
transform 1 0 61100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6643
timestamp 1757982896
transform 1 0 62600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6644
timestamp 1757982896
transform 1 0 64100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6645
timestamp 1757982896
transform 1 0 65600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6646
timestamp 1757982896
transform 1 0 67100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6647
timestamp 1757982896
transform 1 0 68600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6648
timestamp 1757982896
transform 1 0 70100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6649
timestamp 1757982896
transform 1 0 71600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6650
timestamp 1757982896
transform 1 0 73100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6651
timestamp 1757982896
transform 1 0 74600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6652
timestamp 1757982896
transform 1 0 76100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6653
timestamp 1757982896
transform 1 0 77600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6654
timestamp 1757982896
transform 1 0 79100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6655
timestamp 1757982896
transform 1 0 80600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6656
timestamp 1757982896
transform 1 0 82100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6657
timestamp 1757982896
transform 1 0 83600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6658
timestamp 1757982896
transform 1 0 85100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6659
timestamp 1757982896
transform 1 0 86600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6660
timestamp 1757982896
transform 1 0 88100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6661
timestamp 1757982896
transform 1 0 89600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6662
timestamp 1757982896
transform 1 0 91100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6663
timestamp 1757982896
transform 1 0 92600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6664
timestamp 1757982896
transform 1 0 94100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6665
timestamp 1757982896
transform 1 0 95600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6666
timestamp 1757982896
transform 1 0 97100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6667
timestamp 1757982896
transform 1 0 98600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6668
timestamp 1757982896
transform 1 0 100100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6669
timestamp 1757982896
transform 1 0 101600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6670
timestamp 1757982896
transform 1 0 103100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6671
timestamp 1757982896
transform 1 0 104600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6672
timestamp 1757982896
transform 1 0 106100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6673
timestamp 1757982896
transform 1 0 107600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6674
timestamp 1757982896
transform 1 0 109100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6675
timestamp 1757982896
transform 1 0 110600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6676
timestamp 1757982896
transform 1 0 112100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6677
timestamp 1757982896
transform 1 0 113600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6678
timestamp 1757982896
transform 1 0 115100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6679
timestamp 1757982896
transform 1 0 116600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6680
timestamp 1757982896
transform 1 0 118100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6681
timestamp 1757982896
transform 1 0 119600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6682
timestamp 1757982896
transform 1 0 121100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6683
timestamp 1757982896
transform 1 0 122600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6684
timestamp 1757982896
transform 1 0 124100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6685
timestamp 1757982896
transform 1 0 125600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6686
timestamp 1757982896
transform 1 0 127100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6687
timestamp 1757982896
transform 1 0 128600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6688
timestamp 1757982896
transform 1 0 130100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6689
timestamp 1757982896
transform 1 0 131600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6690
timestamp 1757982896
transform 1 0 133100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6691
timestamp 1757982896
transform 1 0 134600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6692
timestamp 1757982896
transform 1 0 136100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6693
timestamp 1757982896
transform 1 0 137600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6694
timestamp 1757982896
transform 1 0 139100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6695
timestamp 1757982896
transform 1 0 140600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6696
timestamp 1757982896
transform 1 0 142100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6697
timestamp 1757982896
transform 1 0 143600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6698
timestamp 1757982896
transform 1 0 145100 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6699
timestamp 1757982896
transform 1 0 146600 0 1 -97650
box 1820 -1430 3480 230
use pixel  pixel_6700
timestamp 1757982896
transform 1 0 -1900 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6701
timestamp 1757982896
transform 1 0 -400 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6702
timestamp 1757982896
transform 1 0 1100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6703
timestamp 1757982896
transform 1 0 2600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6704
timestamp 1757982896
transform 1 0 4100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6705
timestamp 1757982896
transform 1 0 5600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6706
timestamp 1757982896
transform 1 0 7100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6707
timestamp 1757982896
transform 1 0 8600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6708
timestamp 1757982896
transform 1 0 10100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6709
timestamp 1757982896
transform 1 0 11600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6710
timestamp 1757982896
transform 1 0 13100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6711
timestamp 1757982896
transform 1 0 14600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6712
timestamp 1757982896
transform 1 0 16100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6713
timestamp 1757982896
transform 1 0 17600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6714
timestamp 1757982896
transform 1 0 19100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6715
timestamp 1757982896
transform 1 0 20600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6716
timestamp 1757982896
transform 1 0 22100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6717
timestamp 1757982896
transform 1 0 23600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6718
timestamp 1757982896
transform 1 0 25100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6719
timestamp 1757982896
transform 1 0 26600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6720
timestamp 1757982896
transform 1 0 28100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6721
timestamp 1757982896
transform 1 0 29600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6722
timestamp 1757982896
transform 1 0 31100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6723
timestamp 1757982896
transform 1 0 32600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6724
timestamp 1757982896
transform 1 0 34100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6725
timestamp 1757982896
transform 1 0 35600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6726
timestamp 1757982896
transform 1 0 37100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6727
timestamp 1757982896
transform 1 0 38600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6728
timestamp 1757982896
transform 1 0 40100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6729
timestamp 1757982896
transform 1 0 41600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6730
timestamp 1757982896
transform 1 0 43100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6731
timestamp 1757982896
transform 1 0 44600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6732
timestamp 1757982896
transform 1 0 46100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6733
timestamp 1757982896
transform 1 0 47600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6734
timestamp 1757982896
transform 1 0 49100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6735
timestamp 1757982896
transform 1 0 50600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6736
timestamp 1757982896
transform 1 0 52100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6737
timestamp 1757982896
transform 1 0 53600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6738
timestamp 1757982896
transform 1 0 55100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6739
timestamp 1757982896
transform 1 0 56600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6740
timestamp 1757982896
transform 1 0 58100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6741
timestamp 1757982896
transform 1 0 59600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6742
timestamp 1757982896
transform 1 0 61100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6743
timestamp 1757982896
transform 1 0 62600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6744
timestamp 1757982896
transform 1 0 64100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6745
timestamp 1757982896
transform 1 0 65600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6746
timestamp 1757982896
transform 1 0 67100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6747
timestamp 1757982896
transform 1 0 68600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6748
timestamp 1757982896
transform 1 0 70100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6749
timestamp 1757982896
transform 1 0 71600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6750
timestamp 1757982896
transform 1 0 73100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6751
timestamp 1757982896
transform 1 0 74600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6752
timestamp 1757982896
transform 1 0 76100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6753
timestamp 1757982896
transform 1 0 77600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6754
timestamp 1757982896
transform 1 0 79100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6755
timestamp 1757982896
transform 1 0 80600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6756
timestamp 1757982896
transform 1 0 82100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6757
timestamp 1757982896
transform 1 0 83600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6758
timestamp 1757982896
transform 1 0 85100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6759
timestamp 1757982896
transform 1 0 86600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6760
timestamp 1757982896
transform 1 0 88100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6761
timestamp 1757982896
transform 1 0 89600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6762
timestamp 1757982896
transform 1 0 91100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6763
timestamp 1757982896
transform 1 0 92600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6764
timestamp 1757982896
transform 1 0 94100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6765
timestamp 1757982896
transform 1 0 95600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6766
timestamp 1757982896
transform 1 0 97100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6767
timestamp 1757982896
transform 1 0 98600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6768
timestamp 1757982896
transform 1 0 100100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6769
timestamp 1757982896
transform 1 0 101600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6770
timestamp 1757982896
transform 1 0 103100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6771
timestamp 1757982896
transform 1 0 104600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6772
timestamp 1757982896
transform 1 0 106100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6773
timestamp 1757982896
transform 1 0 107600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6774
timestamp 1757982896
transform 1 0 109100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6775
timestamp 1757982896
transform 1 0 110600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6776
timestamp 1757982896
transform 1 0 112100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6777
timestamp 1757982896
transform 1 0 113600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6778
timestamp 1757982896
transform 1 0 115100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6779
timestamp 1757982896
transform 1 0 116600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6780
timestamp 1757982896
transform 1 0 118100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6781
timestamp 1757982896
transform 1 0 119600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6782
timestamp 1757982896
transform 1 0 121100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6783
timestamp 1757982896
transform 1 0 122600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6784
timestamp 1757982896
transform 1 0 124100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6785
timestamp 1757982896
transform 1 0 125600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6786
timestamp 1757982896
transform 1 0 127100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6787
timestamp 1757982896
transform 1 0 128600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6788
timestamp 1757982896
transform 1 0 130100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6789
timestamp 1757982896
transform 1 0 131600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6790
timestamp 1757982896
transform 1 0 133100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6791
timestamp 1757982896
transform 1 0 134600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6792
timestamp 1757982896
transform 1 0 136100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6793
timestamp 1757982896
transform 1 0 137600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6794
timestamp 1757982896
transform 1 0 139100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6795
timestamp 1757982896
transform 1 0 140600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6796
timestamp 1757982896
transform 1 0 142100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6797
timestamp 1757982896
transform 1 0 143600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6798
timestamp 1757982896
transform 1 0 145100 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6799
timestamp 1757982896
transform 1 0 146600 0 1 -99150
box 1820 -1430 3480 230
use pixel  pixel_6800
timestamp 1757982896
transform 1 0 -1900 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6801
timestamp 1757982896
transform 1 0 -400 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6802
timestamp 1757982896
transform 1 0 1100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6803
timestamp 1757982896
transform 1 0 2600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6804
timestamp 1757982896
transform 1 0 4100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6805
timestamp 1757982896
transform 1 0 5600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6806
timestamp 1757982896
transform 1 0 7100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6807
timestamp 1757982896
transform 1 0 8600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6808
timestamp 1757982896
transform 1 0 10100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6809
timestamp 1757982896
transform 1 0 11600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6810
timestamp 1757982896
transform 1 0 13100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6811
timestamp 1757982896
transform 1 0 14600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6812
timestamp 1757982896
transform 1 0 16100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6813
timestamp 1757982896
transform 1 0 17600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6814
timestamp 1757982896
transform 1 0 19100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6815
timestamp 1757982896
transform 1 0 20600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6816
timestamp 1757982896
transform 1 0 22100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6817
timestamp 1757982896
transform 1 0 23600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6818
timestamp 1757982896
transform 1 0 25100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6819
timestamp 1757982896
transform 1 0 26600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6820
timestamp 1757982896
transform 1 0 28100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6821
timestamp 1757982896
transform 1 0 29600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6822
timestamp 1757982896
transform 1 0 31100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6823
timestamp 1757982896
transform 1 0 32600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6824
timestamp 1757982896
transform 1 0 34100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6825
timestamp 1757982896
transform 1 0 35600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6826
timestamp 1757982896
transform 1 0 37100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6827
timestamp 1757982896
transform 1 0 38600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6828
timestamp 1757982896
transform 1 0 40100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6829
timestamp 1757982896
transform 1 0 41600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6830
timestamp 1757982896
transform 1 0 43100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6831
timestamp 1757982896
transform 1 0 44600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6832
timestamp 1757982896
transform 1 0 46100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6833
timestamp 1757982896
transform 1 0 47600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6834
timestamp 1757982896
transform 1 0 49100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6835
timestamp 1757982896
transform 1 0 50600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6836
timestamp 1757982896
transform 1 0 52100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6837
timestamp 1757982896
transform 1 0 53600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6838
timestamp 1757982896
transform 1 0 55100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6839
timestamp 1757982896
transform 1 0 56600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6840
timestamp 1757982896
transform 1 0 58100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6841
timestamp 1757982896
transform 1 0 59600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6842
timestamp 1757982896
transform 1 0 61100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6843
timestamp 1757982896
transform 1 0 62600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6844
timestamp 1757982896
transform 1 0 64100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6845
timestamp 1757982896
transform 1 0 65600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6846
timestamp 1757982896
transform 1 0 67100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6847
timestamp 1757982896
transform 1 0 68600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6848
timestamp 1757982896
transform 1 0 70100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6849
timestamp 1757982896
transform 1 0 71600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6850
timestamp 1757982896
transform 1 0 73100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6851
timestamp 1757982896
transform 1 0 74600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6852
timestamp 1757982896
transform 1 0 76100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6853
timestamp 1757982896
transform 1 0 77600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6854
timestamp 1757982896
transform 1 0 79100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6855
timestamp 1757982896
transform 1 0 80600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6856
timestamp 1757982896
transform 1 0 82100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6857
timestamp 1757982896
transform 1 0 83600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6858
timestamp 1757982896
transform 1 0 85100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6859
timestamp 1757982896
transform 1 0 86600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6860
timestamp 1757982896
transform 1 0 88100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6861
timestamp 1757982896
transform 1 0 89600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6862
timestamp 1757982896
transform 1 0 91100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6863
timestamp 1757982896
transform 1 0 92600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6864
timestamp 1757982896
transform 1 0 94100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6865
timestamp 1757982896
transform 1 0 95600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6866
timestamp 1757982896
transform 1 0 97100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6867
timestamp 1757982896
transform 1 0 98600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6868
timestamp 1757982896
transform 1 0 100100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6869
timestamp 1757982896
transform 1 0 101600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6870
timestamp 1757982896
transform 1 0 103100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6871
timestamp 1757982896
transform 1 0 104600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6872
timestamp 1757982896
transform 1 0 106100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6873
timestamp 1757982896
transform 1 0 107600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6874
timestamp 1757982896
transform 1 0 109100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6875
timestamp 1757982896
transform 1 0 110600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6876
timestamp 1757982896
transform 1 0 112100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6877
timestamp 1757982896
transform 1 0 113600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6878
timestamp 1757982896
transform 1 0 115100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6879
timestamp 1757982896
transform 1 0 116600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6880
timestamp 1757982896
transform 1 0 118100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6881
timestamp 1757982896
transform 1 0 119600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6882
timestamp 1757982896
transform 1 0 121100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6883
timestamp 1757982896
transform 1 0 122600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6884
timestamp 1757982896
transform 1 0 124100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6885
timestamp 1757982896
transform 1 0 125600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6886
timestamp 1757982896
transform 1 0 127100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6887
timestamp 1757982896
transform 1 0 128600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6888
timestamp 1757982896
transform 1 0 130100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6889
timestamp 1757982896
transform 1 0 131600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6890
timestamp 1757982896
transform 1 0 133100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6891
timestamp 1757982896
transform 1 0 134600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6892
timestamp 1757982896
transform 1 0 136100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6893
timestamp 1757982896
transform 1 0 137600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6894
timestamp 1757982896
transform 1 0 139100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6895
timestamp 1757982896
transform 1 0 140600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6896
timestamp 1757982896
transform 1 0 142100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6897
timestamp 1757982896
transform 1 0 143600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6898
timestamp 1757982896
transform 1 0 145100 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6899
timestamp 1757982896
transform 1 0 146600 0 1 -100650
box 1820 -1430 3480 230
use pixel  pixel_6900
timestamp 1757982896
transform 1 0 -1900 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6901
timestamp 1757982896
transform 1 0 -400 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6902
timestamp 1757982896
transform 1 0 1100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6903
timestamp 1757982896
transform 1 0 2600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6904
timestamp 1757982896
transform 1 0 4100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6905
timestamp 1757982896
transform 1 0 5600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6906
timestamp 1757982896
transform 1 0 7100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6907
timestamp 1757982896
transform 1 0 8600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6908
timestamp 1757982896
transform 1 0 10100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6909
timestamp 1757982896
transform 1 0 11600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6910
timestamp 1757982896
transform 1 0 13100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6911
timestamp 1757982896
transform 1 0 14600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6912
timestamp 1757982896
transform 1 0 16100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6913
timestamp 1757982896
transform 1 0 17600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6914
timestamp 1757982896
transform 1 0 19100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6915
timestamp 1757982896
transform 1 0 20600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6916
timestamp 1757982896
transform 1 0 22100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6917
timestamp 1757982896
transform 1 0 23600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6918
timestamp 1757982896
transform 1 0 25100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6919
timestamp 1757982896
transform 1 0 26600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6920
timestamp 1757982896
transform 1 0 28100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6921
timestamp 1757982896
transform 1 0 29600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6922
timestamp 1757982896
transform 1 0 31100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6923
timestamp 1757982896
transform 1 0 32600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6924
timestamp 1757982896
transform 1 0 34100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6925
timestamp 1757982896
transform 1 0 35600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6926
timestamp 1757982896
transform 1 0 37100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6927
timestamp 1757982896
transform 1 0 38600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6928
timestamp 1757982896
transform 1 0 40100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6929
timestamp 1757982896
transform 1 0 41600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6930
timestamp 1757982896
transform 1 0 43100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6931
timestamp 1757982896
transform 1 0 44600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6932
timestamp 1757982896
transform 1 0 46100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6933
timestamp 1757982896
transform 1 0 47600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6934
timestamp 1757982896
transform 1 0 49100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6935
timestamp 1757982896
transform 1 0 50600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6936
timestamp 1757982896
transform 1 0 52100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6937
timestamp 1757982896
transform 1 0 53600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6938
timestamp 1757982896
transform 1 0 55100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6939
timestamp 1757982896
transform 1 0 56600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6940
timestamp 1757982896
transform 1 0 58100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6941
timestamp 1757982896
transform 1 0 59600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6942
timestamp 1757982896
transform 1 0 61100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6943
timestamp 1757982896
transform 1 0 62600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6944
timestamp 1757982896
transform 1 0 64100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6945
timestamp 1757982896
transform 1 0 65600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6946
timestamp 1757982896
transform 1 0 67100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6947
timestamp 1757982896
transform 1 0 68600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6948
timestamp 1757982896
transform 1 0 70100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6949
timestamp 1757982896
transform 1 0 71600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6950
timestamp 1757982896
transform 1 0 73100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6951
timestamp 1757982896
transform 1 0 74600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6952
timestamp 1757982896
transform 1 0 76100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6953
timestamp 1757982896
transform 1 0 77600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6954
timestamp 1757982896
transform 1 0 79100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6955
timestamp 1757982896
transform 1 0 80600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6956
timestamp 1757982896
transform 1 0 82100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6957
timestamp 1757982896
transform 1 0 83600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6958
timestamp 1757982896
transform 1 0 85100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6959
timestamp 1757982896
transform 1 0 86600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6960
timestamp 1757982896
transform 1 0 88100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6961
timestamp 1757982896
transform 1 0 89600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6962
timestamp 1757982896
transform 1 0 91100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6963
timestamp 1757982896
transform 1 0 92600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6964
timestamp 1757982896
transform 1 0 94100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6965
timestamp 1757982896
transform 1 0 95600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6966
timestamp 1757982896
transform 1 0 97100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6967
timestamp 1757982896
transform 1 0 98600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6968
timestamp 1757982896
transform 1 0 100100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6969
timestamp 1757982896
transform 1 0 101600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6970
timestamp 1757982896
transform 1 0 103100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6971
timestamp 1757982896
transform 1 0 104600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6972
timestamp 1757982896
transform 1 0 106100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6973
timestamp 1757982896
transform 1 0 107600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6974
timestamp 1757982896
transform 1 0 109100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6975
timestamp 1757982896
transform 1 0 110600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6976
timestamp 1757982896
transform 1 0 112100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6977
timestamp 1757982896
transform 1 0 113600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6978
timestamp 1757982896
transform 1 0 115100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6979
timestamp 1757982896
transform 1 0 116600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6980
timestamp 1757982896
transform 1 0 118100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6981
timestamp 1757982896
transform 1 0 119600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6982
timestamp 1757982896
transform 1 0 121100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6983
timestamp 1757982896
transform 1 0 122600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6984
timestamp 1757982896
transform 1 0 124100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6985
timestamp 1757982896
transform 1 0 125600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6986
timestamp 1757982896
transform 1 0 127100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6987
timestamp 1757982896
transform 1 0 128600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6988
timestamp 1757982896
transform 1 0 130100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6989
timestamp 1757982896
transform 1 0 131600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6990
timestamp 1757982896
transform 1 0 133100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6991
timestamp 1757982896
transform 1 0 134600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6992
timestamp 1757982896
transform 1 0 136100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6993
timestamp 1757982896
transform 1 0 137600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6994
timestamp 1757982896
transform 1 0 139100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6995
timestamp 1757982896
transform 1 0 140600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6996
timestamp 1757982896
transform 1 0 142100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6997
timestamp 1757982896
transform 1 0 143600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6998
timestamp 1757982896
transform 1 0 145100 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_6999
timestamp 1757982896
transform 1 0 146600 0 1 -102150
box 1820 -1430 3480 230
use pixel  pixel_7000
timestamp 1757982896
transform 1 0 -1900 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7001
timestamp 1757982896
transform 1 0 -400 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7002
timestamp 1757982896
transform 1 0 1100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7003
timestamp 1757982896
transform 1 0 2600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7004
timestamp 1757982896
transform 1 0 4100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7005
timestamp 1757982896
transform 1 0 5600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7006
timestamp 1757982896
transform 1 0 7100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7007
timestamp 1757982896
transform 1 0 8600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7008
timestamp 1757982896
transform 1 0 10100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7009
timestamp 1757982896
transform 1 0 11600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7010
timestamp 1757982896
transform 1 0 13100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7011
timestamp 1757982896
transform 1 0 14600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7012
timestamp 1757982896
transform 1 0 16100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7013
timestamp 1757982896
transform 1 0 17600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7014
timestamp 1757982896
transform 1 0 19100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7015
timestamp 1757982896
transform 1 0 20600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7016
timestamp 1757982896
transform 1 0 22100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7017
timestamp 1757982896
transform 1 0 23600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7018
timestamp 1757982896
transform 1 0 25100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7019
timestamp 1757982896
transform 1 0 26600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7020
timestamp 1757982896
transform 1 0 28100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7021
timestamp 1757982896
transform 1 0 29600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7022
timestamp 1757982896
transform 1 0 31100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7023
timestamp 1757982896
transform 1 0 32600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7024
timestamp 1757982896
transform 1 0 34100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7025
timestamp 1757982896
transform 1 0 35600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7026
timestamp 1757982896
transform 1 0 37100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7027
timestamp 1757982896
transform 1 0 38600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7028
timestamp 1757982896
transform 1 0 40100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7029
timestamp 1757982896
transform 1 0 41600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7030
timestamp 1757982896
transform 1 0 43100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7031
timestamp 1757982896
transform 1 0 44600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7032
timestamp 1757982896
transform 1 0 46100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7033
timestamp 1757982896
transform 1 0 47600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7034
timestamp 1757982896
transform 1 0 49100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7035
timestamp 1757982896
transform 1 0 50600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7036
timestamp 1757982896
transform 1 0 52100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7037
timestamp 1757982896
transform 1 0 53600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7038
timestamp 1757982896
transform 1 0 55100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7039
timestamp 1757982896
transform 1 0 56600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7040
timestamp 1757982896
transform 1 0 58100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7041
timestamp 1757982896
transform 1 0 59600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7042
timestamp 1757982896
transform 1 0 61100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7043
timestamp 1757982896
transform 1 0 62600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7044
timestamp 1757982896
transform 1 0 64100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7045
timestamp 1757982896
transform 1 0 65600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7046
timestamp 1757982896
transform 1 0 67100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7047
timestamp 1757982896
transform 1 0 68600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7048
timestamp 1757982896
transform 1 0 70100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7049
timestamp 1757982896
transform 1 0 71600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7050
timestamp 1757982896
transform 1 0 73100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7051
timestamp 1757982896
transform 1 0 74600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7052
timestamp 1757982896
transform 1 0 76100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7053
timestamp 1757982896
transform 1 0 77600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7054
timestamp 1757982896
transform 1 0 79100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7055
timestamp 1757982896
transform 1 0 80600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7056
timestamp 1757982896
transform 1 0 82100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7057
timestamp 1757982896
transform 1 0 83600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7058
timestamp 1757982896
transform 1 0 85100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7059
timestamp 1757982896
transform 1 0 86600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7060
timestamp 1757982896
transform 1 0 88100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7061
timestamp 1757982896
transform 1 0 89600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7062
timestamp 1757982896
transform 1 0 91100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7063
timestamp 1757982896
transform 1 0 92600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7064
timestamp 1757982896
transform 1 0 94100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7065
timestamp 1757982896
transform 1 0 95600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7066
timestamp 1757982896
transform 1 0 97100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7067
timestamp 1757982896
transform 1 0 98600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7068
timestamp 1757982896
transform 1 0 100100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7069
timestamp 1757982896
transform 1 0 101600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7070
timestamp 1757982896
transform 1 0 103100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7071
timestamp 1757982896
transform 1 0 104600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7072
timestamp 1757982896
transform 1 0 106100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7073
timestamp 1757982896
transform 1 0 107600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7074
timestamp 1757982896
transform 1 0 109100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7075
timestamp 1757982896
transform 1 0 110600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7076
timestamp 1757982896
transform 1 0 112100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7077
timestamp 1757982896
transform 1 0 113600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7078
timestamp 1757982896
transform 1 0 115100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7079
timestamp 1757982896
transform 1 0 116600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7080
timestamp 1757982896
transform 1 0 118100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7081
timestamp 1757982896
transform 1 0 119600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7082
timestamp 1757982896
transform 1 0 121100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7083
timestamp 1757982896
transform 1 0 122600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7084
timestamp 1757982896
transform 1 0 124100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7085
timestamp 1757982896
transform 1 0 125600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7086
timestamp 1757982896
transform 1 0 127100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7087
timestamp 1757982896
transform 1 0 128600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7088
timestamp 1757982896
transform 1 0 130100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7089
timestamp 1757982896
transform 1 0 131600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7090
timestamp 1757982896
transform 1 0 133100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7091
timestamp 1757982896
transform 1 0 134600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7092
timestamp 1757982896
transform 1 0 136100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7093
timestamp 1757982896
transform 1 0 137600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7094
timestamp 1757982896
transform 1 0 139100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7095
timestamp 1757982896
transform 1 0 140600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7096
timestamp 1757982896
transform 1 0 142100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7097
timestamp 1757982896
transform 1 0 143600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7098
timestamp 1757982896
transform 1 0 145100 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7099
timestamp 1757982896
transform 1 0 146600 0 1 -103650
box 1820 -1430 3480 230
use pixel  pixel_7100
timestamp 1757982896
transform 1 0 -1900 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7101
timestamp 1757982896
transform 1 0 -400 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7102
timestamp 1757982896
transform 1 0 1100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7103
timestamp 1757982896
transform 1 0 2600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7104
timestamp 1757982896
transform 1 0 4100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7105
timestamp 1757982896
transform 1 0 5600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7106
timestamp 1757982896
transform 1 0 7100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7107
timestamp 1757982896
transform 1 0 8600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7108
timestamp 1757982896
transform 1 0 10100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7109
timestamp 1757982896
transform 1 0 11600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7110
timestamp 1757982896
transform 1 0 13100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7111
timestamp 1757982896
transform 1 0 14600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7112
timestamp 1757982896
transform 1 0 16100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7113
timestamp 1757982896
transform 1 0 17600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7114
timestamp 1757982896
transform 1 0 19100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7115
timestamp 1757982896
transform 1 0 20600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7116
timestamp 1757982896
transform 1 0 22100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7117
timestamp 1757982896
transform 1 0 23600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7118
timestamp 1757982896
transform 1 0 25100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7119
timestamp 1757982896
transform 1 0 26600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7120
timestamp 1757982896
transform 1 0 28100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7121
timestamp 1757982896
transform 1 0 29600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7122
timestamp 1757982896
transform 1 0 31100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7123
timestamp 1757982896
transform 1 0 32600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7124
timestamp 1757982896
transform 1 0 34100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7125
timestamp 1757982896
transform 1 0 35600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7126
timestamp 1757982896
transform 1 0 37100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7127
timestamp 1757982896
transform 1 0 38600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7128
timestamp 1757982896
transform 1 0 40100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7129
timestamp 1757982896
transform 1 0 41600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7130
timestamp 1757982896
transform 1 0 43100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7131
timestamp 1757982896
transform 1 0 44600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7132
timestamp 1757982896
transform 1 0 46100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7133
timestamp 1757982896
transform 1 0 47600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7134
timestamp 1757982896
transform 1 0 49100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7135
timestamp 1757982896
transform 1 0 50600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7136
timestamp 1757982896
transform 1 0 52100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7137
timestamp 1757982896
transform 1 0 53600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7138
timestamp 1757982896
transform 1 0 55100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7139
timestamp 1757982896
transform 1 0 56600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7140
timestamp 1757982896
transform 1 0 58100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7141
timestamp 1757982896
transform 1 0 59600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7142
timestamp 1757982896
transform 1 0 61100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7143
timestamp 1757982896
transform 1 0 62600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7144
timestamp 1757982896
transform 1 0 64100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7145
timestamp 1757982896
transform 1 0 65600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7146
timestamp 1757982896
transform 1 0 67100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7147
timestamp 1757982896
transform 1 0 68600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7148
timestamp 1757982896
transform 1 0 70100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7149
timestamp 1757982896
transform 1 0 71600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7150
timestamp 1757982896
transform 1 0 73100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7151
timestamp 1757982896
transform 1 0 74600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7152
timestamp 1757982896
transform 1 0 76100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7153
timestamp 1757982896
transform 1 0 77600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7154
timestamp 1757982896
transform 1 0 79100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7155
timestamp 1757982896
transform 1 0 80600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7156
timestamp 1757982896
transform 1 0 82100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7157
timestamp 1757982896
transform 1 0 83600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7158
timestamp 1757982896
transform 1 0 85100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7159
timestamp 1757982896
transform 1 0 86600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7160
timestamp 1757982896
transform 1 0 88100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7161
timestamp 1757982896
transform 1 0 89600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7162
timestamp 1757982896
transform 1 0 91100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7163
timestamp 1757982896
transform 1 0 92600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7164
timestamp 1757982896
transform 1 0 94100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7165
timestamp 1757982896
transform 1 0 95600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7166
timestamp 1757982896
transform 1 0 97100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7167
timestamp 1757982896
transform 1 0 98600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7168
timestamp 1757982896
transform 1 0 100100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7169
timestamp 1757982896
transform 1 0 101600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7170
timestamp 1757982896
transform 1 0 103100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7171
timestamp 1757982896
transform 1 0 104600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7172
timestamp 1757982896
transform 1 0 106100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7173
timestamp 1757982896
transform 1 0 107600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7174
timestamp 1757982896
transform 1 0 109100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7175
timestamp 1757982896
transform 1 0 110600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7176
timestamp 1757982896
transform 1 0 112100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7177
timestamp 1757982896
transform 1 0 113600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7178
timestamp 1757982896
transform 1 0 115100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7179
timestamp 1757982896
transform 1 0 116600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7180
timestamp 1757982896
transform 1 0 118100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7181
timestamp 1757982896
transform 1 0 119600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7182
timestamp 1757982896
transform 1 0 121100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7183
timestamp 1757982896
transform 1 0 122600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7184
timestamp 1757982896
transform 1 0 124100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7185
timestamp 1757982896
transform 1 0 125600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7186
timestamp 1757982896
transform 1 0 127100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7187
timestamp 1757982896
transform 1 0 128600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7188
timestamp 1757982896
transform 1 0 130100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7189
timestamp 1757982896
transform 1 0 131600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7190
timestamp 1757982896
transform 1 0 133100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7191
timestamp 1757982896
transform 1 0 134600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7192
timestamp 1757982896
transform 1 0 136100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7193
timestamp 1757982896
transform 1 0 137600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7194
timestamp 1757982896
transform 1 0 139100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7195
timestamp 1757982896
transform 1 0 140600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7196
timestamp 1757982896
transform 1 0 142100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7197
timestamp 1757982896
transform 1 0 143600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7198
timestamp 1757982896
transform 1 0 145100 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7199
timestamp 1757982896
transform 1 0 146600 0 1 -105150
box 1820 -1430 3480 230
use pixel  pixel_7200
timestamp 1757982896
transform 1 0 -1900 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7201
timestamp 1757982896
transform 1 0 -400 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7202
timestamp 1757982896
transform 1 0 1100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7203
timestamp 1757982896
transform 1 0 2600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7204
timestamp 1757982896
transform 1 0 4100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7205
timestamp 1757982896
transform 1 0 5600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7206
timestamp 1757982896
transform 1 0 7100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7207
timestamp 1757982896
transform 1 0 8600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7208
timestamp 1757982896
transform 1 0 10100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7209
timestamp 1757982896
transform 1 0 11600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7210
timestamp 1757982896
transform 1 0 13100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7211
timestamp 1757982896
transform 1 0 14600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7212
timestamp 1757982896
transform 1 0 16100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7213
timestamp 1757982896
transform 1 0 17600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7214
timestamp 1757982896
transform 1 0 19100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7215
timestamp 1757982896
transform 1 0 20600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7216
timestamp 1757982896
transform 1 0 22100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7217
timestamp 1757982896
transform 1 0 23600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7218
timestamp 1757982896
transform 1 0 25100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7219
timestamp 1757982896
transform 1 0 26600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7220
timestamp 1757982896
transform 1 0 28100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7221
timestamp 1757982896
transform 1 0 29600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7222
timestamp 1757982896
transform 1 0 31100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7223
timestamp 1757982896
transform 1 0 32600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7224
timestamp 1757982896
transform 1 0 34100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7225
timestamp 1757982896
transform 1 0 35600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7226
timestamp 1757982896
transform 1 0 37100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7227
timestamp 1757982896
transform 1 0 38600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7228
timestamp 1757982896
transform 1 0 40100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7229
timestamp 1757982896
transform 1 0 41600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7230
timestamp 1757982896
transform 1 0 43100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7231
timestamp 1757982896
transform 1 0 44600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7232
timestamp 1757982896
transform 1 0 46100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7233
timestamp 1757982896
transform 1 0 47600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7234
timestamp 1757982896
transform 1 0 49100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7235
timestamp 1757982896
transform 1 0 50600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7236
timestamp 1757982896
transform 1 0 52100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7237
timestamp 1757982896
transform 1 0 53600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7238
timestamp 1757982896
transform 1 0 55100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7239
timestamp 1757982896
transform 1 0 56600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7240
timestamp 1757982896
transform 1 0 58100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7241
timestamp 1757982896
transform 1 0 59600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7242
timestamp 1757982896
transform 1 0 61100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7243
timestamp 1757982896
transform 1 0 62600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7244
timestamp 1757982896
transform 1 0 64100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7245
timestamp 1757982896
transform 1 0 65600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7246
timestamp 1757982896
transform 1 0 67100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7247
timestamp 1757982896
transform 1 0 68600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7248
timestamp 1757982896
transform 1 0 70100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7249
timestamp 1757982896
transform 1 0 71600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7250
timestamp 1757982896
transform 1 0 73100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7251
timestamp 1757982896
transform 1 0 74600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7252
timestamp 1757982896
transform 1 0 76100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7253
timestamp 1757982896
transform 1 0 77600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7254
timestamp 1757982896
transform 1 0 79100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7255
timestamp 1757982896
transform 1 0 80600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7256
timestamp 1757982896
transform 1 0 82100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7257
timestamp 1757982896
transform 1 0 83600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7258
timestamp 1757982896
transform 1 0 85100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7259
timestamp 1757982896
transform 1 0 86600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7260
timestamp 1757982896
transform 1 0 88100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7261
timestamp 1757982896
transform 1 0 89600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7262
timestamp 1757982896
transform 1 0 91100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7263
timestamp 1757982896
transform 1 0 92600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7264
timestamp 1757982896
transform 1 0 94100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7265
timestamp 1757982896
transform 1 0 95600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7266
timestamp 1757982896
transform 1 0 97100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7267
timestamp 1757982896
transform 1 0 98600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7268
timestamp 1757982896
transform 1 0 100100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7269
timestamp 1757982896
transform 1 0 101600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7270
timestamp 1757982896
transform 1 0 103100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7271
timestamp 1757982896
transform 1 0 104600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7272
timestamp 1757982896
transform 1 0 106100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7273
timestamp 1757982896
transform 1 0 107600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7274
timestamp 1757982896
transform 1 0 109100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7275
timestamp 1757982896
transform 1 0 110600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7276
timestamp 1757982896
transform 1 0 112100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7277
timestamp 1757982896
transform 1 0 113600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7278
timestamp 1757982896
transform 1 0 115100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7279
timestamp 1757982896
transform 1 0 116600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7280
timestamp 1757982896
transform 1 0 118100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7281
timestamp 1757982896
transform 1 0 119600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7282
timestamp 1757982896
transform 1 0 121100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7283
timestamp 1757982896
transform 1 0 122600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7284
timestamp 1757982896
transform 1 0 124100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7285
timestamp 1757982896
transform 1 0 125600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7286
timestamp 1757982896
transform 1 0 127100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7287
timestamp 1757982896
transform 1 0 128600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7288
timestamp 1757982896
transform 1 0 130100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7289
timestamp 1757982896
transform 1 0 131600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7290
timestamp 1757982896
transform 1 0 133100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7291
timestamp 1757982896
transform 1 0 134600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7292
timestamp 1757982896
transform 1 0 136100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7293
timestamp 1757982896
transform 1 0 137600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7294
timestamp 1757982896
transform 1 0 139100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7295
timestamp 1757982896
transform 1 0 140600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7296
timestamp 1757982896
transform 1 0 142100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7297
timestamp 1757982896
transform 1 0 143600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7298
timestamp 1757982896
transform 1 0 145100 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7299
timestamp 1757982896
transform 1 0 146600 0 1 -106650
box 1820 -1430 3480 230
use pixel  pixel_7300
timestamp 1757982896
transform 1 0 -1900 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7301
timestamp 1757982896
transform 1 0 -400 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7302
timestamp 1757982896
transform 1 0 1100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7303
timestamp 1757982896
transform 1 0 2600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7304
timestamp 1757982896
transform 1 0 4100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7305
timestamp 1757982896
transform 1 0 5600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7306
timestamp 1757982896
transform 1 0 7100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7307
timestamp 1757982896
transform 1 0 8600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7308
timestamp 1757982896
transform 1 0 10100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7309
timestamp 1757982896
transform 1 0 11600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7310
timestamp 1757982896
transform 1 0 13100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7311
timestamp 1757982896
transform 1 0 14600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7312
timestamp 1757982896
transform 1 0 16100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7313
timestamp 1757982896
transform 1 0 17600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7314
timestamp 1757982896
transform 1 0 19100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7315
timestamp 1757982896
transform 1 0 20600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7316
timestamp 1757982896
transform 1 0 22100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7317
timestamp 1757982896
transform 1 0 23600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7318
timestamp 1757982896
transform 1 0 25100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7319
timestamp 1757982896
transform 1 0 26600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7320
timestamp 1757982896
transform 1 0 28100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7321
timestamp 1757982896
transform 1 0 29600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7322
timestamp 1757982896
transform 1 0 31100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7323
timestamp 1757982896
transform 1 0 32600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7324
timestamp 1757982896
transform 1 0 34100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7325
timestamp 1757982896
transform 1 0 35600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7326
timestamp 1757982896
transform 1 0 37100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7327
timestamp 1757982896
transform 1 0 38600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7328
timestamp 1757982896
transform 1 0 40100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7329
timestamp 1757982896
transform 1 0 41600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7330
timestamp 1757982896
transform 1 0 43100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7331
timestamp 1757982896
transform 1 0 44600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7332
timestamp 1757982896
transform 1 0 46100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7333
timestamp 1757982896
transform 1 0 47600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7334
timestamp 1757982896
transform 1 0 49100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7335
timestamp 1757982896
transform 1 0 50600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7336
timestamp 1757982896
transform 1 0 52100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7337
timestamp 1757982896
transform 1 0 53600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7338
timestamp 1757982896
transform 1 0 55100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7339
timestamp 1757982896
transform 1 0 56600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7340
timestamp 1757982896
transform 1 0 58100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7341
timestamp 1757982896
transform 1 0 59600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7342
timestamp 1757982896
transform 1 0 61100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7343
timestamp 1757982896
transform 1 0 62600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7344
timestamp 1757982896
transform 1 0 64100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7345
timestamp 1757982896
transform 1 0 65600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7346
timestamp 1757982896
transform 1 0 67100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7347
timestamp 1757982896
transform 1 0 68600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7348
timestamp 1757982896
transform 1 0 70100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7349
timestamp 1757982896
transform 1 0 71600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7350
timestamp 1757982896
transform 1 0 73100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7351
timestamp 1757982896
transform 1 0 74600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7352
timestamp 1757982896
transform 1 0 76100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7353
timestamp 1757982896
transform 1 0 77600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7354
timestamp 1757982896
transform 1 0 79100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7355
timestamp 1757982896
transform 1 0 80600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7356
timestamp 1757982896
transform 1 0 82100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7357
timestamp 1757982896
transform 1 0 83600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7358
timestamp 1757982896
transform 1 0 85100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7359
timestamp 1757982896
transform 1 0 86600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7360
timestamp 1757982896
transform 1 0 88100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7361
timestamp 1757982896
transform 1 0 89600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7362
timestamp 1757982896
transform 1 0 91100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7363
timestamp 1757982896
transform 1 0 92600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7364
timestamp 1757982896
transform 1 0 94100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7365
timestamp 1757982896
transform 1 0 95600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7366
timestamp 1757982896
transform 1 0 97100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7367
timestamp 1757982896
transform 1 0 98600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7368
timestamp 1757982896
transform 1 0 100100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7369
timestamp 1757982896
transform 1 0 101600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7370
timestamp 1757982896
transform 1 0 103100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7371
timestamp 1757982896
transform 1 0 104600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7372
timestamp 1757982896
transform 1 0 106100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7373
timestamp 1757982896
transform 1 0 107600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7374
timestamp 1757982896
transform 1 0 109100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7375
timestamp 1757982896
transform 1 0 110600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7376
timestamp 1757982896
transform 1 0 112100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7377
timestamp 1757982896
transform 1 0 113600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7378
timestamp 1757982896
transform 1 0 115100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7379
timestamp 1757982896
transform 1 0 116600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7380
timestamp 1757982896
transform 1 0 118100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7381
timestamp 1757982896
transform 1 0 119600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7382
timestamp 1757982896
transform 1 0 121100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7383
timestamp 1757982896
transform 1 0 122600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7384
timestamp 1757982896
transform 1 0 124100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7385
timestamp 1757982896
transform 1 0 125600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7386
timestamp 1757982896
transform 1 0 127100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7387
timestamp 1757982896
transform 1 0 128600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7388
timestamp 1757982896
transform 1 0 130100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7389
timestamp 1757982896
transform 1 0 131600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7390
timestamp 1757982896
transform 1 0 133100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7391
timestamp 1757982896
transform 1 0 134600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7392
timestamp 1757982896
transform 1 0 136100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7393
timestamp 1757982896
transform 1 0 137600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7394
timestamp 1757982896
transform 1 0 139100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7395
timestamp 1757982896
transform 1 0 140600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7396
timestamp 1757982896
transform 1 0 142100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7397
timestamp 1757982896
transform 1 0 143600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7398
timestamp 1757982896
transform 1 0 145100 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7399
timestamp 1757982896
transform 1 0 146600 0 1 -108150
box 1820 -1430 3480 230
use pixel  pixel_7400
timestamp 1757982896
transform 1 0 -1900 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7401
timestamp 1757982896
transform 1 0 -400 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7402
timestamp 1757982896
transform 1 0 1100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7403
timestamp 1757982896
transform 1 0 2600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7404
timestamp 1757982896
transform 1 0 4100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7405
timestamp 1757982896
transform 1 0 5600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7406
timestamp 1757982896
transform 1 0 7100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7407
timestamp 1757982896
transform 1 0 8600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7408
timestamp 1757982896
transform 1 0 10100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7409
timestamp 1757982896
transform 1 0 11600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7410
timestamp 1757982896
transform 1 0 13100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7411
timestamp 1757982896
transform 1 0 14600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7412
timestamp 1757982896
transform 1 0 16100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7413
timestamp 1757982896
transform 1 0 17600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7414
timestamp 1757982896
transform 1 0 19100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7415
timestamp 1757982896
transform 1 0 20600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7416
timestamp 1757982896
transform 1 0 22100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7417
timestamp 1757982896
transform 1 0 23600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7418
timestamp 1757982896
transform 1 0 25100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7419
timestamp 1757982896
transform 1 0 26600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7420
timestamp 1757982896
transform 1 0 28100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7421
timestamp 1757982896
transform 1 0 29600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7422
timestamp 1757982896
transform 1 0 31100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7423
timestamp 1757982896
transform 1 0 32600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7424
timestamp 1757982896
transform 1 0 34100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7425
timestamp 1757982896
transform 1 0 35600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7426
timestamp 1757982896
transform 1 0 37100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7427
timestamp 1757982896
transform 1 0 38600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7428
timestamp 1757982896
transform 1 0 40100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7429
timestamp 1757982896
transform 1 0 41600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7430
timestamp 1757982896
transform 1 0 43100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7431
timestamp 1757982896
transform 1 0 44600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7432
timestamp 1757982896
transform 1 0 46100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7433
timestamp 1757982896
transform 1 0 47600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7434
timestamp 1757982896
transform 1 0 49100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7435
timestamp 1757982896
transform 1 0 50600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7436
timestamp 1757982896
transform 1 0 52100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7437
timestamp 1757982896
transform 1 0 53600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7438
timestamp 1757982896
transform 1 0 55100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7439
timestamp 1757982896
transform 1 0 56600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7440
timestamp 1757982896
transform 1 0 58100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7441
timestamp 1757982896
transform 1 0 59600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7442
timestamp 1757982896
transform 1 0 61100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7443
timestamp 1757982896
transform 1 0 62600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7444
timestamp 1757982896
transform 1 0 64100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7445
timestamp 1757982896
transform 1 0 65600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7446
timestamp 1757982896
transform 1 0 67100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7447
timestamp 1757982896
transform 1 0 68600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7448
timestamp 1757982896
transform 1 0 70100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7449
timestamp 1757982896
transform 1 0 71600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7450
timestamp 1757982896
transform 1 0 73100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7451
timestamp 1757982896
transform 1 0 74600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7452
timestamp 1757982896
transform 1 0 76100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7453
timestamp 1757982896
transform 1 0 77600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7454
timestamp 1757982896
transform 1 0 79100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7455
timestamp 1757982896
transform 1 0 80600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7456
timestamp 1757982896
transform 1 0 82100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7457
timestamp 1757982896
transform 1 0 83600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7458
timestamp 1757982896
transform 1 0 85100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7459
timestamp 1757982896
transform 1 0 86600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7460
timestamp 1757982896
transform 1 0 88100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7461
timestamp 1757982896
transform 1 0 89600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7462
timestamp 1757982896
transform 1 0 91100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7463
timestamp 1757982896
transform 1 0 92600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7464
timestamp 1757982896
transform 1 0 94100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7465
timestamp 1757982896
transform 1 0 95600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7466
timestamp 1757982896
transform 1 0 97100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7467
timestamp 1757982896
transform 1 0 98600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7468
timestamp 1757982896
transform 1 0 100100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7469
timestamp 1757982896
transform 1 0 101600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7470
timestamp 1757982896
transform 1 0 103100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7471
timestamp 1757982896
transform 1 0 104600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7472
timestamp 1757982896
transform 1 0 106100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7473
timestamp 1757982896
transform 1 0 107600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7474
timestamp 1757982896
transform 1 0 109100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7475
timestamp 1757982896
transform 1 0 110600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7476
timestamp 1757982896
transform 1 0 112100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7477
timestamp 1757982896
transform 1 0 113600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7478
timestamp 1757982896
transform 1 0 115100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7479
timestamp 1757982896
transform 1 0 116600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7480
timestamp 1757982896
transform 1 0 118100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7481
timestamp 1757982896
transform 1 0 119600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7482
timestamp 1757982896
transform 1 0 121100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7483
timestamp 1757982896
transform 1 0 122600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7484
timestamp 1757982896
transform 1 0 124100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7485
timestamp 1757982896
transform 1 0 125600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7486
timestamp 1757982896
transform 1 0 127100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7487
timestamp 1757982896
transform 1 0 128600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7488
timestamp 1757982896
transform 1 0 130100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7489
timestamp 1757982896
transform 1 0 131600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7490
timestamp 1757982896
transform 1 0 133100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7491
timestamp 1757982896
transform 1 0 134600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7492
timestamp 1757982896
transform 1 0 136100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7493
timestamp 1757982896
transform 1 0 137600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7494
timestamp 1757982896
transform 1 0 139100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7495
timestamp 1757982896
transform 1 0 140600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7496
timestamp 1757982896
transform 1 0 142100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7497
timestamp 1757982896
transform 1 0 143600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7498
timestamp 1757982896
transform 1 0 145100 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7499
timestamp 1757982896
transform 1 0 146600 0 1 -109650
box 1820 -1430 3480 230
use pixel  pixel_7500
timestamp 1757982896
transform 1 0 -1900 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7501
timestamp 1757982896
transform 1 0 -400 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7502
timestamp 1757982896
transform 1 0 1100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7503
timestamp 1757982896
transform 1 0 2600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7504
timestamp 1757982896
transform 1 0 4100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7505
timestamp 1757982896
transform 1 0 5600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7506
timestamp 1757982896
transform 1 0 7100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7507
timestamp 1757982896
transform 1 0 8600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7508
timestamp 1757982896
transform 1 0 10100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7509
timestamp 1757982896
transform 1 0 11600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7510
timestamp 1757982896
transform 1 0 13100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7511
timestamp 1757982896
transform 1 0 14600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7512
timestamp 1757982896
transform 1 0 16100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7513
timestamp 1757982896
transform 1 0 17600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7514
timestamp 1757982896
transform 1 0 19100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7515
timestamp 1757982896
transform 1 0 20600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7516
timestamp 1757982896
transform 1 0 22100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7517
timestamp 1757982896
transform 1 0 23600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7518
timestamp 1757982896
transform 1 0 25100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7519
timestamp 1757982896
transform 1 0 26600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7520
timestamp 1757982896
transform 1 0 28100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7521
timestamp 1757982896
transform 1 0 29600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7522
timestamp 1757982896
transform 1 0 31100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7523
timestamp 1757982896
transform 1 0 32600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7524
timestamp 1757982896
transform 1 0 34100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7525
timestamp 1757982896
transform 1 0 35600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7526
timestamp 1757982896
transform 1 0 37100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7527
timestamp 1757982896
transform 1 0 38600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7528
timestamp 1757982896
transform 1 0 40100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7529
timestamp 1757982896
transform 1 0 41600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7530
timestamp 1757982896
transform 1 0 43100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7531
timestamp 1757982896
transform 1 0 44600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7532
timestamp 1757982896
transform 1 0 46100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7533
timestamp 1757982896
transform 1 0 47600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7534
timestamp 1757982896
transform 1 0 49100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7535
timestamp 1757982896
transform 1 0 50600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7536
timestamp 1757982896
transform 1 0 52100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7537
timestamp 1757982896
transform 1 0 53600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7538
timestamp 1757982896
transform 1 0 55100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7539
timestamp 1757982896
transform 1 0 56600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7540
timestamp 1757982896
transform 1 0 58100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7541
timestamp 1757982896
transform 1 0 59600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7542
timestamp 1757982896
transform 1 0 61100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7543
timestamp 1757982896
transform 1 0 62600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7544
timestamp 1757982896
transform 1 0 64100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7545
timestamp 1757982896
transform 1 0 65600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7546
timestamp 1757982896
transform 1 0 67100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7547
timestamp 1757982896
transform 1 0 68600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7548
timestamp 1757982896
transform 1 0 70100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7549
timestamp 1757982896
transform 1 0 71600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7550
timestamp 1757982896
transform 1 0 73100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7551
timestamp 1757982896
transform 1 0 74600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7552
timestamp 1757982896
transform 1 0 76100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7553
timestamp 1757982896
transform 1 0 77600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7554
timestamp 1757982896
transform 1 0 79100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7555
timestamp 1757982896
transform 1 0 80600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7556
timestamp 1757982896
transform 1 0 82100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7557
timestamp 1757982896
transform 1 0 83600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7558
timestamp 1757982896
transform 1 0 85100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7559
timestamp 1757982896
transform 1 0 86600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7560
timestamp 1757982896
transform 1 0 88100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7561
timestamp 1757982896
transform 1 0 89600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7562
timestamp 1757982896
transform 1 0 91100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7563
timestamp 1757982896
transform 1 0 92600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7564
timestamp 1757982896
transform 1 0 94100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7565
timestamp 1757982896
transform 1 0 95600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7566
timestamp 1757982896
transform 1 0 97100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7567
timestamp 1757982896
transform 1 0 98600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7568
timestamp 1757982896
transform 1 0 100100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7569
timestamp 1757982896
transform 1 0 101600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7570
timestamp 1757982896
transform 1 0 103100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7571
timestamp 1757982896
transform 1 0 104600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7572
timestamp 1757982896
transform 1 0 106100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7573
timestamp 1757982896
transform 1 0 107600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7574
timestamp 1757982896
transform 1 0 109100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7575
timestamp 1757982896
transform 1 0 110600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7576
timestamp 1757982896
transform 1 0 112100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7577
timestamp 1757982896
transform 1 0 113600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7578
timestamp 1757982896
transform 1 0 115100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7579
timestamp 1757982896
transform 1 0 116600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7580
timestamp 1757982896
transform 1 0 118100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7581
timestamp 1757982896
transform 1 0 119600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7582
timestamp 1757982896
transform 1 0 121100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7583
timestamp 1757982896
transform 1 0 122600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7584
timestamp 1757982896
transform 1 0 124100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7585
timestamp 1757982896
transform 1 0 125600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7586
timestamp 1757982896
transform 1 0 127100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7587
timestamp 1757982896
transform 1 0 128600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7588
timestamp 1757982896
transform 1 0 130100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7589
timestamp 1757982896
transform 1 0 131600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7590
timestamp 1757982896
transform 1 0 133100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7591
timestamp 1757982896
transform 1 0 134600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7592
timestamp 1757982896
transform 1 0 136100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7593
timestamp 1757982896
transform 1 0 137600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7594
timestamp 1757982896
transform 1 0 139100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7595
timestamp 1757982896
transform 1 0 140600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7596
timestamp 1757982896
transform 1 0 142100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7597
timestamp 1757982896
transform 1 0 143600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7598
timestamp 1757982896
transform 1 0 145100 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7599
timestamp 1757982896
transform 1 0 146600 0 1 -111150
box 1820 -1430 3480 230
use pixel  pixel_7600
timestamp 1757982896
transform 1 0 -1900 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7601
timestamp 1757982896
transform 1 0 -400 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7602
timestamp 1757982896
transform 1 0 1100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7603
timestamp 1757982896
transform 1 0 2600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7604
timestamp 1757982896
transform 1 0 4100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7605
timestamp 1757982896
transform 1 0 5600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7606
timestamp 1757982896
transform 1 0 7100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7607
timestamp 1757982896
transform 1 0 8600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7608
timestamp 1757982896
transform 1 0 10100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7609
timestamp 1757982896
transform 1 0 11600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7610
timestamp 1757982896
transform 1 0 13100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7611
timestamp 1757982896
transform 1 0 14600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7612
timestamp 1757982896
transform 1 0 16100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7613
timestamp 1757982896
transform 1 0 17600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7614
timestamp 1757982896
transform 1 0 19100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7615
timestamp 1757982896
transform 1 0 20600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7616
timestamp 1757982896
transform 1 0 22100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7617
timestamp 1757982896
transform 1 0 23600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7618
timestamp 1757982896
transform 1 0 25100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7619
timestamp 1757982896
transform 1 0 26600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7620
timestamp 1757982896
transform 1 0 28100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7621
timestamp 1757982896
transform 1 0 29600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7622
timestamp 1757982896
transform 1 0 31100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7623
timestamp 1757982896
transform 1 0 32600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7624
timestamp 1757982896
transform 1 0 34100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7625
timestamp 1757982896
transform 1 0 35600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7626
timestamp 1757982896
transform 1 0 37100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7627
timestamp 1757982896
transform 1 0 38600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7628
timestamp 1757982896
transform 1 0 40100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7629
timestamp 1757982896
transform 1 0 41600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7630
timestamp 1757982896
transform 1 0 43100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7631
timestamp 1757982896
transform 1 0 44600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7632
timestamp 1757982896
transform 1 0 46100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7633
timestamp 1757982896
transform 1 0 47600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7634
timestamp 1757982896
transform 1 0 49100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7635
timestamp 1757982896
transform 1 0 50600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7636
timestamp 1757982896
transform 1 0 52100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7637
timestamp 1757982896
transform 1 0 53600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7638
timestamp 1757982896
transform 1 0 55100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7639
timestamp 1757982896
transform 1 0 56600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7640
timestamp 1757982896
transform 1 0 58100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7641
timestamp 1757982896
transform 1 0 59600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7642
timestamp 1757982896
transform 1 0 61100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7643
timestamp 1757982896
transform 1 0 62600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7644
timestamp 1757982896
transform 1 0 64100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7645
timestamp 1757982896
transform 1 0 65600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7646
timestamp 1757982896
transform 1 0 67100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7647
timestamp 1757982896
transform 1 0 68600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7648
timestamp 1757982896
transform 1 0 70100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7649
timestamp 1757982896
transform 1 0 71600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7650
timestamp 1757982896
transform 1 0 73100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7651
timestamp 1757982896
transform 1 0 74600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7652
timestamp 1757982896
transform 1 0 76100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7653
timestamp 1757982896
transform 1 0 77600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7654
timestamp 1757982896
transform 1 0 79100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7655
timestamp 1757982896
transform 1 0 80600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7656
timestamp 1757982896
transform 1 0 82100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7657
timestamp 1757982896
transform 1 0 83600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7658
timestamp 1757982896
transform 1 0 85100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7659
timestamp 1757982896
transform 1 0 86600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7660
timestamp 1757982896
transform 1 0 88100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7661
timestamp 1757982896
transform 1 0 89600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7662
timestamp 1757982896
transform 1 0 91100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7663
timestamp 1757982896
transform 1 0 92600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7664
timestamp 1757982896
transform 1 0 94100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7665
timestamp 1757982896
transform 1 0 95600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7666
timestamp 1757982896
transform 1 0 97100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7667
timestamp 1757982896
transform 1 0 98600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7668
timestamp 1757982896
transform 1 0 100100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7669
timestamp 1757982896
transform 1 0 101600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7670
timestamp 1757982896
transform 1 0 103100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7671
timestamp 1757982896
transform 1 0 104600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7672
timestamp 1757982896
transform 1 0 106100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7673
timestamp 1757982896
transform 1 0 107600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7674
timestamp 1757982896
transform 1 0 109100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7675
timestamp 1757982896
transform 1 0 110600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7676
timestamp 1757982896
transform 1 0 112100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7677
timestamp 1757982896
transform 1 0 113600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7678
timestamp 1757982896
transform 1 0 115100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7679
timestamp 1757982896
transform 1 0 116600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7680
timestamp 1757982896
transform 1 0 118100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7681
timestamp 1757982896
transform 1 0 119600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7682
timestamp 1757982896
transform 1 0 121100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7683
timestamp 1757982896
transform 1 0 122600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7684
timestamp 1757982896
transform 1 0 124100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7685
timestamp 1757982896
transform 1 0 125600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7686
timestamp 1757982896
transform 1 0 127100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7687
timestamp 1757982896
transform 1 0 128600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7688
timestamp 1757982896
transform 1 0 130100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7689
timestamp 1757982896
transform 1 0 131600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7690
timestamp 1757982896
transform 1 0 133100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7691
timestamp 1757982896
transform 1 0 134600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7692
timestamp 1757982896
transform 1 0 136100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7693
timestamp 1757982896
transform 1 0 137600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7694
timestamp 1757982896
transform 1 0 139100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7695
timestamp 1757982896
transform 1 0 140600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7696
timestamp 1757982896
transform 1 0 142100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7697
timestamp 1757982896
transform 1 0 143600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7698
timestamp 1757982896
transform 1 0 145100 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7699
timestamp 1757982896
transform 1 0 146600 0 1 -112650
box 1820 -1430 3480 230
use pixel  pixel_7700
timestamp 1757982896
transform 1 0 -1900 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7701
timestamp 1757982896
transform 1 0 -400 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7702
timestamp 1757982896
transform 1 0 1100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7703
timestamp 1757982896
transform 1 0 2600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7704
timestamp 1757982896
transform 1 0 4100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7705
timestamp 1757982896
transform 1 0 5600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7706
timestamp 1757982896
transform 1 0 7100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7707
timestamp 1757982896
transform 1 0 8600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7708
timestamp 1757982896
transform 1 0 10100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7709
timestamp 1757982896
transform 1 0 11600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7710
timestamp 1757982896
transform 1 0 13100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7711
timestamp 1757982896
transform 1 0 14600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7712
timestamp 1757982896
transform 1 0 16100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7713
timestamp 1757982896
transform 1 0 17600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7714
timestamp 1757982896
transform 1 0 19100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7715
timestamp 1757982896
transform 1 0 20600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7716
timestamp 1757982896
transform 1 0 22100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7717
timestamp 1757982896
transform 1 0 23600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7718
timestamp 1757982896
transform 1 0 25100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7719
timestamp 1757982896
transform 1 0 26600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7720
timestamp 1757982896
transform 1 0 28100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7721
timestamp 1757982896
transform 1 0 29600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7722
timestamp 1757982896
transform 1 0 31100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7723
timestamp 1757982896
transform 1 0 32600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7724
timestamp 1757982896
transform 1 0 34100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7725
timestamp 1757982896
transform 1 0 35600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7726
timestamp 1757982896
transform 1 0 37100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7727
timestamp 1757982896
transform 1 0 38600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7728
timestamp 1757982896
transform 1 0 40100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7729
timestamp 1757982896
transform 1 0 41600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7730
timestamp 1757982896
transform 1 0 43100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7731
timestamp 1757982896
transform 1 0 44600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7732
timestamp 1757982896
transform 1 0 46100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7733
timestamp 1757982896
transform 1 0 47600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7734
timestamp 1757982896
transform 1 0 49100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7735
timestamp 1757982896
transform 1 0 50600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7736
timestamp 1757982896
transform 1 0 52100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7737
timestamp 1757982896
transform 1 0 53600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7738
timestamp 1757982896
transform 1 0 55100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7739
timestamp 1757982896
transform 1 0 56600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7740
timestamp 1757982896
transform 1 0 58100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7741
timestamp 1757982896
transform 1 0 59600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7742
timestamp 1757982896
transform 1 0 61100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7743
timestamp 1757982896
transform 1 0 62600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7744
timestamp 1757982896
transform 1 0 64100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7745
timestamp 1757982896
transform 1 0 65600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7746
timestamp 1757982896
transform 1 0 67100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7747
timestamp 1757982896
transform 1 0 68600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7748
timestamp 1757982896
transform 1 0 70100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7749
timestamp 1757982896
transform 1 0 71600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7750
timestamp 1757982896
transform 1 0 73100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7751
timestamp 1757982896
transform 1 0 74600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7752
timestamp 1757982896
transform 1 0 76100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7753
timestamp 1757982896
transform 1 0 77600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7754
timestamp 1757982896
transform 1 0 79100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7755
timestamp 1757982896
transform 1 0 80600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7756
timestamp 1757982896
transform 1 0 82100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7757
timestamp 1757982896
transform 1 0 83600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7758
timestamp 1757982896
transform 1 0 85100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7759
timestamp 1757982896
transform 1 0 86600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7760
timestamp 1757982896
transform 1 0 88100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7761
timestamp 1757982896
transform 1 0 89600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7762
timestamp 1757982896
transform 1 0 91100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7763
timestamp 1757982896
transform 1 0 92600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7764
timestamp 1757982896
transform 1 0 94100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7765
timestamp 1757982896
transform 1 0 95600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7766
timestamp 1757982896
transform 1 0 97100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7767
timestamp 1757982896
transform 1 0 98600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7768
timestamp 1757982896
transform 1 0 100100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7769
timestamp 1757982896
transform 1 0 101600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7770
timestamp 1757982896
transform 1 0 103100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7771
timestamp 1757982896
transform 1 0 104600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7772
timestamp 1757982896
transform 1 0 106100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7773
timestamp 1757982896
transform 1 0 107600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7774
timestamp 1757982896
transform 1 0 109100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7775
timestamp 1757982896
transform 1 0 110600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7776
timestamp 1757982896
transform 1 0 112100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7777
timestamp 1757982896
transform 1 0 113600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7778
timestamp 1757982896
transform 1 0 115100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7779
timestamp 1757982896
transform 1 0 116600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7780
timestamp 1757982896
transform 1 0 118100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7781
timestamp 1757982896
transform 1 0 119600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7782
timestamp 1757982896
transform 1 0 121100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7783
timestamp 1757982896
transform 1 0 122600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7784
timestamp 1757982896
transform 1 0 124100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7785
timestamp 1757982896
transform 1 0 125600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7786
timestamp 1757982896
transform 1 0 127100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7787
timestamp 1757982896
transform 1 0 128600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7788
timestamp 1757982896
transform 1 0 130100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7789
timestamp 1757982896
transform 1 0 131600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7790
timestamp 1757982896
transform 1 0 133100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7791
timestamp 1757982896
transform 1 0 134600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7792
timestamp 1757982896
transform 1 0 136100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7793
timestamp 1757982896
transform 1 0 137600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7794
timestamp 1757982896
transform 1 0 139100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7795
timestamp 1757982896
transform 1 0 140600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7796
timestamp 1757982896
transform 1 0 142100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7797
timestamp 1757982896
transform 1 0 143600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7798
timestamp 1757982896
transform 1 0 145100 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7799
timestamp 1757982896
transform 1 0 146600 0 1 -114150
box 1820 -1430 3480 230
use pixel  pixel_7800
timestamp 1757982896
transform 1 0 -1900 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7801
timestamp 1757982896
transform 1 0 -400 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7802
timestamp 1757982896
transform 1 0 1100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7803
timestamp 1757982896
transform 1 0 2600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7804
timestamp 1757982896
transform 1 0 4100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7805
timestamp 1757982896
transform 1 0 5600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7806
timestamp 1757982896
transform 1 0 7100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7807
timestamp 1757982896
transform 1 0 8600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7808
timestamp 1757982896
transform 1 0 10100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7809
timestamp 1757982896
transform 1 0 11600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7810
timestamp 1757982896
transform 1 0 13100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7811
timestamp 1757982896
transform 1 0 14600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7812
timestamp 1757982896
transform 1 0 16100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7813
timestamp 1757982896
transform 1 0 17600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7814
timestamp 1757982896
transform 1 0 19100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7815
timestamp 1757982896
transform 1 0 20600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7816
timestamp 1757982896
transform 1 0 22100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7817
timestamp 1757982896
transform 1 0 23600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7818
timestamp 1757982896
transform 1 0 25100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7819
timestamp 1757982896
transform 1 0 26600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7820
timestamp 1757982896
transform 1 0 28100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7821
timestamp 1757982896
transform 1 0 29600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7822
timestamp 1757982896
transform 1 0 31100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7823
timestamp 1757982896
transform 1 0 32600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7824
timestamp 1757982896
transform 1 0 34100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7825
timestamp 1757982896
transform 1 0 35600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7826
timestamp 1757982896
transform 1 0 37100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7827
timestamp 1757982896
transform 1 0 38600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7828
timestamp 1757982896
transform 1 0 40100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7829
timestamp 1757982896
transform 1 0 41600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7830
timestamp 1757982896
transform 1 0 43100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7831
timestamp 1757982896
transform 1 0 44600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7832
timestamp 1757982896
transform 1 0 46100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7833
timestamp 1757982896
transform 1 0 47600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7834
timestamp 1757982896
transform 1 0 49100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7835
timestamp 1757982896
transform 1 0 50600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7836
timestamp 1757982896
transform 1 0 52100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7837
timestamp 1757982896
transform 1 0 53600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7838
timestamp 1757982896
transform 1 0 55100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7839
timestamp 1757982896
transform 1 0 56600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7840
timestamp 1757982896
transform 1 0 58100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7841
timestamp 1757982896
transform 1 0 59600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7842
timestamp 1757982896
transform 1 0 61100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7843
timestamp 1757982896
transform 1 0 62600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7844
timestamp 1757982896
transform 1 0 64100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7845
timestamp 1757982896
transform 1 0 65600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7846
timestamp 1757982896
transform 1 0 67100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7847
timestamp 1757982896
transform 1 0 68600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7848
timestamp 1757982896
transform 1 0 70100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7849
timestamp 1757982896
transform 1 0 71600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7850
timestamp 1757982896
transform 1 0 73100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7851
timestamp 1757982896
transform 1 0 74600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7852
timestamp 1757982896
transform 1 0 76100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7853
timestamp 1757982896
transform 1 0 77600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7854
timestamp 1757982896
transform 1 0 79100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7855
timestamp 1757982896
transform 1 0 80600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7856
timestamp 1757982896
transform 1 0 82100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7857
timestamp 1757982896
transform 1 0 83600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7858
timestamp 1757982896
transform 1 0 85100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7859
timestamp 1757982896
transform 1 0 86600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7860
timestamp 1757982896
transform 1 0 88100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7861
timestamp 1757982896
transform 1 0 89600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7862
timestamp 1757982896
transform 1 0 91100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7863
timestamp 1757982896
transform 1 0 92600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7864
timestamp 1757982896
transform 1 0 94100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7865
timestamp 1757982896
transform 1 0 95600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7866
timestamp 1757982896
transform 1 0 97100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7867
timestamp 1757982896
transform 1 0 98600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7868
timestamp 1757982896
transform 1 0 100100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7869
timestamp 1757982896
transform 1 0 101600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7870
timestamp 1757982896
transform 1 0 103100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7871
timestamp 1757982896
transform 1 0 104600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7872
timestamp 1757982896
transform 1 0 106100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7873
timestamp 1757982896
transform 1 0 107600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7874
timestamp 1757982896
transform 1 0 109100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7875
timestamp 1757982896
transform 1 0 110600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7876
timestamp 1757982896
transform 1 0 112100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7877
timestamp 1757982896
transform 1 0 113600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7878
timestamp 1757982896
transform 1 0 115100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7879
timestamp 1757982896
transform 1 0 116600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7880
timestamp 1757982896
transform 1 0 118100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7881
timestamp 1757982896
transform 1 0 119600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7882
timestamp 1757982896
transform 1 0 121100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7883
timestamp 1757982896
transform 1 0 122600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7884
timestamp 1757982896
transform 1 0 124100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7885
timestamp 1757982896
transform 1 0 125600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7886
timestamp 1757982896
transform 1 0 127100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7887
timestamp 1757982896
transform 1 0 128600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7888
timestamp 1757982896
transform 1 0 130100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7889
timestamp 1757982896
transform 1 0 131600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7890
timestamp 1757982896
transform 1 0 133100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7891
timestamp 1757982896
transform 1 0 134600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7892
timestamp 1757982896
transform 1 0 136100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7893
timestamp 1757982896
transform 1 0 137600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7894
timestamp 1757982896
transform 1 0 139100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7895
timestamp 1757982896
transform 1 0 140600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7896
timestamp 1757982896
transform 1 0 142100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7897
timestamp 1757982896
transform 1 0 143600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7898
timestamp 1757982896
transform 1 0 145100 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7899
timestamp 1757982896
transform 1 0 146600 0 1 -115650
box 1820 -1430 3480 230
use pixel  pixel_7900
timestamp 1757982896
transform 1 0 -1900 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7901
timestamp 1757982896
transform 1 0 -400 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7902
timestamp 1757982896
transform 1 0 1100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7903
timestamp 1757982896
transform 1 0 2600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7904
timestamp 1757982896
transform 1 0 4100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7905
timestamp 1757982896
transform 1 0 5600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7906
timestamp 1757982896
transform 1 0 7100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7907
timestamp 1757982896
transform 1 0 8600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7908
timestamp 1757982896
transform 1 0 10100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7909
timestamp 1757982896
transform 1 0 11600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7910
timestamp 1757982896
transform 1 0 13100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7911
timestamp 1757982896
transform 1 0 14600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7912
timestamp 1757982896
transform 1 0 16100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7913
timestamp 1757982896
transform 1 0 17600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7914
timestamp 1757982896
transform 1 0 19100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7915
timestamp 1757982896
transform 1 0 20600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7916
timestamp 1757982896
transform 1 0 22100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7917
timestamp 1757982896
transform 1 0 23600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7918
timestamp 1757982896
transform 1 0 25100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7919
timestamp 1757982896
transform 1 0 26600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7920
timestamp 1757982896
transform 1 0 28100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7921
timestamp 1757982896
transform 1 0 29600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7922
timestamp 1757982896
transform 1 0 31100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7923
timestamp 1757982896
transform 1 0 32600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7924
timestamp 1757982896
transform 1 0 34100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7925
timestamp 1757982896
transform 1 0 35600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7926
timestamp 1757982896
transform 1 0 37100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7927
timestamp 1757982896
transform 1 0 38600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7928
timestamp 1757982896
transform 1 0 40100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7929
timestamp 1757982896
transform 1 0 41600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7930
timestamp 1757982896
transform 1 0 43100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7931
timestamp 1757982896
transform 1 0 44600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7932
timestamp 1757982896
transform 1 0 46100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7933
timestamp 1757982896
transform 1 0 47600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7934
timestamp 1757982896
transform 1 0 49100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7935
timestamp 1757982896
transform 1 0 50600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7936
timestamp 1757982896
transform 1 0 52100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7937
timestamp 1757982896
transform 1 0 53600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7938
timestamp 1757982896
transform 1 0 55100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7939
timestamp 1757982896
transform 1 0 56600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7940
timestamp 1757982896
transform 1 0 58100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7941
timestamp 1757982896
transform 1 0 59600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7942
timestamp 1757982896
transform 1 0 61100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7943
timestamp 1757982896
transform 1 0 62600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7944
timestamp 1757982896
transform 1 0 64100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7945
timestamp 1757982896
transform 1 0 65600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7946
timestamp 1757982896
transform 1 0 67100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7947
timestamp 1757982896
transform 1 0 68600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7948
timestamp 1757982896
transform 1 0 70100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7949
timestamp 1757982896
transform 1 0 71600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7950
timestamp 1757982896
transform 1 0 73100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7951
timestamp 1757982896
transform 1 0 74600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7952
timestamp 1757982896
transform 1 0 76100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7953
timestamp 1757982896
transform 1 0 77600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7954
timestamp 1757982896
transform 1 0 79100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7955
timestamp 1757982896
transform 1 0 80600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7956
timestamp 1757982896
transform 1 0 82100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7957
timestamp 1757982896
transform 1 0 83600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7958
timestamp 1757982896
transform 1 0 85100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7959
timestamp 1757982896
transform 1 0 86600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7960
timestamp 1757982896
transform 1 0 88100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7961
timestamp 1757982896
transform 1 0 89600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7962
timestamp 1757982896
transform 1 0 91100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7963
timestamp 1757982896
transform 1 0 92600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7964
timestamp 1757982896
transform 1 0 94100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7965
timestamp 1757982896
transform 1 0 95600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7966
timestamp 1757982896
transform 1 0 97100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7967
timestamp 1757982896
transform 1 0 98600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7968
timestamp 1757982896
transform 1 0 100100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7969
timestamp 1757982896
transform 1 0 101600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7970
timestamp 1757982896
transform 1 0 103100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7971
timestamp 1757982896
transform 1 0 104600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7972
timestamp 1757982896
transform 1 0 106100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7973
timestamp 1757982896
transform 1 0 107600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7974
timestamp 1757982896
transform 1 0 109100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7975
timestamp 1757982896
transform 1 0 110600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7976
timestamp 1757982896
transform 1 0 112100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7977
timestamp 1757982896
transform 1 0 113600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7978
timestamp 1757982896
transform 1 0 115100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7979
timestamp 1757982896
transform 1 0 116600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7980
timestamp 1757982896
transform 1 0 118100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7981
timestamp 1757982896
transform 1 0 119600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7982
timestamp 1757982896
transform 1 0 121100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7983
timestamp 1757982896
transform 1 0 122600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7984
timestamp 1757982896
transform 1 0 124100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7985
timestamp 1757982896
transform 1 0 125600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7986
timestamp 1757982896
transform 1 0 127100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7987
timestamp 1757982896
transform 1 0 128600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7988
timestamp 1757982896
transform 1 0 130100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7989
timestamp 1757982896
transform 1 0 131600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7990
timestamp 1757982896
transform 1 0 133100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7991
timestamp 1757982896
transform 1 0 134600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7992
timestamp 1757982896
transform 1 0 136100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7993
timestamp 1757982896
transform 1 0 137600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7994
timestamp 1757982896
transform 1 0 139100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7995
timestamp 1757982896
transform 1 0 140600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7996
timestamp 1757982896
transform 1 0 142100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7997
timestamp 1757982896
transform 1 0 143600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7998
timestamp 1757982896
transform 1 0 145100 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_7999
timestamp 1757982896
transform 1 0 146600 0 1 -117150
box 1820 -1430 3480 230
use pixel  pixel_8000
timestamp 1757982896
transform 1 0 -1900 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8001
timestamp 1757982896
transform 1 0 -400 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8002
timestamp 1757982896
transform 1 0 1100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8003
timestamp 1757982896
transform 1 0 2600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8004
timestamp 1757982896
transform 1 0 4100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8005
timestamp 1757982896
transform 1 0 5600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8006
timestamp 1757982896
transform 1 0 7100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8007
timestamp 1757982896
transform 1 0 8600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8008
timestamp 1757982896
transform 1 0 10100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8009
timestamp 1757982896
transform 1 0 11600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8010
timestamp 1757982896
transform 1 0 13100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8011
timestamp 1757982896
transform 1 0 14600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8012
timestamp 1757982896
transform 1 0 16100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8013
timestamp 1757982896
transform 1 0 17600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8014
timestamp 1757982896
transform 1 0 19100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8015
timestamp 1757982896
transform 1 0 20600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8016
timestamp 1757982896
transform 1 0 22100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8017
timestamp 1757982896
transform 1 0 23600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8018
timestamp 1757982896
transform 1 0 25100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8019
timestamp 1757982896
transform 1 0 26600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8020
timestamp 1757982896
transform 1 0 28100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8021
timestamp 1757982896
transform 1 0 29600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8022
timestamp 1757982896
transform 1 0 31100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8023
timestamp 1757982896
transform 1 0 32600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8024
timestamp 1757982896
transform 1 0 34100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8025
timestamp 1757982896
transform 1 0 35600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8026
timestamp 1757982896
transform 1 0 37100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8027
timestamp 1757982896
transform 1 0 38600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8028
timestamp 1757982896
transform 1 0 40100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8029
timestamp 1757982896
transform 1 0 41600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8030
timestamp 1757982896
transform 1 0 43100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8031
timestamp 1757982896
transform 1 0 44600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8032
timestamp 1757982896
transform 1 0 46100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8033
timestamp 1757982896
transform 1 0 47600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8034
timestamp 1757982896
transform 1 0 49100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8035
timestamp 1757982896
transform 1 0 50600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8036
timestamp 1757982896
transform 1 0 52100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8037
timestamp 1757982896
transform 1 0 53600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8038
timestamp 1757982896
transform 1 0 55100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8039
timestamp 1757982896
transform 1 0 56600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8040
timestamp 1757982896
transform 1 0 58100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8041
timestamp 1757982896
transform 1 0 59600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8042
timestamp 1757982896
transform 1 0 61100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8043
timestamp 1757982896
transform 1 0 62600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8044
timestamp 1757982896
transform 1 0 64100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8045
timestamp 1757982896
transform 1 0 65600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8046
timestamp 1757982896
transform 1 0 67100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8047
timestamp 1757982896
transform 1 0 68600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8048
timestamp 1757982896
transform 1 0 70100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8049
timestamp 1757982896
transform 1 0 71600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8050
timestamp 1757982896
transform 1 0 73100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8051
timestamp 1757982896
transform 1 0 74600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8052
timestamp 1757982896
transform 1 0 76100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8053
timestamp 1757982896
transform 1 0 77600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8054
timestamp 1757982896
transform 1 0 79100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8055
timestamp 1757982896
transform 1 0 80600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8056
timestamp 1757982896
transform 1 0 82100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8057
timestamp 1757982896
transform 1 0 83600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8058
timestamp 1757982896
transform 1 0 85100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8059
timestamp 1757982896
transform 1 0 86600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8060
timestamp 1757982896
transform 1 0 88100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8061
timestamp 1757982896
transform 1 0 89600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8062
timestamp 1757982896
transform 1 0 91100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8063
timestamp 1757982896
transform 1 0 92600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8064
timestamp 1757982896
transform 1 0 94100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8065
timestamp 1757982896
transform 1 0 95600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8066
timestamp 1757982896
transform 1 0 97100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8067
timestamp 1757982896
transform 1 0 98600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8068
timestamp 1757982896
transform 1 0 100100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8069
timestamp 1757982896
transform 1 0 101600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8070
timestamp 1757982896
transform 1 0 103100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8071
timestamp 1757982896
transform 1 0 104600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8072
timestamp 1757982896
transform 1 0 106100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8073
timestamp 1757982896
transform 1 0 107600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8074
timestamp 1757982896
transform 1 0 109100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8075
timestamp 1757982896
transform 1 0 110600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8076
timestamp 1757982896
transform 1 0 112100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8077
timestamp 1757982896
transform 1 0 113600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8078
timestamp 1757982896
transform 1 0 115100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8079
timestamp 1757982896
transform 1 0 116600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8080
timestamp 1757982896
transform 1 0 118100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8081
timestamp 1757982896
transform 1 0 119600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8082
timestamp 1757982896
transform 1 0 121100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8083
timestamp 1757982896
transform 1 0 122600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8084
timestamp 1757982896
transform 1 0 124100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8085
timestamp 1757982896
transform 1 0 125600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8086
timestamp 1757982896
transform 1 0 127100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8087
timestamp 1757982896
transform 1 0 128600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8088
timestamp 1757982896
transform 1 0 130100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8089
timestamp 1757982896
transform 1 0 131600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8090
timestamp 1757982896
transform 1 0 133100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8091
timestamp 1757982896
transform 1 0 134600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8092
timestamp 1757982896
transform 1 0 136100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8093
timestamp 1757982896
transform 1 0 137600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8094
timestamp 1757982896
transform 1 0 139100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8095
timestamp 1757982896
transform 1 0 140600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8096
timestamp 1757982896
transform 1 0 142100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8097
timestamp 1757982896
transform 1 0 143600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8098
timestamp 1757982896
transform 1 0 145100 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8099
timestamp 1757982896
transform 1 0 146600 0 1 -118650
box 1820 -1430 3480 230
use pixel  pixel_8100
timestamp 1757982896
transform 1 0 -1900 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8101
timestamp 1757982896
transform 1 0 -400 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8102
timestamp 1757982896
transform 1 0 1100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8103
timestamp 1757982896
transform 1 0 2600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8104
timestamp 1757982896
transform 1 0 4100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8105
timestamp 1757982896
transform 1 0 5600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8106
timestamp 1757982896
transform 1 0 7100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8107
timestamp 1757982896
transform 1 0 8600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8108
timestamp 1757982896
transform 1 0 10100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8109
timestamp 1757982896
transform 1 0 11600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8110
timestamp 1757982896
transform 1 0 13100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8111
timestamp 1757982896
transform 1 0 14600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8112
timestamp 1757982896
transform 1 0 16100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8113
timestamp 1757982896
transform 1 0 17600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8114
timestamp 1757982896
transform 1 0 19100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8115
timestamp 1757982896
transform 1 0 20600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8116
timestamp 1757982896
transform 1 0 22100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8117
timestamp 1757982896
transform 1 0 23600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8118
timestamp 1757982896
transform 1 0 25100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8119
timestamp 1757982896
transform 1 0 26600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8120
timestamp 1757982896
transform 1 0 28100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8121
timestamp 1757982896
transform 1 0 29600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8122
timestamp 1757982896
transform 1 0 31100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8123
timestamp 1757982896
transform 1 0 32600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8124
timestamp 1757982896
transform 1 0 34100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8125
timestamp 1757982896
transform 1 0 35600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8126
timestamp 1757982896
transform 1 0 37100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8127
timestamp 1757982896
transform 1 0 38600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8128
timestamp 1757982896
transform 1 0 40100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8129
timestamp 1757982896
transform 1 0 41600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8130
timestamp 1757982896
transform 1 0 43100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8131
timestamp 1757982896
transform 1 0 44600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8132
timestamp 1757982896
transform 1 0 46100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8133
timestamp 1757982896
transform 1 0 47600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8134
timestamp 1757982896
transform 1 0 49100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8135
timestamp 1757982896
transform 1 0 50600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8136
timestamp 1757982896
transform 1 0 52100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8137
timestamp 1757982896
transform 1 0 53600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8138
timestamp 1757982896
transform 1 0 55100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8139
timestamp 1757982896
transform 1 0 56600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8140
timestamp 1757982896
transform 1 0 58100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8141
timestamp 1757982896
transform 1 0 59600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8142
timestamp 1757982896
transform 1 0 61100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8143
timestamp 1757982896
transform 1 0 62600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8144
timestamp 1757982896
transform 1 0 64100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8145
timestamp 1757982896
transform 1 0 65600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8146
timestamp 1757982896
transform 1 0 67100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8147
timestamp 1757982896
transform 1 0 68600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8148
timestamp 1757982896
transform 1 0 70100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8149
timestamp 1757982896
transform 1 0 71600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8150
timestamp 1757982896
transform 1 0 73100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8151
timestamp 1757982896
transform 1 0 74600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8152
timestamp 1757982896
transform 1 0 76100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8153
timestamp 1757982896
transform 1 0 77600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8154
timestamp 1757982896
transform 1 0 79100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8155
timestamp 1757982896
transform 1 0 80600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8156
timestamp 1757982896
transform 1 0 82100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8157
timestamp 1757982896
transform 1 0 83600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8158
timestamp 1757982896
transform 1 0 85100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8159
timestamp 1757982896
transform 1 0 86600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8160
timestamp 1757982896
transform 1 0 88100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8161
timestamp 1757982896
transform 1 0 89600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8162
timestamp 1757982896
transform 1 0 91100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8163
timestamp 1757982896
transform 1 0 92600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8164
timestamp 1757982896
transform 1 0 94100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8165
timestamp 1757982896
transform 1 0 95600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8166
timestamp 1757982896
transform 1 0 97100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8167
timestamp 1757982896
transform 1 0 98600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8168
timestamp 1757982896
transform 1 0 100100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8169
timestamp 1757982896
transform 1 0 101600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8170
timestamp 1757982896
transform 1 0 103100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8171
timestamp 1757982896
transform 1 0 104600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8172
timestamp 1757982896
transform 1 0 106100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8173
timestamp 1757982896
transform 1 0 107600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8174
timestamp 1757982896
transform 1 0 109100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8175
timestamp 1757982896
transform 1 0 110600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8176
timestamp 1757982896
transform 1 0 112100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8177
timestamp 1757982896
transform 1 0 113600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8178
timestamp 1757982896
transform 1 0 115100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8179
timestamp 1757982896
transform 1 0 116600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8180
timestamp 1757982896
transform 1 0 118100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8181
timestamp 1757982896
transform 1 0 119600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8182
timestamp 1757982896
transform 1 0 121100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8183
timestamp 1757982896
transform 1 0 122600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8184
timestamp 1757982896
transform 1 0 124100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8185
timestamp 1757982896
transform 1 0 125600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8186
timestamp 1757982896
transform 1 0 127100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8187
timestamp 1757982896
transform 1 0 128600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8188
timestamp 1757982896
transform 1 0 130100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8189
timestamp 1757982896
transform 1 0 131600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8190
timestamp 1757982896
transform 1 0 133100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8191
timestamp 1757982896
transform 1 0 134600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8192
timestamp 1757982896
transform 1 0 136100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8193
timestamp 1757982896
transform 1 0 137600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8194
timestamp 1757982896
transform 1 0 139100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8195
timestamp 1757982896
transform 1 0 140600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8196
timestamp 1757982896
transform 1 0 142100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8197
timestamp 1757982896
transform 1 0 143600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8198
timestamp 1757982896
transform 1 0 145100 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8199
timestamp 1757982896
transform 1 0 146600 0 1 -120150
box 1820 -1430 3480 230
use pixel  pixel_8200
timestamp 1757982896
transform 1 0 -1900 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8201
timestamp 1757982896
transform 1 0 -400 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8202
timestamp 1757982896
transform 1 0 1100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8203
timestamp 1757982896
transform 1 0 2600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8204
timestamp 1757982896
transform 1 0 4100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8205
timestamp 1757982896
transform 1 0 5600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8206
timestamp 1757982896
transform 1 0 7100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8207
timestamp 1757982896
transform 1 0 8600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8208
timestamp 1757982896
transform 1 0 10100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8209
timestamp 1757982896
transform 1 0 11600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8210
timestamp 1757982896
transform 1 0 13100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8211
timestamp 1757982896
transform 1 0 14600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8212
timestamp 1757982896
transform 1 0 16100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8213
timestamp 1757982896
transform 1 0 17600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8214
timestamp 1757982896
transform 1 0 19100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8215
timestamp 1757982896
transform 1 0 20600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8216
timestamp 1757982896
transform 1 0 22100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8217
timestamp 1757982896
transform 1 0 23600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8218
timestamp 1757982896
transform 1 0 25100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8219
timestamp 1757982896
transform 1 0 26600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8220
timestamp 1757982896
transform 1 0 28100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8221
timestamp 1757982896
transform 1 0 29600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8222
timestamp 1757982896
transform 1 0 31100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8223
timestamp 1757982896
transform 1 0 32600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8224
timestamp 1757982896
transform 1 0 34100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8225
timestamp 1757982896
transform 1 0 35600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8226
timestamp 1757982896
transform 1 0 37100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8227
timestamp 1757982896
transform 1 0 38600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8228
timestamp 1757982896
transform 1 0 40100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8229
timestamp 1757982896
transform 1 0 41600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8230
timestamp 1757982896
transform 1 0 43100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8231
timestamp 1757982896
transform 1 0 44600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8232
timestamp 1757982896
transform 1 0 46100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8233
timestamp 1757982896
transform 1 0 47600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8234
timestamp 1757982896
transform 1 0 49100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8235
timestamp 1757982896
transform 1 0 50600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8236
timestamp 1757982896
transform 1 0 52100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8237
timestamp 1757982896
transform 1 0 53600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8238
timestamp 1757982896
transform 1 0 55100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8239
timestamp 1757982896
transform 1 0 56600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8240
timestamp 1757982896
transform 1 0 58100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8241
timestamp 1757982896
transform 1 0 59600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8242
timestamp 1757982896
transform 1 0 61100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8243
timestamp 1757982896
transform 1 0 62600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8244
timestamp 1757982896
transform 1 0 64100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8245
timestamp 1757982896
transform 1 0 65600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8246
timestamp 1757982896
transform 1 0 67100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8247
timestamp 1757982896
transform 1 0 68600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8248
timestamp 1757982896
transform 1 0 70100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8249
timestamp 1757982896
transform 1 0 71600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8250
timestamp 1757982896
transform 1 0 73100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8251
timestamp 1757982896
transform 1 0 74600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8252
timestamp 1757982896
transform 1 0 76100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8253
timestamp 1757982896
transform 1 0 77600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8254
timestamp 1757982896
transform 1 0 79100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8255
timestamp 1757982896
transform 1 0 80600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8256
timestamp 1757982896
transform 1 0 82100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8257
timestamp 1757982896
transform 1 0 83600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8258
timestamp 1757982896
transform 1 0 85100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8259
timestamp 1757982896
transform 1 0 86600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8260
timestamp 1757982896
transform 1 0 88100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8261
timestamp 1757982896
transform 1 0 89600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8262
timestamp 1757982896
transform 1 0 91100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8263
timestamp 1757982896
transform 1 0 92600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8264
timestamp 1757982896
transform 1 0 94100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8265
timestamp 1757982896
transform 1 0 95600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8266
timestamp 1757982896
transform 1 0 97100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8267
timestamp 1757982896
transform 1 0 98600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8268
timestamp 1757982896
transform 1 0 100100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8269
timestamp 1757982896
transform 1 0 101600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8270
timestamp 1757982896
transform 1 0 103100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8271
timestamp 1757982896
transform 1 0 104600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8272
timestamp 1757982896
transform 1 0 106100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8273
timestamp 1757982896
transform 1 0 107600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8274
timestamp 1757982896
transform 1 0 109100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8275
timestamp 1757982896
transform 1 0 110600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8276
timestamp 1757982896
transform 1 0 112100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8277
timestamp 1757982896
transform 1 0 113600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8278
timestamp 1757982896
transform 1 0 115100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8279
timestamp 1757982896
transform 1 0 116600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8280
timestamp 1757982896
transform 1 0 118100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8281
timestamp 1757982896
transform 1 0 119600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8282
timestamp 1757982896
transform 1 0 121100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8283
timestamp 1757982896
transform 1 0 122600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8284
timestamp 1757982896
transform 1 0 124100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8285
timestamp 1757982896
transform 1 0 125600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8286
timestamp 1757982896
transform 1 0 127100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8287
timestamp 1757982896
transform 1 0 128600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8288
timestamp 1757982896
transform 1 0 130100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8289
timestamp 1757982896
transform 1 0 131600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8290
timestamp 1757982896
transform 1 0 133100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8291
timestamp 1757982896
transform 1 0 134600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8292
timestamp 1757982896
transform 1 0 136100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8293
timestamp 1757982896
transform 1 0 137600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8294
timestamp 1757982896
transform 1 0 139100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8295
timestamp 1757982896
transform 1 0 140600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8296
timestamp 1757982896
transform 1 0 142100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8297
timestamp 1757982896
transform 1 0 143600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8298
timestamp 1757982896
transform 1 0 145100 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8299
timestamp 1757982896
transform 1 0 146600 0 1 -121650
box 1820 -1430 3480 230
use pixel  pixel_8300
timestamp 1757982896
transform 1 0 -1900 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8301
timestamp 1757982896
transform 1 0 -400 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8302
timestamp 1757982896
transform 1 0 1100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8303
timestamp 1757982896
transform 1 0 2600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8304
timestamp 1757982896
transform 1 0 4100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8305
timestamp 1757982896
transform 1 0 5600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8306
timestamp 1757982896
transform 1 0 7100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8307
timestamp 1757982896
transform 1 0 8600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8308
timestamp 1757982896
transform 1 0 10100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8309
timestamp 1757982896
transform 1 0 11600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8310
timestamp 1757982896
transform 1 0 13100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8311
timestamp 1757982896
transform 1 0 14600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8312
timestamp 1757982896
transform 1 0 16100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8313
timestamp 1757982896
transform 1 0 17600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8314
timestamp 1757982896
transform 1 0 19100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8315
timestamp 1757982896
transform 1 0 20600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8316
timestamp 1757982896
transform 1 0 22100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8317
timestamp 1757982896
transform 1 0 23600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8318
timestamp 1757982896
transform 1 0 25100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8319
timestamp 1757982896
transform 1 0 26600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8320
timestamp 1757982896
transform 1 0 28100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8321
timestamp 1757982896
transform 1 0 29600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8322
timestamp 1757982896
transform 1 0 31100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8323
timestamp 1757982896
transform 1 0 32600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8324
timestamp 1757982896
transform 1 0 34100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8325
timestamp 1757982896
transform 1 0 35600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8326
timestamp 1757982896
transform 1 0 37100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8327
timestamp 1757982896
transform 1 0 38600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8328
timestamp 1757982896
transform 1 0 40100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8329
timestamp 1757982896
transform 1 0 41600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8330
timestamp 1757982896
transform 1 0 43100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8331
timestamp 1757982896
transform 1 0 44600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8332
timestamp 1757982896
transform 1 0 46100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8333
timestamp 1757982896
transform 1 0 47600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8334
timestamp 1757982896
transform 1 0 49100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8335
timestamp 1757982896
transform 1 0 50600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8336
timestamp 1757982896
transform 1 0 52100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8337
timestamp 1757982896
transform 1 0 53600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8338
timestamp 1757982896
transform 1 0 55100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8339
timestamp 1757982896
transform 1 0 56600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8340
timestamp 1757982896
transform 1 0 58100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8341
timestamp 1757982896
transform 1 0 59600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8342
timestamp 1757982896
transform 1 0 61100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8343
timestamp 1757982896
transform 1 0 62600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8344
timestamp 1757982896
transform 1 0 64100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8345
timestamp 1757982896
transform 1 0 65600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8346
timestamp 1757982896
transform 1 0 67100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8347
timestamp 1757982896
transform 1 0 68600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8348
timestamp 1757982896
transform 1 0 70100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8349
timestamp 1757982896
transform 1 0 71600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8350
timestamp 1757982896
transform 1 0 73100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8351
timestamp 1757982896
transform 1 0 74600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8352
timestamp 1757982896
transform 1 0 76100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8353
timestamp 1757982896
transform 1 0 77600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8354
timestamp 1757982896
transform 1 0 79100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8355
timestamp 1757982896
transform 1 0 80600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8356
timestamp 1757982896
transform 1 0 82100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8357
timestamp 1757982896
transform 1 0 83600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8358
timestamp 1757982896
transform 1 0 85100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8359
timestamp 1757982896
transform 1 0 86600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8360
timestamp 1757982896
transform 1 0 88100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8361
timestamp 1757982896
transform 1 0 89600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8362
timestamp 1757982896
transform 1 0 91100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8363
timestamp 1757982896
transform 1 0 92600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8364
timestamp 1757982896
transform 1 0 94100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8365
timestamp 1757982896
transform 1 0 95600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8366
timestamp 1757982896
transform 1 0 97100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8367
timestamp 1757982896
transform 1 0 98600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8368
timestamp 1757982896
transform 1 0 100100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8369
timestamp 1757982896
transform 1 0 101600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8370
timestamp 1757982896
transform 1 0 103100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8371
timestamp 1757982896
transform 1 0 104600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8372
timestamp 1757982896
transform 1 0 106100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8373
timestamp 1757982896
transform 1 0 107600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8374
timestamp 1757982896
transform 1 0 109100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8375
timestamp 1757982896
transform 1 0 110600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8376
timestamp 1757982896
transform 1 0 112100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8377
timestamp 1757982896
transform 1 0 113600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8378
timestamp 1757982896
transform 1 0 115100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8379
timestamp 1757982896
transform 1 0 116600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8380
timestamp 1757982896
transform 1 0 118100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8381
timestamp 1757982896
transform 1 0 119600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8382
timestamp 1757982896
transform 1 0 121100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8383
timestamp 1757982896
transform 1 0 122600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8384
timestamp 1757982896
transform 1 0 124100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8385
timestamp 1757982896
transform 1 0 125600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8386
timestamp 1757982896
transform 1 0 127100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8387
timestamp 1757982896
transform 1 0 128600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8388
timestamp 1757982896
transform 1 0 130100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8389
timestamp 1757982896
transform 1 0 131600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8390
timestamp 1757982896
transform 1 0 133100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8391
timestamp 1757982896
transform 1 0 134600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8392
timestamp 1757982896
transform 1 0 136100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8393
timestamp 1757982896
transform 1 0 137600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8394
timestamp 1757982896
transform 1 0 139100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8395
timestamp 1757982896
transform 1 0 140600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8396
timestamp 1757982896
transform 1 0 142100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8397
timestamp 1757982896
transform 1 0 143600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8398
timestamp 1757982896
transform 1 0 145100 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8399
timestamp 1757982896
transform 1 0 146600 0 1 -123150
box 1820 -1430 3480 230
use pixel  pixel_8400
timestamp 1757982896
transform 1 0 -1900 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8401
timestamp 1757982896
transform 1 0 -400 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8402
timestamp 1757982896
transform 1 0 1100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8403
timestamp 1757982896
transform 1 0 2600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8404
timestamp 1757982896
transform 1 0 4100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8405
timestamp 1757982896
transform 1 0 5600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8406
timestamp 1757982896
transform 1 0 7100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8407
timestamp 1757982896
transform 1 0 8600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8408
timestamp 1757982896
transform 1 0 10100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8409
timestamp 1757982896
transform 1 0 11600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8410
timestamp 1757982896
transform 1 0 13100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8411
timestamp 1757982896
transform 1 0 14600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8412
timestamp 1757982896
transform 1 0 16100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8413
timestamp 1757982896
transform 1 0 17600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8414
timestamp 1757982896
transform 1 0 19100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8415
timestamp 1757982896
transform 1 0 20600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8416
timestamp 1757982896
transform 1 0 22100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8417
timestamp 1757982896
transform 1 0 23600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8418
timestamp 1757982896
transform 1 0 25100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8419
timestamp 1757982896
transform 1 0 26600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8420
timestamp 1757982896
transform 1 0 28100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8421
timestamp 1757982896
transform 1 0 29600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8422
timestamp 1757982896
transform 1 0 31100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8423
timestamp 1757982896
transform 1 0 32600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8424
timestamp 1757982896
transform 1 0 34100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8425
timestamp 1757982896
transform 1 0 35600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8426
timestamp 1757982896
transform 1 0 37100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8427
timestamp 1757982896
transform 1 0 38600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8428
timestamp 1757982896
transform 1 0 40100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8429
timestamp 1757982896
transform 1 0 41600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8430
timestamp 1757982896
transform 1 0 43100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8431
timestamp 1757982896
transform 1 0 44600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8432
timestamp 1757982896
transform 1 0 46100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8433
timestamp 1757982896
transform 1 0 47600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8434
timestamp 1757982896
transform 1 0 49100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8435
timestamp 1757982896
transform 1 0 50600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8436
timestamp 1757982896
transform 1 0 52100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8437
timestamp 1757982896
transform 1 0 53600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8438
timestamp 1757982896
transform 1 0 55100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8439
timestamp 1757982896
transform 1 0 56600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8440
timestamp 1757982896
transform 1 0 58100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8441
timestamp 1757982896
transform 1 0 59600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8442
timestamp 1757982896
transform 1 0 61100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8443
timestamp 1757982896
transform 1 0 62600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8444
timestamp 1757982896
transform 1 0 64100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8445
timestamp 1757982896
transform 1 0 65600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8446
timestamp 1757982896
transform 1 0 67100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8447
timestamp 1757982896
transform 1 0 68600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8448
timestamp 1757982896
transform 1 0 70100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8449
timestamp 1757982896
transform 1 0 71600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8450
timestamp 1757982896
transform 1 0 73100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8451
timestamp 1757982896
transform 1 0 74600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8452
timestamp 1757982896
transform 1 0 76100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8453
timestamp 1757982896
transform 1 0 77600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8454
timestamp 1757982896
transform 1 0 79100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8455
timestamp 1757982896
transform 1 0 80600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8456
timestamp 1757982896
transform 1 0 82100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8457
timestamp 1757982896
transform 1 0 83600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8458
timestamp 1757982896
transform 1 0 85100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8459
timestamp 1757982896
transform 1 0 86600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8460
timestamp 1757982896
transform 1 0 88100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8461
timestamp 1757982896
transform 1 0 89600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8462
timestamp 1757982896
transform 1 0 91100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8463
timestamp 1757982896
transform 1 0 92600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8464
timestamp 1757982896
transform 1 0 94100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8465
timestamp 1757982896
transform 1 0 95600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8466
timestamp 1757982896
transform 1 0 97100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8467
timestamp 1757982896
transform 1 0 98600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8468
timestamp 1757982896
transform 1 0 100100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8469
timestamp 1757982896
transform 1 0 101600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8470
timestamp 1757982896
transform 1 0 103100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8471
timestamp 1757982896
transform 1 0 104600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8472
timestamp 1757982896
transform 1 0 106100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8473
timestamp 1757982896
transform 1 0 107600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8474
timestamp 1757982896
transform 1 0 109100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8475
timestamp 1757982896
transform 1 0 110600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8476
timestamp 1757982896
transform 1 0 112100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8477
timestamp 1757982896
transform 1 0 113600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8478
timestamp 1757982896
transform 1 0 115100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8479
timestamp 1757982896
transform 1 0 116600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8480
timestamp 1757982896
transform 1 0 118100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8481
timestamp 1757982896
transform 1 0 119600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8482
timestamp 1757982896
transform 1 0 121100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8483
timestamp 1757982896
transform 1 0 122600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8484
timestamp 1757982896
transform 1 0 124100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8485
timestamp 1757982896
transform 1 0 125600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8486
timestamp 1757982896
transform 1 0 127100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8487
timestamp 1757982896
transform 1 0 128600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8488
timestamp 1757982896
transform 1 0 130100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8489
timestamp 1757982896
transform 1 0 131600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8490
timestamp 1757982896
transform 1 0 133100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8491
timestamp 1757982896
transform 1 0 134600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8492
timestamp 1757982896
transform 1 0 136100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8493
timestamp 1757982896
transform 1 0 137600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8494
timestamp 1757982896
transform 1 0 139100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8495
timestamp 1757982896
transform 1 0 140600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8496
timestamp 1757982896
transform 1 0 142100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8497
timestamp 1757982896
transform 1 0 143600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8498
timestamp 1757982896
transform 1 0 145100 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8499
timestamp 1757982896
transform 1 0 146600 0 1 -124650
box 1820 -1430 3480 230
use pixel  pixel_8500
timestamp 1757982896
transform 1 0 -1900 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8501
timestamp 1757982896
transform 1 0 -400 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8502
timestamp 1757982896
transform 1 0 1100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8503
timestamp 1757982896
transform 1 0 2600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8504
timestamp 1757982896
transform 1 0 4100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8505
timestamp 1757982896
transform 1 0 5600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8506
timestamp 1757982896
transform 1 0 7100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8507
timestamp 1757982896
transform 1 0 8600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8508
timestamp 1757982896
transform 1 0 10100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8509
timestamp 1757982896
transform 1 0 11600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8510
timestamp 1757982896
transform 1 0 13100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8511
timestamp 1757982896
transform 1 0 14600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8512
timestamp 1757982896
transform 1 0 16100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8513
timestamp 1757982896
transform 1 0 17600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8514
timestamp 1757982896
transform 1 0 19100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8515
timestamp 1757982896
transform 1 0 20600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8516
timestamp 1757982896
transform 1 0 22100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8517
timestamp 1757982896
transform 1 0 23600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8518
timestamp 1757982896
transform 1 0 25100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8519
timestamp 1757982896
transform 1 0 26600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8520
timestamp 1757982896
transform 1 0 28100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8521
timestamp 1757982896
transform 1 0 29600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8522
timestamp 1757982896
transform 1 0 31100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8523
timestamp 1757982896
transform 1 0 32600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8524
timestamp 1757982896
transform 1 0 34100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8525
timestamp 1757982896
transform 1 0 35600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8526
timestamp 1757982896
transform 1 0 37100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8527
timestamp 1757982896
transform 1 0 38600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8528
timestamp 1757982896
transform 1 0 40100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8529
timestamp 1757982896
transform 1 0 41600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8530
timestamp 1757982896
transform 1 0 43100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8531
timestamp 1757982896
transform 1 0 44600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8532
timestamp 1757982896
transform 1 0 46100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8533
timestamp 1757982896
transform 1 0 47600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8534
timestamp 1757982896
transform 1 0 49100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8535
timestamp 1757982896
transform 1 0 50600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8536
timestamp 1757982896
transform 1 0 52100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8537
timestamp 1757982896
transform 1 0 53600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8538
timestamp 1757982896
transform 1 0 55100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8539
timestamp 1757982896
transform 1 0 56600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8540
timestamp 1757982896
transform 1 0 58100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8541
timestamp 1757982896
transform 1 0 59600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8542
timestamp 1757982896
transform 1 0 61100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8543
timestamp 1757982896
transform 1 0 62600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8544
timestamp 1757982896
transform 1 0 64100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8545
timestamp 1757982896
transform 1 0 65600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8546
timestamp 1757982896
transform 1 0 67100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8547
timestamp 1757982896
transform 1 0 68600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8548
timestamp 1757982896
transform 1 0 70100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8549
timestamp 1757982896
transform 1 0 71600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8550
timestamp 1757982896
transform 1 0 73100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8551
timestamp 1757982896
transform 1 0 74600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8552
timestamp 1757982896
transform 1 0 76100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8553
timestamp 1757982896
transform 1 0 77600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8554
timestamp 1757982896
transform 1 0 79100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8555
timestamp 1757982896
transform 1 0 80600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8556
timestamp 1757982896
transform 1 0 82100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8557
timestamp 1757982896
transform 1 0 83600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8558
timestamp 1757982896
transform 1 0 85100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8559
timestamp 1757982896
transform 1 0 86600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8560
timestamp 1757982896
transform 1 0 88100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8561
timestamp 1757982896
transform 1 0 89600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8562
timestamp 1757982896
transform 1 0 91100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8563
timestamp 1757982896
transform 1 0 92600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8564
timestamp 1757982896
transform 1 0 94100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8565
timestamp 1757982896
transform 1 0 95600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8566
timestamp 1757982896
transform 1 0 97100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8567
timestamp 1757982896
transform 1 0 98600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8568
timestamp 1757982896
transform 1 0 100100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8569
timestamp 1757982896
transform 1 0 101600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8570
timestamp 1757982896
transform 1 0 103100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8571
timestamp 1757982896
transform 1 0 104600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8572
timestamp 1757982896
transform 1 0 106100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8573
timestamp 1757982896
transform 1 0 107600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8574
timestamp 1757982896
transform 1 0 109100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8575
timestamp 1757982896
transform 1 0 110600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8576
timestamp 1757982896
transform 1 0 112100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8577
timestamp 1757982896
transform 1 0 113600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8578
timestamp 1757982896
transform 1 0 115100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8579
timestamp 1757982896
transform 1 0 116600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8580
timestamp 1757982896
transform 1 0 118100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8581
timestamp 1757982896
transform 1 0 119600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8582
timestamp 1757982896
transform 1 0 121100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8583
timestamp 1757982896
transform 1 0 122600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8584
timestamp 1757982896
transform 1 0 124100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8585
timestamp 1757982896
transform 1 0 125600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8586
timestamp 1757982896
transform 1 0 127100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8587
timestamp 1757982896
transform 1 0 128600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8588
timestamp 1757982896
transform 1 0 130100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8589
timestamp 1757982896
transform 1 0 131600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8590
timestamp 1757982896
transform 1 0 133100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8591
timestamp 1757982896
transform 1 0 134600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8592
timestamp 1757982896
transform 1 0 136100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8593
timestamp 1757982896
transform 1 0 137600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8594
timestamp 1757982896
transform 1 0 139100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8595
timestamp 1757982896
transform 1 0 140600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8596
timestamp 1757982896
transform 1 0 142100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8597
timestamp 1757982896
transform 1 0 143600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8598
timestamp 1757982896
transform 1 0 145100 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8599
timestamp 1757982896
transform 1 0 146600 0 1 -126150
box 1820 -1430 3480 230
use pixel  pixel_8600
timestamp 1757982896
transform 1 0 -1900 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8601
timestamp 1757982896
transform 1 0 -400 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8602
timestamp 1757982896
transform 1 0 1100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8603
timestamp 1757982896
transform 1 0 2600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8604
timestamp 1757982896
transform 1 0 4100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8605
timestamp 1757982896
transform 1 0 5600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8606
timestamp 1757982896
transform 1 0 7100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8607
timestamp 1757982896
transform 1 0 8600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8608
timestamp 1757982896
transform 1 0 10100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8609
timestamp 1757982896
transform 1 0 11600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8610
timestamp 1757982896
transform 1 0 13100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8611
timestamp 1757982896
transform 1 0 14600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8612
timestamp 1757982896
transform 1 0 16100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8613
timestamp 1757982896
transform 1 0 17600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8614
timestamp 1757982896
transform 1 0 19100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8615
timestamp 1757982896
transform 1 0 20600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8616
timestamp 1757982896
transform 1 0 22100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8617
timestamp 1757982896
transform 1 0 23600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8618
timestamp 1757982896
transform 1 0 25100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8619
timestamp 1757982896
transform 1 0 26600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8620
timestamp 1757982896
transform 1 0 28100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8621
timestamp 1757982896
transform 1 0 29600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8622
timestamp 1757982896
transform 1 0 31100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8623
timestamp 1757982896
transform 1 0 32600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8624
timestamp 1757982896
transform 1 0 34100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8625
timestamp 1757982896
transform 1 0 35600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8626
timestamp 1757982896
transform 1 0 37100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8627
timestamp 1757982896
transform 1 0 38600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8628
timestamp 1757982896
transform 1 0 40100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8629
timestamp 1757982896
transform 1 0 41600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8630
timestamp 1757982896
transform 1 0 43100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8631
timestamp 1757982896
transform 1 0 44600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8632
timestamp 1757982896
transform 1 0 46100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8633
timestamp 1757982896
transform 1 0 47600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8634
timestamp 1757982896
transform 1 0 49100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8635
timestamp 1757982896
transform 1 0 50600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8636
timestamp 1757982896
transform 1 0 52100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8637
timestamp 1757982896
transform 1 0 53600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8638
timestamp 1757982896
transform 1 0 55100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8639
timestamp 1757982896
transform 1 0 56600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8640
timestamp 1757982896
transform 1 0 58100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8641
timestamp 1757982896
transform 1 0 59600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8642
timestamp 1757982896
transform 1 0 61100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8643
timestamp 1757982896
transform 1 0 62600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8644
timestamp 1757982896
transform 1 0 64100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8645
timestamp 1757982896
transform 1 0 65600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8646
timestamp 1757982896
transform 1 0 67100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8647
timestamp 1757982896
transform 1 0 68600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8648
timestamp 1757982896
transform 1 0 70100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8649
timestamp 1757982896
transform 1 0 71600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8650
timestamp 1757982896
transform 1 0 73100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8651
timestamp 1757982896
transform 1 0 74600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8652
timestamp 1757982896
transform 1 0 76100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8653
timestamp 1757982896
transform 1 0 77600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8654
timestamp 1757982896
transform 1 0 79100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8655
timestamp 1757982896
transform 1 0 80600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8656
timestamp 1757982896
transform 1 0 82100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8657
timestamp 1757982896
transform 1 0 83600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8658
timestamp 1757982896
transform 1 0 85100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8659
timestamp 1757982896
transform 1 0 86600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8660
timestamp 1757982896
transform 1 0 88100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8661
timestamp 1757982896
transform 1 0 89600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8662
timestamp 1757982896
transform 1 0 91100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8663
timestamp 1757982896
transform 1 0 92600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8664
timestamp 1757982896
transform 1 0 94100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8665
timestamp 1757982896
transform 1 0 95600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8666
timestamp 1757982896
transform 1 0 97100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8667
timestamp 1757982896
transform 1 0 98600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8668
timestamp 1757982896
transform 1 0 100100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8669
timestamp 1757982896
transform 1 0 101600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8670
timestamp 1757982896
transform 1 0 103100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8671
timestamp 1757982896
transform 1 0 104600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8672
timestamp 1757982896
transform 1 0 106100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8673
timestamp 1757982896
transform 1 0 107600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8674
timestamp 1757982896
transform 1 0 109100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8675
timestamp 1757982896
transform 1 0 110600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8676
timestamp 1757982896
transform 1 0 112100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8677
timestamp 1757982896
transform 1 0 113600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8678
timestamp 1757982896
transform 1 0 115100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8679
timestamp 1757982896
transform 1 0 116600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8680
timestamp 1757982896
transform 1 0 118100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8681
timestamp 1757982896
transform 1 0 119600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8682
timestamp 1757982896
transform 1 0 121100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8683
timestamp 1757982896
transform 1 0 122600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8684
timestamp 1757982896
transform 1 0 124100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8685
timestamp 1757982896
transform 1 0 125600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8686
timestamp 1757982896
transform 1 0 127100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8687
timestamp 1757982896
transform 1 0 128600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8688
timestamp 1757982896
transform 1 0 130100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8689
timestamp 1757982896
transform 1 0 131600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8690
timestamp 1757982896
transform 1 0 133100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8691
timestamp 1757982896
transform 1 0 134600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8692
timestamp 1757982896
transform 1 0 136100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8693
timestamp 1757982896
transform 1 0 137600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8694
timestamp 1757982896
transform 1 0 139100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8695
timestamp 1757982896
transform 1 0 140600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8696
timestamp 1757982896
transform 1 0 142100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8697
timestamp 1757982896
transform 1 0 143600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8698
timestamp 1757982896
transform 1 0 145100 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8699
timestamp 1757982896
transform 1 0 146600 0 1 -127650
box 1820 -1430 3480 230
use pixel  pixel_8700
timestamp 1757982896
transform 1 0 -1900 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8701
timestamp 1757982896
transform 1 0 -400 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8702
timestamp 1757982896
transform 1 0 1100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8703
timestamp 1757982896
transform 1 0 2600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8704
timestamp 1757982896
transform 1 0 4100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8705
timestamp 1757982896
transform 1 0 5600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8706
timestamp 1757982896
transform 1 0 7100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8707
timestamp 1757982896
transform 1 0 8600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8708
timestamp 1757982896
transform 1 0 10100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8709
timestamp 1757982896
transform 1 0 11600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8710
timestamp 1757982896
transform 1 0 13100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8711
timestamp 1757982896
transform 1 0 14600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8712
timestamp 1757982896
transform 1 0 16100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8713
timestamp 1757982896
transform 1 0 17600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8714
timestamp 1757982896
transform 1 0 19100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8715
timestamp 1757982896
transform 1 0 20600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8716
timestamp 1757982896
transform 1 0 22100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8717
timestamp 1757982896
transform 1 0 23600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8718
timestamp 1757982896
transform 1 0 25100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8719
timestamp 1757982896
transform 1 0 26600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8720
timestamp 1757982896
transform 1 0 28100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8721
timestamp 1757982896
transform 1 0 29600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8722
timestamp 1757982896
transform 1 0 31100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8723
timestamp 1757982896
transform 1 0 32600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8724
timestamp 1757982896
transform 1 0 34100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8725
timestamp 1757982896
transform 1 0 35600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8726
timestamp 1757982896
transform 1 0 37100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8727
timestamp 1757982896
transform 1 0 38600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8728
timestamp 1757982896
transform 1 0 40100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8729
timestamp 1757982896
transform 1 0 41600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8730
timestamp 1757982896
transform 1 0 43100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8731
timestamp 1757982896
transform 1 0 44600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8732
timestamp 1757982896
transform 1 0 46100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8733
timestamp 1757982896
transform 1 0 47600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8734
timestamp 1757982896
transform 1 0 49100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8735
timestamp 1757982896
transform 1 0 50600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8736
timestamp 1757982896
transform 1 0 52100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8737
timestamp 1757982896
transform 1 0 53600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8738
timestamp 1757982896
transform 1 0 55100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8739
timestamp 1757982896
transform 1 0 56600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8740
timestamp 1757982896
transform 1 0 58100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8741
timestamp 1757982896
transform 1 0 59600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8742
timestamp 1757982896
transform 1 0 61100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8743
timestamp 1757982896
transform 1 0 62600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8744
timestamp 1757982896
transform 1 0 64100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8745
timestamp 1757982896
transform 1 0 65600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8746
timestamp 1757982896
transform 1 0 67100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8747
timestamp 1757982896
transform 1 0 68600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8748
timestamp 1757982896
transform 1 0 70100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8749
timestamp 1757982896
transform 1 0 71600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8750
timestamp 1757982896
transform 1 0 73100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8751
timestamp 1757982896
transform 1 0 74600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8752
timestamp 1757982896
transform 1 0 76100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8753
timestamp 1757982896
transform 1 0 77600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8754
timestamp 1757982896
transform 1 0 79100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8755
timestamp 1757982896
transform 1 0 80600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8756
timestamp 1757982896
transform 1 0 82100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8757
timestamp 1757982896
transform 1 0 83600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8758
timestamp 1757982896
transform 1 0 85100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8759
timestamp 1757982896
transform 1 0 86600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8760
timestamp 1757982896
transform 1 0 88100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8761
timestamp 1757982896
transform 1 0 89600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8762
timestamp 1757982896
transform 1 0 91100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8763
timestamp 1757982896
transform 1 0 92600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8764
timestamp 1757982896
transform 1 0 94100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8765
timestamp 1757982896
transform 1 0 95600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8766
timestamp 1757982896
transform 1 0 97100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8767
timestamp 1757982896
transform 1 0 98600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8768
timestamp 1757982896
transform 1 0 100100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8769
timestamp 1757982896
transform 1 0 101600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8770
timestamp 1757982896
transform 1 0 103100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8771
timestamp 1757982896
transform 1 0 104600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8772
timestamp 1757982896
transform 1 0 106100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8773
timestamp 1757982896
transform 1 0 107600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8774
timestamp 1757982896
transform 1 0 109100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8775
timestamp 1757982896
transform 1 0 110600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8776
timestamp 1757982896
transform 1 0 112100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8777
timestamp 1757982896
transform 1 0 113600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8778
timestamp 1757982896
transform 1 0 115100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8779
timestamp 1757982896
transform 1 0 116600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8780
timestamp 1757982896
transform 1 0 118100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8781
timestamp 1757982896
transform 1 0 119600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8782
timestamp 1757982896
transform 1 0 121100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8783
timestamp 1757982896
transform 1 0 122600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8784
timestamp 1757982896
transform 1 0 124100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8785
timestamp 1757982896
transform 1 0 125600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8786
timestamp 1757982896
transform 1 0 127100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8787
timestamp 1757982896
transform 1 0 128600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8788
timestamp 1757982896
transform 1 0 130100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8789
timestamp 1757982896
transform 1 0 131600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8790
timestamp 1757982896
transform 1 0 133100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8791
timestamp 1757982896
transform 1 0 134600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8792
timestamp 1757982896
transform 1 0 136100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8793
timestamp 1757982896
transform 1 0 137600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8794
timestamp 1757982896
transform 1 0 139100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8795
timestamp 1757982896
transform 1 0 140600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8796
timestamp 1757982896
transform 1 0 142100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8797
timestamp 1757982896
transform 1 0 143600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8798
timestamp 1757982896
transform 1 0 145100 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8799
timestamp 1757982896
transform 1 0 146600 0 1 -129150
box 1820 -1430 3480 230
use pixel  pixel_8800
timestamp 1757982896
transform 1 0 -1900 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8801
timestamp 1757982896
transform 1 0 -400 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8802
timestamp 1757982896
transform 1 0 1100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8803
timestamp 1757982896
transform 1 0 2600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8804
timestamp 1757982896
transform 1 0 4100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8805
timestamp 1757982896
transform 1 0 5600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8806
timestamp 1757982896
transform 1 0 7100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8807
timestamp 1757982896
transform 1 0 8600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8808
timestamp 1757982896
transform 1 0 10100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8809
timestamp 1757982896
transform 1 0 11600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8810
timestamp 1757982896
transform 1 0 13100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8811
timestamp 1757982896
transform 1 0 14600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8812
timestamp 1757982896
transform 1 0 16100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8813
timestamp 1757982896
transform 1 0 17600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8814
timestamp 1757982896
transform 1 0 19100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8815
timestamp 1757982896
transform 1 0 20600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8816
timestamp 1757982896
transform 1 0 22100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8817
timestamp 1757982896
transform 1 0 23600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8818
timestamp 1757982896
transform 1 0 25100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8819
timestamp 1757982896
transform 1 0 26600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8820
timestamp 1757982896
transform 1 0 28100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8821
timestamp 1757982896
transform 1 0 29600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8822
timestamp 1757982896
transform 1 0 31100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8823
timestamp 1757982896
transform 1 0 32600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8824
timestamp 1757982896
transform 1 0 34100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8825
timestamp 1757982896
transform 1 0 35600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8826
timestamp 1757982896
transform 1 0 37100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8827
timestamp 1757982896
transform 1 0 38600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8828
timestamp 1757982896
transform 1 0 40100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8829
timestamp 1757982896
transform 1 0 41600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8830
timestamp 1757982896
transform 1 0 43100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8831
timestamp 1757982896
transform 1 0 44600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8832
timestamp 1757982896
transform 1 0 46100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8833
timestamp 1757982896
transform 1 0 47600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8834
timestamp 1757982896
transform 1 0 49100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8835
timestamp 1757982896
transform 1 0 50600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8836
timestamp 1757982896
transform 1 0 52100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8837
timestamp 1757982896
transform 1 0 53600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8838
timestamp 1757982896
transform 1 0 55100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8839
timestamp 1757982896
transform 1 0 56600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8840
timestamp 1757982896
transform 1 0 58100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8841
timestamp 1757982896
transform 1 0 59600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8842
timestamp 1757982896
transform 1 0 61100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8843
timestamp 1757982896
transform 1 0 62600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8844
timestamp 1757982896
transform 1 0 64100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8845
timestamp 1757982896
transform 1 0 65600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8846
timestamp 1757982896
transform 1 0 67100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8847
timestamp 1757982896
transform 1 0 68600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8848
timestamp 1757982896
transform 1 0 70100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8849
timestamp 1757982896
transform 1 0 71600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8850
timestamp 1757982896
transform 1 0 73100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8851
timestamp 1757982896
transform 1 0 74600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8852
timestamp 1757982896
transform 1 0 76100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8853
timestamp 1757982896
transform 1 0 77600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8854
timestamp 1757982896
transform 1 0 79100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8855
timestamp 1757982896
transform 1 0 80600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8856
timestamp 1757982896
transform 1 0 82100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8857
timestamp 1757982896
transform 1 0 83600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8858
timestamp 1757982896
transform 1 0 85100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8859
timestamp 1757982896
transform 1 0 86600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8860
timestamp 1757982896
transform 1 0 88100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8861
timestamp 1757982896
transform 1 0 89600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8862
timestamp 1757982896
transform 1 0 91100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8863
timestamp 1757982896
transform 1 0 92600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8864
timestamp 1757982896
transform 1 0 94100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8865
timestamp 1757982896
transform 1 0 95600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8866
timestamp 1757982896
transform 1 0 97100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8867
timestamp 1757982896
transform 1 0 98600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8868
timestamp 1757982896
transform 1 0 100100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8869
timestamp 1757982896
transform 1 0 101600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8870
timestamp 1757982896
transform 1 0 103100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8871
timestamp 1757982896
transform 1 0 104600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8872
timestamp 1757982896
transform 1 0 106100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8873
timestamp 1757982896
transform 1 0 107600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8874
timestamp 1757982896
transform 1 0 109100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8875
timestamp 1757982896
transform 1 0 110600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8876
timestamp 1757982896
transform 1 0 112100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8877
timestamp 1757982896
transform 1 0 113600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8878
timestamp 1757982896
transform 1 0 115100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8879
timestamp 1757982896
transform 1 0 116600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8880
timestamp 1757982896
transform 1 0 118100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8881
timestamp 1757982896
transform 1 0 119600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8882
timestamp 1757982896
transform 1 0 121100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8883
timestamp 1757982896
transform 1 0 122600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8884
timestamp 1757982896
transform 1 0 124100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8885
timestamp 1757982896
transform 1 0 125600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8886
timestamp 1757982896
transform 1 0 127100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8887
timestamp 1757982896
transform 1 0 128600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8888
timestamp 1757982896
transform 1 0 130100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8889
timestamp 1757982896
transform 1 0 131600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8890
timestamp 1757982896
transform 1 0 133100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8891
timestamp 1757982896
transform 1 0 134600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8892
timestamp 1757982896
transform 1 0 136100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8893
timestamp 1757982896
transform 1 0 137600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8894
timestamp 1757982896
transform 1 0 139100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8895
timestamp 1757982896
transform 1 0 140600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8896
timestamp 1757982896
transform 1 0 142100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8897
timestamp 1757982896
transform 1 0 143600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8898
timestamp 1757982896
transform 1 0 145100 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8899
timestamp 1757982896
transform 1 0 146600 0 1 -130650
box 1820 -1430 3480 230
use pixel  pixel_8900
timestamp 1757982896
transform 1 0 -1900 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8901
timestamp 1757982896
transform 1 0 -400 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8902
timestamp 1757982896
transform 1 0 1100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8903
timestamp 1757982896
transform 1 0 2600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8904
timestamp 1757982896
transform 1 0 4100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8905
timestamp 1757982896
transform 1 0 5600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8906
timestamp 1757982896
transform 1 0 7100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8907
timestamp 1757982896
transform 1 0 8600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8908
timestamp 1757982896
transform 1 0 10100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8909
timestamp 1757982896
transform 1 0 11600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8910
timestamp 1757982896
transform 1 0 13100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8911
timestamp 1757982896
transform 1 0 14600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8912
timestamp 1757982896
transform 1 0 16100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8913
timestamp 1757982896
transform 1 0 17600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8914
timestamp 1757982896
transform 1 0 19100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8915
timestamp 1757982896
transform 1 0 20600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8916
timestamp 1757982896
transform 1 0 22100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8917
timestamp 1757982896
transform 1 0 23600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8918
timestamp 1757982896
transform 1 0 25100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8919
timestamp 1757982896
transform 1 0 26600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8920
timestamp 1757982896
transform 1 0 28100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8921
timestamp 1757982896
transform 1 0 29600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8922
timestamp 1757982896
transform 1 0 31100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8923
timestamp 1757982896
transform 1 0 32600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8924
timestamp 1757982896
transform 1 0 34100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8925
timestamp 1757982896
transform 1 0 35600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8926
timestamp 1757982896
transform 1 0 37100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8927
timestamp 1757982896
transform 1 0 38600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8928
timestamp 1757982896
transform 1 0 40100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8929
timestamp 1757982896
transform 1 0 41600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8930
timestamp 1757982896
transform 1 0 43100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8931
timestamp 1757982896
transform 1 0 44600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8932
timestamp 1757982896
transform 1 0 46100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8933
timestamp 1757982896
transform 1 0 47600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8934
timestamp 1757982896
transform 1 0 49100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8935
timestamp 1757982896
transform 1 0 50600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8936
timestamp 1757982896
transform 1 0 52100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8937
timestamp 1757982896
transform 1 0 53600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8938
timestamp 1757982896
transform 1 0 55100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8939
timestamp 1757982896
transform 1 0 56600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8940
timestamp 1757982896
transform 1 0 58100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8941
timestamp 1757982896
transform 1 0 59600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8942
timestamp 1757982896
transform 1 0 61100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8943
timestamp 1757982896
transform 1 0 62600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8944
timestamp 1757982896
transform 1 0 64100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8945
timestamp 1757982896
transform 1 0 65600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8946
timestamp 1757982896
transform 1 0 67100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8947
timestamp 1757982896
transform 1 0 68600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8948
timestamp 1757982896
transform 1 0 70100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8949
timestamp 1757982896
transform 1 0 71600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8950
timestamp 1757982896
transform 1 0 73100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8951
timestamp 1757982896
transform 1 0 74600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8952
timestamp 1757982896
transform 1 0 76100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8953
timestamp 1757982896
transform 1 0 77600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8954
timestamp 1757982896
transform 1 0 79100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8955
timestamp 1757982896
transform 1 0 80600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8956
timestamp 1757982896
transform 1 0 82100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8957
timestamp 1757982896
transform 1 0 83600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8958
timestamp 1757982896
transform 1 0 85100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8959
timestamp 1757982896
transform 1 0 86600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8960
timestamp 1757982896
transform 1 0 88100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8961
timestamp 1757982896
transform 1 0 89600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8962
timestamp 1757982896
transform 1 0 91100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8963
timestamp 1757982896
transform 1 0 92600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8964
timestamp 1757982896
transform 1 0 94100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8965
timestamp 1757982896
transform 1 0 95600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8966
timestamp 1757982896
transform 1 0 97100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8967
timestamp 1757982896
transform 1 0 98600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8968
timestamp 1757982896
transform 1 0 100100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8969
timestamp 1757982896
transform 1 0 101600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8970
timestamp 1757982896
transform 1 0 103100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8971
timestamp 1757982896
transform 1 0 104600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8972
timestamp 1757982896
transform 1 0 106100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8973
timestamp 1757982896
transform 1 0 107600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8974
timestamp 1757982896
transform 1 0 109100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8975
timestamp 1757982896
transform 1 0 110600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8976
timestamp 1757982896
transform 1 0 112100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8977
timestamp 1757982896
transform 1 0 113600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8978
timestamp 1757982896
transform 1 0 115100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8979
timestamp 1757982896
transform 1 0 116600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8980
timestamp 1757982896
transform 1 0 118100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8981
timestamp 1757982896
transform 1 0 119600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8982
timestamp 1757982896
transform 1 0 121100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8983
timestamp 1757982896
transform 1 0 122600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8984
timestamp 1757982896
transform 1 0 124100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8985
timestamp 1757982896
transform 1 0 125600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8986
timestamp 1757982896
transform 1 0 127100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8987
timestamp 1757982896
transform 1 0 128600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8988
timestamp 1757982896
transform 1 0 130100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8989
timestamp 1757982896
transform 1 0 131600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8990
timestamp 1757982896
transform 1 0 133100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8991
timestamp 1757982896
transform 1 0 134600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8992
timestamp 1757982896
transform 1 0 136100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8993
timestamp 1757982896
transform 1 0 137600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8994
timestamp 1757982896
transform 1 0 139100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8995
timestamp 1757982896
transform 1 0 140600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8996
timestamp 1757982896
transform 1 0 142100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8997
timestamp 1757982896
transform 1 0 143600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8998
timestamp 1757982896
transform 1 0 145100 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_8999
timestamp 1757982896
transform 1 0 146600 0 1 -132150
box 1820 -1430 3480 230
use pixel  pixel_9000
timestamp 1757982896
transform 1 0 -1900 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9001
timestamp 1757982896
transform 1 0 -400 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9002
timestamp 1757982896
transform 1 0 1100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9003
timestamp 1757982896
transform 1 0 2600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9004
timestamp 1757982896
transform 1 0 4100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9005
timestamp 1757982896
transform 1 0 5600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9006
timestamp 1757982896
transform 1 0 7100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9007
timestamp 1757982896
transform 1 0 8600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9008
timestamp 1757982896
transform 1 0 10100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9009
timestamp 1757982896
transform 1 0 11600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9010
timestamp 1757982896
transform 1 0 13100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9011
timestamp 1757982896
transform 1 0 14600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9012
timestamp 1757982896
transform 1 0 16100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9013
timestamp 1757982896
transform 1 0 17600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9014
timestamp 1757982896
transform 1 0 19100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9015
timestamp 1757982896
transform 1 0 20600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9016
timestamp 1757982896
transform 1 0 22100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9017
timestamp 1757982896
transform 1 0 23600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9018
timestamp 1757982896
transform 1 0 25100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9019
timestamp 1757982896
transform 1 0 26600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9020
timestamp 1757982896
transform 1 0 28100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9021
timestamp 1757982896
transform 1 0 29600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9022
timestamp 1757982896
transform 1 0 31100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9023
timestamp 1757982896
transform 1 0 32600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9024
timestamp 1757982896
transform 1 0 34100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9025
timestamp 1757982896
transform 1 0 35600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9026
timestamp 1757982896
transform 1 0 37100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9027
timestamp 1757982896
transform 1 0 38600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9028
timestamp 1757982896
transform 1 0 40100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9029
timestamp 1757982896
transform 1 0 41600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9030
timestamp 1757982896
transform 1 0 43100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9031
timestamp 1757982896
transform 1 0 44600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9032
timestamp 1757982896
transform 1 0 46100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9033
timestamp 1757982896
transform 1 0 47600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9034
timestamp 1757982896
transform 1 0 49100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9035
timestamp 1757982896
transform 1 0 50600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9036
timestamp 1757982896
transform 1 0 52100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9037
timestamp 1757982896
transform 1 0 53600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9038
timestamp 1757982896
transform 1 0 55100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9039
timestamp 1757982896
transform 1 0 56600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9040
timestamp 1757982896
transform 1 0 58100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9041
timestamp 1757982896
transform 1 0 59600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9042
timestamp 1757982896
transform 1 0 61100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9043
timestamp 1757982896
transform 1 0 62600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9044
timestamp 1757982896
transform 1 0 64100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9045
timestamp 1757982896
transform 1 0 65600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9046
timestamp 1757982896
transform 1 0 67100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9047
timestamp 1757982896
transform 1 0 68600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9048
timestamp 1757982896
transform 1 0 70100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9049
timestamp 1757982896
transform 1 0 71600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9050
timestamp 1757982896
transform 1 0 73100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9051
timestamp 1757982896
transform 1 0 74600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9052
timestamp 1757982896
transform 1 0 76100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9053
timestamp 1757982896
transform 1 0 77600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9054
timestamp 1757982896
transform 1 0 79100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9055
timestamp 1757982896
transform 1 0 80600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9056
timestamp 1757982896
transform 1 0 82100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9057
timestamp 1757982896
transform 1 0 83600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9058
timestamp 1757982896
transform 1 0 85100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9059
timestamp 1757982896
transform 1 0 86600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9060
timestamp 1757982896
transform 1 0 88100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9061
timestamp 1757982896
transform 1 0 89600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9062
timestamp 1757982896
transform 1 0 91100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9063
timestamp 1757982896
transform 1 0 92600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9064
timestamp 1757982896
transform 1 0 94100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9065
timestamp 1757982896
transform 1 0 95600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9066
timestamp 1757982896
transform 1 0 97100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9067
timestamp 1757982896
transform 1 0 98600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9068
timestamp 1757982896
transform 1 0 100100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9069
timestamp 1757982896
transform 1 0 101600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9070
timestamp 1757982896
transform 1 0 103100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9071
timestamp 1757982896
transform 1 0 104600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9072
timestamp 1757982896
transform 1 0 106100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9073
timestamp 1757982896
transform 1 0 107600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9074
timestamp 1757982896
transform 1 0 109100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9075
timestamp 1757982896
transform 1 0 110600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9076
timestamp 1757982896
transform 1 0 112100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9077
timestamp 1757982896
transform 1 0 113600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9078
timestamp 1757982896
transform 1 0 115100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9079
timestamp 1757982896
transform 1 0 116600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9080
timestamp 1757982896
transform 1 0 118100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9081
timestamp 1757982896
transform 1 0 119600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9082
timestamp 1757982896
transform 1 0 121100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9083
timestamp 1757982896
transform 1 0 122600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9084
timestamp 1757982896
transform 1 0 124100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9085
timestamp 1757982896
transform 1 0 125600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9086
timestamp 1757982896
transform 1 0 127100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9087
timestamp 1757982896
transform 1 0 128600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9088
timestamp 1757982896
transform 1 0 130100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9089
timestamp 1757982896
transform 1 0 131600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9090
timestamp 1757982896
transform 1 0 133100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9091
timestamp 1757982896
transform 1 0 134600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9092
timestamp 1757982896
transform 1 0 136100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9093
timestamp 1757982896
transform 1 0 137600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9094
timestamp 1757982896
transform 1 0 139100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9095
timestamp 1757982896
transform 1 0 140600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9096
timestamp 1757982896
transform 1 0 142100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9097
timestamp 1757982896
transform 1 0 143600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9098
timestamp 1757982896
transform 1 0 145100 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9099
timestamp 1757982896
transform 1 0 146600 0 1 -133650
box 1820 -1430 3480 230
use pixel  pixel_9100
timestamp 1757982896
transform 1 0 -1900 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9101
timestamp 1757982896
transform 1 0 -400 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9102
timestamp 1757982896
transform 1 0 1100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9103
timestamp 1757982896
transform 1 0 2600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9104
timestamp 1757982896
transform 1 0 4100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9105
timestamp 1757982896
transform 1 0 5600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9106
timestamp 1757982896
transform 1 0 7100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9107
timestamp 1757982896
transform 1 0 8600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9108
timestamp 1757982896
transform 1 0 10100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9109
timestamp 1757982896
transform 1 0 11600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9110
timestamp 1757982896
transform 1 0 13100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9111
timestamp 1757982896
transform 1 0 14600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9112
timestamp 1757982896
transform 1 0 16100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9113
timestamp 1757982896
transform 1 0 17600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9114
timestamp 1757982896
transform 1 0 19100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9115
timestamp 1757982896
transform 1 0 20600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9116
timestamp 1757982896
transform 1 0 22100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9117
timestamp 1757982896
transform 1 0 23600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9118
timestamp 1757982896
transform 1 0 25100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9119
timestamp 1757982896
transform 1 0 26600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9120
timestamp 1757982896
transform 1 0 28100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9121
timestamp 1757982896
transform 1 0 29600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9122
timestamp 1757982896
transform 1 0 31100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9123
timestamp 1757982896
transform 1 0 32600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9124
timestamp 1757982896
transform 1 0 34100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9125
timestamp 1757982896
transform 1 0 35600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9126
timestamp 1757982896
transform 1 0 37100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9127
timestamp 1757982896
transform 1 0 38600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9128
timestamp 1757982896
transform 1 0 40100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9129
timestamp 1757982896
transform 1 0 41600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9130
timestamp 1757982896
transform 1 0 43100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9131
timestamp 1757982896
transform 1 0 44600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9132
timestamp 1757982896
transform 1 0 46100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9133
timestamp 1757982896
transform 1 0 47600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9134
timestamp 1757982896
transform 1 0 49100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9135
timestamp 1757982896
transform 1 0 50600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9136
timestamp 1757982896
transform 1 0 52100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9137
timestamp 1757982896
transform 1 0 53600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9138
timestamp 1757982896
transform 1 0 55100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9139
timestamp 1757982896
transform 1 0 56600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9140
timestamp 1757982896
transform 1 0 58100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9141
timestamp 1757982896
transform 1 0 59600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9142
timestamp 1757982896
transform 1 0 61100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9143
timestamp 1757982896
transform 1 0 62600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9144
timestamp 1757982896
transform 1 0 64100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9145
timestamp 1757982896
transform 1 0 65600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9146
timestamp 1757982896
transform 1 0 67100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9147
timestamp 1757982896
transform 1 0 68600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9148
timestamp 1757982896
transform 1 0 70100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9149
timestamp 1757982896
transform 1 0 71600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9150
timestamp 1757982896
transform 1 0 73100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9151
timestamp 1757982896
transform 1 0 74600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9152
timestamp 1757982896
transform 1 0 76100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9153
timestamp 1757982896
transform 1 0 77600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9154
timestamp 1757982896
transform 1 0 79100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9155
timestamp 1757982896
transform 1 0 80600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9156
timestamp 1757982896
transform 1 0 82100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9157
timestamp 1757982896
transform 1 0 83600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9158
timestamp 1757982896
transform 1 0 85100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9159
timestamp 1757982896
transform 1 0 86600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9160
timestamp 1757982896
transform 1 0 88100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9161
timestamp 1757982896
transform 1 0 89600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9162
timestamp 1757982896
transform 1 0 91100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9163
timestamp 1757982896
transform 1 0 92600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9164
timestamp 1757982896
transform 1 0 94100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9165
timestamp 1757982896
transform 1 0 95600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9166
timestamp 1757982896
transform 1 0 97100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9167
timestamp 1757982896
transform 1 0 98600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9168
timestamp 1757982896
transform 1 0 100100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9169
timestamp 1757982896
transform 1 0 101600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9170
timestamp 1757982896
transform 1 0 103100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9171
timestamp 1757982896
transform 1 0 104600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9172
timestamp 1757982896
transform 1 0 106100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9173
timestamp 1757982896
transform 1 0 107600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9174
timestamp 1757982896
transform 1 0 109100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9175
timestamp 1757982896
transform 1 0 110600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9176
timestamp 1757982896
transform 1 0 112100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9177
timestamp 1757982896
transform 1 0 113600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9178
timestamp 1757982896
transform 1 0 115100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9179
timestamp 1757982896
transform 1 0 116600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9180
timestamp 1757982896
transform 1 0 118100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9181
timestamp 1757982896
transform 1 0 119600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9182
timestamp 1757982896
transform 1 0 121100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9183
timestamp 1757982896
transform 1 0 122600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9184
timestamp 1757982896
transform 1 0 124100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9185
timestamp 1757982896
transform 1 0 125600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9186
timestamp 1757982896
transform 1 0 127100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9187
timestamp 1757982896
transform 1 0 128600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9188
timestamp 1757982896
transform 1 0 130100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9189
timestamp 1757982896
transform 1 0 131600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9190
timestamp 1757982896
transform 1 0 133100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9191
timestamp 1757982896
transform 1 0 134600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9192
timestamp 1757982896
transform 1 0 136100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9193
timestamp 1757982896
transform 1 0 137600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9194
timestamp 1757982896
transform 1 0 139100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9195
timestamp 1757982896
transform 1 0 140600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9196
timestamp 1757982896
transform 1 0 142100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9197
timestamp 1757982896
transform 1 0 143600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9198
timestamp 1757982896
transform 1 0 145100 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9199
timestamp 1757982896
transform 1 0 146600 0 1 -135150
box 1820 -1430 3480 230
use pixel  pixel_9200
timestamp 1757982896
transform 1 0 -1900 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9201
timestamp 1757982896
transform 1 0 -400 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9202
timestamp 1757982896
transform 1 0 1100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9203
timestamp 1757982896
transform 1 0 2600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9204
timestamp 1757982896
transform 1 0 4100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9205
timestamp 1757982896
transform 1 0 5600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9206
timestamp 1757982896
transform 1 0 7100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9207
timestamp 1757982896
transform 1 0 8600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9208
timestamp 1757982896
transform 1 0 10100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9209
timestamp 1757982896
transform 1 0 11600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9210
timestamp 1757982896
transform 1 0 13100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9211
timestamp 1757982896
transform 1 0 14600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9212
timestamp 1757982896
transform 1 0 16100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9213
timestamp 1757982896
transform 1 0 17600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9214
timestamp 1757982896
transform 1 0 19100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9215
timestamp 1757982896
transform 1 0 20600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9216
timestamp 1757982896
transform 1 0 22100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9217
timestamp 1757982896
transform 1 0 23600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9218
timestamp 1757982896
transform 1 0 25100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9219
timestamp 1757982896
transform 1 0 26600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9220
timestamp 1757982896
transform 1 0 28100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9221
timestamp 1757982896
transform 1 0 29600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9222
timestamp 1757982896
transform 1 0 31100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9223
timestamp 1757982896
transform 1 0 32600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9224
timestamp 1757982896
transform 1 0 34100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9225
timestamp 1757982896
transform 1 0 35600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9226
timestamp 1757982896
transform 1 0 37100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9227
timestamp 1757982896
transform 1 0 38600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9228
timestamp 1757982896
transform 1 0 40100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9229
timestamp 1757982896
transform 1 0 41600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9230
timestamp 1757982896
transform 1 0 43100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9231
timestamp 1757982896
transform 1 0 44600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9232
timestamp 1757982896
transform 1 0 46100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9233
timestamp 1757982896
transform 1 0 47600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9234
timestamp 1757982896
transform 1 0 49100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9235
timestamp 1757982896
transform 1 0 50600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9236
timestamp 1757982896
transform 1 0 52100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9237
timestamp 1757982896
transform 1 0 53600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9238
timestamp 1757982896
transform 1 0 55100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9239
timestamp 1757982896
transform 1 0 56600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9240
timestamp 1757982896
transform 1 0 58100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9241
timestamp 1757982896
transform 1 0 59600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9242
timestamp 1757982896
transform 1 0 61100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9243
timestamp 1757982896
transform 1 0 62600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9244
timestamp 1757982896
transform 1 0 64100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9245
timestamp 1757982896
transform 1 0 65600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9246
timestamp 1757982896
transform 1 0 67100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9247
timestamp 1757982896
transform 1 0 68600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9248
timestamp 1757982896
transform 1 0 70100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9249
timestamp 1757982896
transform 1 0 71600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9250
timestamp 1757982896
transform 1 0 73100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9251
timestamp 1757982896
transform 1 0 74600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9252
timestamp 1757982896
transform 1 0 76100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9253
timestamp 1757982896
transform 1 0 77600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9254
timestamp 1757982896
transform 1 0 79100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9255
timestamp 1757982896
transform 1 0 80600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9256
timestamp 1757982896
transform 1 0 82100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9257
timestamp 1757982896
transform 1 0 83600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9258
timestamp 1757982896
transform 1 0 85100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9259
timestamp 1757982896
transform 1 0 86600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9260
timestamp 1757982896
transform 1 0 88100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9261
timestamp 1757982896
transform 1 0 89600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9262
timestamp 1757982896
transform 1 0 91100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9263
timestamp 1757982896
transform 1 0 92600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9264
timestamp 1757982896
transform 1 0 94100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9265
timestamp 1757982896
transform 1 0 95600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9266
timestamp 1757982896
transform 1 0 97100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9267
timestamp 1757982896
transform 1 0 98600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9268
timestamp 1757982896
transform 1 0 100100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9269
timestamp 1757982896
transform 1 0 101600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9270
timestamp 1757982896
transform 1 0 103100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9271
timestamp 1757982896
transform 1 0 104600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9272
timestamp 1757982896
transform 1 0 106100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9273
timestamp 1757982896
transform 1 0 107600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9274
timestamp 1757982896
transform 1 0 109100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9275
timestamp 1757982896
transform 1 0 110600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9276
timestamp 1757982896
transform 1 0 112100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9277
timestamp 1757982896
transform 1 0 113600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9278
timestamp 1757982896
transform 1 0 115100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9279
timestamp 1757982896
transform 1 0 116600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9280
timestamp 1757982896
transform 1 0 118100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9281
timestamp 1757982896
transform 1 0 119600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9282
timestamp 1757982896
transform 1 0 121100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9283
timestamp 1757982896
transform 1 0 122600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9284
timestamp 1757982896
transform 1 0 124100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9285
timestamp 1757982896
transform 1 0 125600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9286
timestamp 1757982896
transform 1 0 127100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9287
timestamp 1757982896
transform 1 0 128600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9288
timestamp 1757982896
transform 1 0 130100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9289
timestamp 1757982896
transform 1 0 131600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9290
timestamp 1757982896
transform 1 0 133100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9291
timestamp 1757982896
transform 1 0 134600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9292
timestamp 1757982896
transform 1 0 136100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9293
timestamp 1757982896
transform 1 0 137600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9294
timestamp 1757982896
transform 1 0 139100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9295
timestamp 1757982896
transform 1 0 140600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9296
timestamp 1757982896
transform 1 0 142100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9297
timestamp 1757982896
transform 1 0 143600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9298
timestamp 1757982896
transform 1 0 145100 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9299
timestamp 1757982896
transform 1 0 146600 0 1 -136650
box 1820 -1430 3480 230
use pixel  pixel_9300
timestamp 1757982896
transform 1 0 -1900 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9301
timestamp 1757982896
transform 1 0 -400 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9302
timestamp 1757982896
transform 1 0 1100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9303
timestamp 1757982896
transform 1 0 2600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9304
timestamp 1757982896
transform 1 0 4100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9305
timestamp 1757982896
transform 1 0 5600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9306
timestamp 1757982896
transform 1 0 7100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9307
timestamp 1757982896
transform 1 0 8600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9308
timestamp 1757982896
transform 1 0 10100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9309
timestamp 1757982896
transform 1 0 11600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9310
timestamp 1757982896
transform 1 0 13100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9311
timestamp 1757982896
transform 1 0 14600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9312
timestamp 1757982896
transform 1 0 16100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9313
timestamp 1757982896
transform 1 0 17600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9314
timestamp 1757982896
transform 1 0 19100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9315
timestamp 1757982896
transform 1 0 20600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9316
timestamp 1757982896
transform 1 0 22100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9317
timestamp 1757982896
transform 1 0 23600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9318
timestamp 1757982896
transform 1 0 25100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9319
timestamp 1757982896
transform 1 0 26600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9320
timestamp 1757982896
transform 1 0 28100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9321
timestamp 1757982896
transform 1 0 29600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9322
timestamp 1757982896
transform 1 0 31100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9323
timestamp 1757982896
transform 1 0 32600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9324
timestamp 1757982896
transform 1 0 34100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9325
timestamp 1757982896
transform 1 0 35600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9326
timestamp 1757982896
transform 1 0 37100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9327
timestamp 1757982896
transform 1 0 38600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9328
timestamp 1757982896
transform 1 0 40100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9329
timestamp 1757982896
transform 1 0 41600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9330
timestamp 1757982896
transform 1 0 43100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9331
timestamp 1757982896
transform 1 0 44600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9332
timestamp 1757982896
transform 1 0 46100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9333
timestamp 1757982896
transform 1 0 47600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9334
timestamp 1757982896
transform 1 0 49100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9335
timestamp 1757982896
transform 1 0 50600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9336
timestamp 1757982896
transform 1 0 52100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9337
timestamp 1757982896
transform 1 0 53600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9338
timestamp 1757982896
transform 1 0 55100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9339
timestamp 1757982896
transform 1 0 56600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9340
timestamp 1757982896
transform 1 0 58100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9341
timestamp 1757982896
transform 1 0 59600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9342
timestamp 1757982896
transform 1 0 61100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9343
timestamp 1757982896
transform 1 0 62600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9344
timestamp 1757982896
transform 1 0 64100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9345
timestamp 1757982896
transform 1 0 65600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9346
timestamp 1757982896
transform 1 0 67100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9347
timestamp 1757982896
transform 1 0 68600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9348
timestamp 1757982896
transform 1 0 70100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9349
timestamp 1757982896
transform 1 0 71600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9350
timestamp 1757982896
transform 1 0 73100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9351
timestamp 1757982896
transform 1 0 74600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9352
timestamp 1757982896
transform 1 0 76100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9353
timestamp 1757982896
transform 1 0 77600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9354
timestamp 1757982896
transform 1 0 79100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9355
timestamp 1757982896
transform 1 0 80600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9356
timestamp 1757982896
transform 1 0 82100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9357
timestamp 1757982896
transform 1 0 83600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9358
timestamp 1757982896
transform 1 0 85100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9359
timestamp 1757982896
transform 1 0 86600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9360
timestamp 1757982896
transform 1 0 88100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9361
timestamp 1757982896
transform 1 0 89600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9362
timestamp 1757982896
transform 1 0 91100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9363
timestamp 1757982896
transform 1 0 92600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9364
timestamp 1757982896
transform 1 0 94100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9365
timestamp 1757982896
transform 1 0 95600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9366
timestamp 1757982896
transform 1 0 97100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9367
timestamp 1757982896
transform 1 0 98600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9368
timestamp 1757982896
transform 1 0 100100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9369
timestamp 1757982896
transform 1 0 101600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9370
timestamp 1757982896
transform 1 0 103100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9371
timestamp 1757982896
transform 1 0 104600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9372
timestamp 1757982896
transform 1 0 106100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9373
timestamp 1757982896
transform 1 0 107600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9374
timestamp 1757982896
transform 1 0 109100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9375
timestamp 1757982896
transform 1 0 110600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9376
timestamp 1757982896
transform 1 0 112100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9377
timestamp 1757982896
transform 1 0 113600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9378
timestamp 1757982896
transform 1 0 115100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9379
timestamp 1757982896
transform 1 0 116600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9380
timestamp 1757982896
transform 1 0 118100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9381
timestamp 1757982896
transform 1 0 119600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9382
timestamp 1757982896
transform 1 0 121100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9383
timestamp 1757982896
transform 1 0 122600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9384
timestamp 1757982896
transform 1 0 124100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9385
timestamp 1757982896
transform 1 0 125600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9386
timestamp 1757982896
transform 1 0 127100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9387
timestamp 1757982896
transform 1 0 128600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9388
timestamp 1757982896
transform 1 0 130100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9389
timestamp 1757982896
transform 1 0 131600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9390
timestamp 1757982896
transform 1 0 133100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9391
timestamp 1757982896
transform 1 0 134600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9392
timestamp 1757982896
transform 1 0 136100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9393
timestamp 1757982896
transform 1 0 137600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9394
timestamp 1757982896
transform 1 0 139100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9395
timestamp 1757982896
transform 1 0 140600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9396
timestamp 1757982896
transform 1 0 142100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9397
timestamp 1757982896
transform 1 0 143600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9398
timestamp 1757982896
transform 1 0 145100 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9399
timestamp 1757982896
transform 1 0 146600 0 1 -138150
box 1820 -1430 3480 230
use pixel  pixel_9400
timestamp 1757982896
transform 1 0 -1900 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9401
timestamp 1757982896
transform 1 0 -400 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9402
timestamp 1757982896
transform 1 0 1100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9403
timestamp 1757982896
transform 1 0 2600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9404
timestamp 1757982896
transform 1 0 4100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9405
timestamp 1757982896
transform 1 0 5600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9406
timestamp 1757982896
transform 1 0 7100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9407
timestamp 1757982896
transform 1 0 8600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9408
timestamp 1757982896
transform 1 0 10100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9409
timestamp 1757982896
transform 1 0 11600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9410
timestamp 1757982896
transform 1 0 13100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9411
timestamp 1757982896
transform 1 0 14600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9412
timestamp 1757982896
transform 1 0 16100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9413
timestamp 1757982896
transform 1 0 17600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9414
timestamp 1757982896
transform 1 0 19100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9415
timestamp 1757982896
transform 1 0 20600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9416
timestamp 1757982896
transform 1 0 22100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9417
timestamp 1757982896
transform 1 0 23600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9418
timestamp 1757982896
transform 1 0 25100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9419
timestamp 1757982896
transform 1 0 26600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9420
timestamp 1757982896
transform 1 0 28100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9421
timestamp 1757982896
transform 1 0 29600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9422
timestamp 1757982896
transform 1 0 31100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9423
timestamp 1757982896
transform 1 0 32600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9424
timestamp 1757982896
transform 1 0 34100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9425
timestamp 1757982896
transform 1 0 35600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9426
timestamp 1757982896
transform 1 0 37100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9427
timestamp 1757982896
transform 1 0 38600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9428
timestamp 1757982896
transform 1 0 40100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9429
timestamp 1757982896
transform 1 0 41600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9430
timestamp 1757982896
transform 1 0 43100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9431
timestamp 1757982896
transform 1 0 44600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9432
timestamp 1757982896
transform 1 0 46100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9433
timestamp 1757982896
transform 1 0 47600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9434
timestamp 1757982896
transform 1 0 49100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9435
timestamp 1757982896
transform 1 0 50600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9436
timestamp 1757982896
transform 1 0 52100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9437
timestamp 1757982896
transform 1 0 53600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9438
timestamp 1757982896
transform 1 0 55100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9439
timestamp 1757982896
transform 1 0 56600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9440
timestamp 1757982896
transform 1 0 58100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9441
timestamp 1757982896
transform 1 0 59600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9442
timestamp 1757982896
transform 1 0 61100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9443
timestamp 1757982896
transform 1 0 62600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9444
timestamp 1757982896
transform 1 0 64100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9445
timestamp 1757982896
transform 1 0 65600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9446
timestamp 1757982896
transform 1 0 67100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9447
timestamp 1757982896
transform 1 0 68600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9448
timestamp 1757982896
transform 1 0 70100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9449
timestamp 1757982896
transform 1 0 71600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9450
timestamp 1757982896
transform 1 0 73100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9451
timestamp 1757982896
transform 1 0 74600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9452
timestamp 1757982896
transform 1 0 76100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9453
timestamp 1757982896
transform 1 0 77600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9454
timestamp 1757982896
transform 1 0 79100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9455
timestamp 1757982896
transform 1 0 80600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9456
timestamp 1757982896
transform 1 0 82100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9457
timestamp 1757982896
transform 1 0 83600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9458
timestamp 1757982896
transform 1 0 85100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9459
timestamp 1757982896
transform 1 0 86600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9460
timestamp 1757982896
transform 1 0 88100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9461
timestamp 1757982896
transform 1 0 89600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9462
timestamp 1757982896
transform 1 0 91100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9463
timestamp 1757982896
transform 1 0 92600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9464
timestamp 1757982896
transform 1 0 94100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9465
timestamp 1757982896
transform 1 0 95600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9466
timestamp 1757982896
transform 1 0 97100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9467
timestamp 1757982896
transform 1 0 98600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9468
timestamp 1757982896
transform 1 0 100100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9469
timestamp 1757982896
transform 1 0 101600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9470
timestamp 1757982896
transform 1 0 103100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9471
timestamp 1757982896
transform 1 0 104600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9472
timestamp 1757982896
transform 1 0 106100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9473
timestamp 1757982896
transform 1 0 107600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9474
timestamp 1757982896
transform 1 0 109100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9475
timestamp 1757982896
transform 1 0 110600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9476
timestamp 1757982896
transform 1 0 112100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9477
timestamp 1757982896
transform 1 0 113600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9478
timestamp 1757982896
transform 1 0 115100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9479
timestamp 1757982896
transform 1 0 116600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9480
timestamp 1757982896
transform 1 0 118100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9481
timestamp 1757982896
transform 1 0 119600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9482
timestamp 1757982896
transform 1 0 121100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9483
timestamp 1757982896
transform 1 0 122600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9484
timestamp 1757982896
transform 1 0 124100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9485
timestamp 1757982896
transform 1 0 125600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9486
timestamp 1757982896
transform 1 0 127100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9487
timestamp 1757982896
transform 1 0 128600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9488
timestamp 1757982896
transform 1 0 130100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9489
timestamp 1757982896
transform 1 0 131600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9490
timestamp 1757982896
transform 1 0 133100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9491
timestamp 1757982896
transform 1 0 134600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9492
timestamp 1757982896
transform 1 0 136100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9493
timestamp 1757982896
transform 1 0 137600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9494
timestamp 1757982896
transform 1 0 139100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9495
timestamp 1757982896
transform 1 0 140600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9496
timestamp 1757982896
transform 1 0 142100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9497
timestamp 1757982896
transform 1 0 143600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9498
timestamp 1757982896
transform 1 0 145100 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9499
timestamp 1757982896
transform 1 0 146600 0 1 -139650
box 1820 -1430 3480 230
use pixel  pixel_9500
timestamp 1757982896
transform 1 0 -1900 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9501
timestamp 1757982896
transform 1 0 -400 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9502
timestamp 1757982896
transform 1 0 1100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9503
timestamp 1757982896
transform 1 0 2600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9504
timestamp 1757982896
transform 1 0 4100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9505
timestamp 1757982896
transform 1 0 5600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9506
timestamp 1757982896
transform 1 0 7100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9507
timestamp 1757982896
transform 1 0 8600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9508
timestamp 1757982896
transform 1 0 10100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9509
timestamp 1757982896
transform 1 0 11600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9510
timestamp 1757982896
transform 1 0 13100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9511
timestamp 1757982896
transform 1 0 14600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9512
timestamp 1757982896
transform 1 0 16100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9513
timestamp 1757982896
transform 1 0 17600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9514
timestamp 1757982896
transform 1 0 19100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9515
timestamp 1757982896
transform 1 0 20600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9516
timestamp 1757982896
transform 1 0 22100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9517
timestamp 1757982896
transform 1 0 23600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9518
timestamp 1757982896
transform 1 0 25100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9519
timestamp 1757982896
transform 1 0 26600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9520
timestamp 1757982896
transform 1 0 28100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9521
timestamp 1757982896
transform 1 0 29600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9522
timestamp 1757982896
transform 1 0 31100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9523
timestamp 1757982896
transform 1 0 32600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9524
timestamp 1757982896
transform 1 0 34100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9525
timestamp 1757982896
transform 1 0 35600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9526
timestamp 1757982896
transform 1 0 37100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9527
timestamp 1757982896
transform 1 0 38600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9528
timestamp 1757982896
transform 1 0 40100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9529
timestamp 1757982896
transform 1 0 41600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9530
timestamp 1757982896
transform 1 0 43100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9531
timestamp 1757982896
transform 1 0 44600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9532
timestamp 1757982896
transform 1 0 46100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9533
timestamp 1757982896
transform 1 0 47600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9534
timestamp 1757982896
transform 1 0 49100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9535
timestamp 1757982896
transform 1 0 50600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9536
timestamp 1757982896
transform 1 0 52100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9537
timestamp 1757982896
transform 1 0 53600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9538
timestamp 1757982896
transform 1 0 55100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9539
timestamp 1757982896
transform 1 0 56600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9540
timestamp 1757982896
transform 1 0 58100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9541
timestamp 1757982896
transform 1 0 59600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9542
timestamp 1757982896
transform 1 0 61100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9543
timestamp 1757982896
transform 1 0 62600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9544
timestamp 1757982896
transform 1 0 64100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9545
timestamp 1757982896
transform 1 0 65600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9546
timestamp 1757982896
transform 1 0 67100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9547
timestamp 1757982896
transform 1 0 68600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9548
timestamp 1757982896
transform 1 0 70100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9549
timestamp 1757982896
transform 1 0 71600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9550
timestamp 1757982896
transform 1 0 73100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9551
timestamp 1757982896
transform 1 0 74600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9552
timestamp 1757982896
transform 1 0 76100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9553
timestamp 1757982896
transform 1 0 77600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9554
timestamp 1757982896
transform 1 0 79100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9555
timestamp 1757982896
transform 1 0 80600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9556
timestamp 1757982896
transform 1 0 82100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9557
timestamp 1757982896
transform 1 0 83600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9558
timestamp 1757982896
transform 1 0 85100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9559
timestamp 1757982896
transform 1 0 86600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9560
timestamp 1757982896
transform 1 0 88100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9561
timestamp 1757982896
transform 1 0 89600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9562
timestamp 1757982896
transform 1 0 91100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9563
timestamp 1757982896
transform 1 0 92600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9564
timestamp 1757982896
transform 1 0 94100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9565
timestamp 1757982896
transform 1 0 95600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9566
timestamp 1757982896
transform 1 0 97100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9567
timestamp 1757982896
transform 1 0 98600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9568
timestamp 1757982896
transform 1 0 100100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9569
timestamp 1757982896
transform 1 0 101600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9570
timestamp 1757982896
transform 1 0 103100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9571
timestamp 1757982896
transform 1 0 104600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9572
timestamp 1757982896
transform 1 0 106100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9573
timestamp 1757982896
transform 1 0 107600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9574
timestamp 1757982896
transform 1 0 109100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9575
timestamp 1757982896
transform 1 0 110600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9576
timestamp 1757982896
transform 1 0 112100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9577
timestamp 1757982896
transform 1 0 113600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9578
timestamp 1757982896
transform 1 0 115100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9579
timestamp 1757982896
transform 1 0 116600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9580
timestamp 1757982896
transform 1 0 118100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9581
timestamp 1757982896
transform 1 0 119600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9582
timestamp 1757982896
transform 1 0 121100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9583
timestamp 1757982896
transform 1 0 122600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9584
timestamp 1757982896
transform 1 0 124100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9585
timestamp 1757982896
transform 1 0 125600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9586
timestamp 1757982896
transform 1 0 127100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9587
timestamp 1757982896
transform 1 0 128600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9588
timestamp 1757982896
transform 1 0 130100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9589
timestamp 1757982896
transform 1 0 131600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9590
timestamp 1757982896
transform 1 0 133100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9591
timestamp 1757982896
transform 1 0 134600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9592
timestamp 1757982896
transform 1 0 136100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9593
timestamp 1757982896
transform 1 0 137600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9594
timestamp 1757982896
transform 1 0 139100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9595
timestamp 1757982896
transform 1 0 140600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9596
timestamp 1757982896
transform 1 0 142100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9597
timestamp 1757982896
transform 1 0 143600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9598
timestamp 1757982896
transform 1 0 145100 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9599
timestamp 1757982896
transform 1 0 146600 0 1 -141150
box 1820 -1430 3480 230
use pixel  pixel_9600
timestamp 1757982896
transform 1 0 -1900 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9601
timestamp 1757982896
transform 1 0 -400 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9602
timestamp 1757982896
transform 1 0 1100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9603
timestamp 1757982896
transform 1 0 2600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9604
timestamp 1757982896
transform 1 0 4100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9605
timestamp 1757982896
transform 1 0 5600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9606
timestamp 1757982896
transform 1 0 7100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9607
timestamp 1757982896
transform 1 0 8600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9608
timestamp 1757982896
transform 1 0 10100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9609
timestamp 1757982896
transform 1 0 11600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9610
timestamp 1757982896
transform 1 0 13100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9611
timestamp 1757982896
transform 1 0 14600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9612
timestamp 1757982896
transform 1 0 16100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9613
timestamp 1757982896
transform 1 0 17600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9614
timestamp 1757982896
transform 1 0 19100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9615
timestamp 1757982896
transform 1 0 20600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9616
timestamp 1757982896
transform 1 0 22100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9617
timestamp 1757982896
transform 1 0 23600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9618
timestamp 1757982896
transform 1 0 25100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9619
timestamp 1757982896
transform 1 0 26600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9620
timestamp 1757982896
transform 1 0 28100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9621
timestamp 1757982896
transform 1 0 29600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9622
timestamp 1757982896
transform 1 0 31100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9623
timestamp 1757982896
transform 1 0 32600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9624
timestamp 1757982896
transform 1 0 34100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9625
timestamp 1757982896
transform 1 0 35600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9626
timestamp 1757982896
transform 1 0 37100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9627
timestamp 1757982896
transform 1 0 38600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9628
timestamp 1757982896
transform 1 0 40100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9629
timestamp 1757982896
transform 1 0 41600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9630
timestamp 1757982896
transform 1 0 43100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9631
timestamp 1757982896
transform 1 0 44600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9632
timestamp 1757982896
transform 1 0 46100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9633
timestamp 1757982896
transform 1 0 47600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9634
timestamp 1757982896
transform 1 0 49100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9635
timestamp 1757982896
transform 1 0 50600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9636
timestamp 1757982896
transform 1 0 52100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9637
timestamp 1757982896
transform 1 0 53600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9638
timestamp 1757982896
transform 1 0 55100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9639
timestamp 1757982896
transform 1 0 56600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9640
timestamp 1757982896
transform 1 0 58100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9641
timestamp 1757982896
transform 1 0 59600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9642
timestamp 1757982896
transform 1 0 61100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9643
timestamp 1757982896
transform 1 0 62600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9644
timestamp 1757982896
transform 1 0 64100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9645
timestamp 1757982896
transform 1 0 65600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9646
timestamp 1757982896
transform 1 0 67100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9647
timestamp 1757982896
transform 1 0 68600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9648
timestamp 1757982896
transform 1 0 70100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9649
timestamp 1757982896
transform 1 0 71600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9650
timestamp 1757982896
transform 1 0 73100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9651
timestamp 1757982896
transform 1 0 74600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9652
timestamp 1757982896
transform 1 0 76100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9653
timestamp 1757982896
transform 1 0 77600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9654
timestamp 1757982896
transform 1 0 79100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9655
timestamp 1757982896
transform 1 0 80600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9656
timestamp 1757982896
transform 1 0 82100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9657
timestamp 1757982896
transform 1 0 83600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9658
timestamp 1757982896
transform 1 0 85100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9659
timestamp 1757982896
transform 1 0 86600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9660
timestamp 1757982896
transform 1 0 88100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9661
timestamp 1757982896
transform 1 0 89600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9662
timestamp 1757982896
transform 1 0 91100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9663
timestamp 1757982896
transform 1 0 92600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9664
timestamp 1757982896
transform 1 0 94100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9665
timestamp 1757982896
transform 1 0 95600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9666
timestamp 1757982896
transform 1 0 97100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9667
timestamp 1757982896
transform 1 0 98600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9668
timestamp 1757982896
transform 1 0 100100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9669
timestamp 1757982896
transform 1 0 101600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9670
timestamp 1757982896
transform 1 0 103100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9671
timestamp 1757982896
transform 1 0 104600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9672
timestamp 1757982896
transform 1 0 106100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9673
timestamp 1757982896
transform 1 0 107600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9674
timestamp 1757982896
transform 1 0 109100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9675
timestamp 1757982896
transform 1 0 110600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9676
timestamp 1757982896
transform 1 0 112100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9677
timestamp 1757982896
transform 1 0 113600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9678
timestamp 1757982896
transform 1 0 115100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9679
timestamp 1757982896
transform 1 0 116600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9680
timestamp 1757982896
transform 1 0 118100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9681
timestamp 1757982896
transform 1 0 119600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9682
timestamp 1757982896
transform 1 0 121100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9683
timestamp 1757982896
transform 1 0 122600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9684
timestamp 1757982896
transform 1 0 124100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9685
timestamp 1757982896
transform 1 0 125600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9686
timestamp 1757982896
transform 1 0 127100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9687
timestamp 1757982896
transform 1 0 128600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9688
timestamp 1757982896
transform 1 0 130100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9689
timestamp 1757982896
transform 1 0 131600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9690
timestamp 1757982896
transform 1 0 133100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9691
timestamp 1757982896
transform 1 0 134600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9692
timestamp 1757982896
transform 1 0 136100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9693
timestamp 1757982896
transform 1 0 137600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9694
timestamp 1757982896
transform 1 0 139100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9695
timestamp 1757982896
transform 1 0 140600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9696
timestamp 1757982896
transform 1 0 142100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9697
timestamp 1757982896
transform 1 0 143600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9698
timestamp 1757982896
transform 1 0 145100 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9699
timestamp 1757982896
transform 1 0 146600 0 1 -142650
box 1820 -1430 3480 230
use pixel  pixel_9700
timestamp 1757982896
transform 1 0 -1900 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9701
timestamp 1757982896
transform 1 0 -400 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9702
timestamp 1757982896
transform 1 0 1100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9703
timestamp 1757982896
transform 1 0 2600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9704
timestamp 1757982896
transform 1 0 4100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9705
timestamp 1757982896
transform 1 0 5600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9706
timestamp 1757982896
transform 1 0 7100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9707
timestamp 1757982896
transform 1 0 8600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9708
timestamp 1757982896
transform 1 0 10100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9709
timestamp 1757982896
transform 1 0 11600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9710
timestamp 1757982896
transform 1 0 13100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9711
timestamp 1757982896
transform 1 0 14600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9712
timestamp 1757982896
transform 1 0 16100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9713
timestamp 1757982896
transform 1 0 17600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9714
timestamp 1757982896
transform 1 0 19100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9715
timestamp 1757982896
transform 1 0 20600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9716
timestamp 1757982896
transform 1 0 22100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9717
timestamp 1757982896
transform 1 0 23600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9718
timestamp 1757982896
transform 1 0 25100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9719
timestamp 1757982896
transform 1 0 26600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9720
timestamp 1757982896
transform 1 0 28100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9721
timestamp 1757982896
transform 1 0 29600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9722
timestamp 1757982896
transform 1 0 31100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9723
timestamp 1757982896
transform 1 0 32600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9724
timestamp 1757982896
transform 1 0 34100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9725
timestamp 1757982896
transform 1 0 35600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9726
timestamp 1757982896
transform 1 0 37100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9727
timestamp 1757982896
transform 1 0 38600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9728
timestamp 1757982896
transform 1 0 40100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9729
timestamp 1757982896
transform 1 0 41600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9730
timestamp 1757982896
transform 1 0 43100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9731
timestamp 1757982896
transform 1 0 44600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9732
timestamp 1757982896
transform 1 0 46100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9733
timestamp 1757982896
transform 1 0 47600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9734
timestamp 1757982896
transform 1 0 49100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9735
timestamp 1757982896
transform 1 0 50600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9736
timestamp 1757982896
transform 1 0 52100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9737
timestamp 1757982896
transform 1 0 53600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9738
timestamp 1757982896
transform 1 0 55100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9739
timestamp 1757982896
transform 1 0 56600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9740
timestamp 1757982896
transform 1 0 58100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9741
timestamp 1757982896
transform 1 0 59600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9742
timestamp 1757982896
transform 1 0 61100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9743
timestamp 1757982896
transform 1 0 62600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9744
timestamp 1757982896
transform 1 0 64100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9745
timestamp 1757982896
transform 1 0 65600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9746
timestamp 1757982896
transform 1 0 67100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9747
timestamp 1757982896
transform 1 0 68600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9748
timestamp 1757982896
transform 1 0 70100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9749
timestamp 1757982896
transform 1 0 71600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9750
timestamp 1757982896
transform 1 0 73100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9751
timestamp 1757982896
transform 1 0 74600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9752
timestamp 1757982896
transform 1 0 76100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9753
timestamp 1757982896
transform 1 0 77600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9754
timestamp 1757982896
transform 1 0 79100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9755
timestamp 1757982896
transform 1 0 80600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9756
timestamp 1757982896
transform 1 0 82100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9757
timestamp 1757982896
transform 1 0 83600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9758
timestamp 1757982896
transform 1 0 85100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9759
timestamp 1757982896
transform 1 0 86600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9760
timestamp 1757982896
transform 1 0 88100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9761
timestamp 1757982896
transform 1 0 89600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9762
timestamp 1757982896
transform 1 0 91100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9763
timestamp 1757982896
transform 1 0 92600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9764
timestamp 1757982896
transform 1 0 94100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9765
timestamp 1757982896
transform 1 0 95600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9766
timestamp 1757982896
transform 1 0 97100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9767
timestamp 1757982896
transform 1 0 98600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9768
timestamp 1757982896
transform 1 0 100100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9769
timestamp 1757982896
transform 1 0 101600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9770
timestamp 1757982896
transform 1 0 103100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9771
timestamp 1757982896
transform 1 0 104600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9772
timestamp 1757982896
transform 1 0 106100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9773
timestamp 1757982896
transform 1 0 107600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9774
timestamp 1757982896
transform 1 0 109100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9775
timestamp 1757982896
transform 1 0 110600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9776
timestamp 1757982896
transform 1 0 112100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9777
timestamp 1757982896
transform 1 0 113600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9778
timestamp 1757982896
transform 1 0 115100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9779
timestamp 1757982896
transform 1 0 116600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9780
timestamp 1757982896
transform 1 0 118100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9781
timestamp 1757982896
transform 1 0 119600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9782
timestamp 1757982896
transform 1 0 121100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9783
timestamp 1757982896
transform 1 0 122600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9784
timestamp 1757982896
transform 1 0 124100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9785
timestamp 1757982896
transform 1 0 125600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9786
timestamp 1757982896
transform 1 0 127100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9787
timestamp 1757982896
transform 1 0 128600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9788
timestamp 1757982896
transform 1 0 130100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9789
timestamp 1757982896
transform 1 0 131600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9790
timestamp 1757982896
transform 1 0 133100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9791
timestamp 1757982896
transform 1 0 134600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9792
timestamp 1757982896
transform 1 0 136100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9793
timestamp 1757982896
transform 1 0 137600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9794
timestamp 1757982896
transform 1 0 139100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9795
timestamp 1757982896
transform 1 0 140600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9796
timestamp 1757982896
transform 1 0 142100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9797
timestamp 1757982896
transform 1 0 143600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9798
timestamp 1757982896
transform 1 0 145100 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9799
timestamp 1757982896
transform 1 0 146600 0 1 -144150
box 1820 -1430 3480 230
use pixel  pixel_9800
timestamp 1757982896
transform 1 0 -1900 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9801
timestamp 1757982896
transform 1 0 -400 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9802
timestamp 1757982896
transform 1 0 1100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9803
timestamp 1757982896
transform 1 0 2600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9804
timestamp 1757982896
transform 1 0 4100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9805
timestamp 1757982896
transform 1 0 5600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9806
timestamp 1757982896
transform 1 0 7100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9807
timestamp 1757982896
transform 1 0 8600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9808
timestamp 1757982896
transform 1 0 10100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9809
timestamp 1757982896
transform 1 0 11600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9810
timestamp 1757982896
transform 1 0 13100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9811
timestamp 1757982896
transform 1 0 14600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9812
timestamp 1757982896
transform 1 0 16100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9813
timestamp 1757982896
transform 1 0 17600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9814
timestamp 1757982896
transform 1 0 19100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9815
timestamp 1757982896
transform 1 0 20600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9816
timestamp 1757982896
transform 1 0 22100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9817
timestamp 1757982896
transform 1 0 23600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9818
timestamp 1757982896
transform 1 0 25100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9819
timestamp 1757982896
transform 1 0 26600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9820
timestamp 1757982896
transform 1 0 28100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9821
timestamp 1757982896
transform 1 0 29600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9822
timestamp 1757982896
transform 1 0 31100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9823
timestamp 1757982896
transform 1 0 32600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9824
timestamp 1757982896
transform 1 0 34100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9825
timestamp 1757982896
transform 1 0 35600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9826
timestamp 1757982896
transform 1 0 37100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9827
timestamp 1757982896
transform 1 0 38600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9828
timestamp 1757982896
transform 1 0 40100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9829
timestamp 1757982896
transform 1 0 41600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9830
timestamp 1757982896
transform 1 0 43100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9831
timestamp 1757982896
transform 1 0 44600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9832
timestamp 1757982896
transform 1 0 46100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9833
timestamp 1757982896
transform 1 0 47600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9834
timestamp 1757982896
transform 1 0 49100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9835
timestamp 1757982896
transform 1 0 50600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9836
timestamp 1757982896
transform 1 0 52100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9837
timestamp 1757982896
transform 1 0 53600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9838
timestamp 1757982896
transform 1 0 55100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9839
timestamp 1757982896
transform 1 0 56600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9840
timestamp 1757982896
transform 1 0 58100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9841
timestamp 1757982896
transform 1 0 59600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9842
timestamp 1757982896
transform 1 0 61100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9843
timestamp 1757982896
transform 1 0 62600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9844
timestamp 1757982896
transform 1 0 64100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9845
timestamp 1757982896
transform 1 0 65600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9846
timestamp 1757982896
transform 1 0 67100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9847
timestamp 1757982896
transform 1 0 68600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9848
timestamp 1757982896
transform 1 0 70100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9849
timestamp 1757982896
transform 1 0 71600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9850
timestamp 1757982896
transform 1 0 73100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9851
timestamp 1757982896
transform 1 0 74600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9852
timestamp 1757982896
transform 1 0 76100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9853
timestamp 1757982896
transform 1 0 77600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9854
timestamp 1757982896
transform 1 0 79100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9855
timestamp 1757982896
transform 1 0 80600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9856
timestamp 1757982896
transform 1 0 82100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9857
timestamp 1757982896
transform 1 0 83600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9858
timestamp 1757982896
transform 1 0 85100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9859
timestamp 1757982896
transform 1 0 86600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9860
timestamp 1757982896
transform 1 0 88100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9861
timestamp 1757982896
transform 1 0 89600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9862
timestamp 1757982896
transform 1 0 91100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9863
timestamp 1757982896
transform 1 0 92600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9864
timestamp 1757982896
transform 1 0 94100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9865
timestamp 1757982896
transform 1 0 95600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9866
timestamp 1757982896
transform 1 0 97100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9867
timestamp 1757982896
transform 1 0 98600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9868
timestamp 1757982896
transform 1 0 100100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9869
timestamp 1757982896
transform 1 0 101600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9870
timestamp 1757982896
transform 1 0 103100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9871
timestamp 1757982896
transform 1 0 104600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9872
timestamp 1757982896
transform 1 0 106100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9873
timestamp 1757982896
transform 1 0 107600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9874
timestamp 1757982896
transform 1 0 109100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9875
timestamp 1757982896
transform 1 0 110600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9876
timestamp 1757982896
transform 1 0 112100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9877
timestamp 1757982896
transform 1 0 113600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9878
timestamp 1757982896
transform 1 0 115100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9879
timestamp 1757982896
transform 1 0 116600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9880
timestamp 1757982896
transform 1 0 118100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9881
timestamp 1757982896
transform 1 0 119600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9882
timestamp 1757982896
transform 1 0 121100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9883
timestamp 1757982896
transform 1 0 122600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9884
timestamp 1757982896
transform 1 0 124100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9885
timestamp 1757982896
transform 1 0 125600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9886
timestamp 1757982896
transform 1 0 127100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9887
timestamp 1757982896
transform 1 0 128600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9888
timestamp 1757982896
transform 1 0 130100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9889
timestamp 1757982896
transform 1 0 131600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9890
timestamp 1757982896
transform 1 0 133100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9891
timestamp 1757982896
transform 1 0 134600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9892
timestamp 1757982896
transform 1 0 136100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9893
timestamp 1757982896
transform 1 0 137600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9894
timestamp 1757982896
transform 1 0 139100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9895
timestamp 1757982896
transform 1 0 140600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9896
timestamp 1757982896
transform 1 0 142100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9897
timestamp 1757982896
transform 1 0 143600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9898
timestamp 1757982896
transform 1 0 145100 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9899
timestamp 1757982896
transform 1 0 146600 0 1 -145650
box 1820 -1430 3480 230
use pixel  pixel_9900
timestamp 1757982896
transform 1 0 -1900 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9901
timestamp 1757982896
transform 1 0 -400 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9902
timestamp 1757982896
transform 1 0 1100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9903
timestamp 1757982896
transform 1 0 2600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9904
timestamp 1757982896
transform 1 0 4100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9905
timestamp 1757982896
transform 1 0 5600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9906
timestamp 1757982896
transform 1 0 7100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9907
timestamp 1757982896
transform 1 0 8600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9908
timestamp 1757982896
transform 1 0 10100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9909
timestamp 1757982896
transform 1 0 11600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9910
timestamp 1757982896
transform 1 0 13100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9911
timestamp 1757982896
transform 1 0 14600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9912
timestamp 1757982896
transform 1 0 16100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9913
timestamp 1757982896
transform 1 0 17600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9914
timestamp 1757982896
transform 1 0 19100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9915
timestamp 1757982896
transform 1 0 20600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9916
timestamp 1757982896
transform 1 0 22100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9917
timestamp 1757982896
transform 1 0 23600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9918
timestamp 1757982896
transform 1 0 25100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9919
timestamp 1757982896
transform 1 0 26600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9920
timestamp 1757982896
transform 1 0 28100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9921
timestamp 1757982896
transform 1 0 29600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9922
timestamp 1757982896
transform 1 0 31100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9923
timestamp 1757982896
transform 1 0 32600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9924
timestamp 1757982896
transform 1 0 34100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9925
timestamp 1757982896
transform 1 0 35600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9926
timestamp 1757982896
transform 1 0 37100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9927
timestamp 1757982896
transform 1 0 38600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9928
timestamp 1757982896
transform 1 0 40100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9929
timestamp 1757982896
transform 1 0 41600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9930
timestamp 1757982896
transform 1 0 43100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9931
timestamp 1757982896
transform 1 0 44600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9932
timestamp 1757982896
transform 1 0 46100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9933
timestamp 1757982896
transform 1 0 47600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9934
timestamp 1757982896
transform 1 0 49100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9935
timestamp 1757982896
transform 1 0 50600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9936
timestamp 1757982896
transform 1 0 52100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9937
timestamp 1757982896
transform 1 0 53600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9938
timestamp 1757982896
transform 1 0 55100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9939
timestamp 1757982896
transform 1 0 56600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9940
timestamp 1757982896
transform 1 0 58100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9941
timestamp 1757982896
transform 1 0 59600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9942
timestamp 1757982896
transform 1 0 61100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9943
timestamp 1757982896
transform 1 0 62600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9944
timestamp 1757982896
transform 1 0 64100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9945
timestamp 1757982896
transform 1 0 65600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9946
timestamp 1757982896
transform 1 0 67100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9947
timestamp 1757982896
transform 1 0 68600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9948
timestamp 1757982896
transform 1 0 70100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9949
timestamp 1757982896
transform 1 0 71600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9950
timestamp 1757982896
transform 1 0 73100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9951
timestamp 1757982896
transform 1 0 74600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9952
timestamp 1757982896
transform 1 0 76100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9953
timestamp 1757982896
transform 1 0 77600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9954
timestamp 1757982896
transform 1 0 79100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9955
timestamp 1757982896
transform 1 0 80600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9956
timestamp 1757982896
transform 1 0 82100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9957
timestamp 1757982896
transform 1 0 83600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9958
timestamp 1757982896
transform 1 0 85100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9959
timestamp 1757982896
transform 1 0 86600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9960
timestamp 1757982896
transform 1 0 88100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9961
timestamp 1757982896
transform 1 0 89600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9962
timestamp 1757982896
transform 1 0 91100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9963
timestamp 1757982896
transform 1 0 92600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9964
timestamp 1757982896
transform 1 0 94100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9965
timestamp 1757982896
transform 1 0 95600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9966
timestamp 1757982896
transform 1 0 97100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9967
timestamp 1757982896
transform 1 0 98600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9968
timestamp 1757982896
transform 1 0 100100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9969
timestamp 1757982896
transform 1 0 101600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9970
timestamp 1757982896
transform 1 0 103100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9971
timestamp 1757982896
transform 1 0 104600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9972
timestamp 1757982896
transform 1 0 106100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9973
timestamp 1757982896
transform 1 0 107600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9974
timestamp 1757982896
transform 1 0 109100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9975
timestamp 1757982896
transform 1 0 110600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9976
timestamp 1757982896
transform 1 0 112100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9977
timestamp 1757982896
transform 1 0 113600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9978
timestamp 1757982896
transform 1 0 115100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9979
timestamp 1757982896
transform 1 0 116600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9980
timestamp 1757982896
transform 1 0 118100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9981
timestamp 1757982896
transform 1 0 119600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9982
timestamp 1757982896
transform 1 0 121100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9983
timestamp 1757982896
transform 1 0 122600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9984
timestamp 1757982896
transform 1 0 124100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9985
timestamp 1757982896
transform 1 0 125600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9986
timestamp 1757982896
transform 1 0 127100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9987
timestamp 1757982896
transform 1 0 128600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9988
timestamp 1757982896
transform 1 0 130100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9989
timestamp 1757982896
transform 1 0 131600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9990
timestamp 1757982896
transform 1 0 133100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9991
timestamp 1757982896
transform 1 0 134600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9992
timestamp 1757982896
transform 1 0 136100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9993
timestamp 1757982896
transform 1 0 137600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9994
timestamp 1757982896
transform 1 0 139100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9995
timestamp 1757982896
transform 1 0 140600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9996
timestamp 1757982896
transform 1 0 142100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9997
timestamp 1757982896
transform 1 0 143600 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9998
timestamp 1757982896
transform 1 0 145100 0 1 -147150
box 1820 -1430 3480 230
use pixel  pixel_9999
timestamp 1757982896
transform 1 0 146600 0 1 -147150
box 1820 -1430 3480 230
<< labels >>
rlabel metal4 -1500 1775 -1500 1830 1 VBIAS
port 2 n
rlabel metal2 -1500 1675 -1500 1725 3 VREF
port 3 e
rlabel metal2 0 2020 0 2020 1 NB2
port 4 n
rlabel metal1 -1000 0 -1000 0 1 VDD
port 5 n
rlabel metal2 -370 1780 -370 1780 1 NB1
port 7 n
rlabel metal2 -1500 740 -1500 785 3 ROW_SEL[0]
port 8 e
rlabel metal5 -1000 1420 -1000 1420 1 GRING
port 9 n
rlabel metal1 150200 15 150200 15 1 GND
port 109 n
rlabel metal2 -1500 -760 -1500 -715 3 ROW_SEL[1]
port 111 e
rlabel metal2 -1500 -2260 -1500 -2215 3 ROW_SEL[2]
port 212 e
rlabel metal2 -1500 -3760 -1500 -3715 3 ROW_SEL[3]
port 313 e
rlabel metal2 -1500 -5260 -1500 -5215 3 ROW_SEL[4]
port 414 e
rlabel metal2 -1500 -6760 -1500 -6715 3 ROW_SEL[5]
port 515 e
rlabel metal2 -1500 -8260 -1500 -8215 3 ROW_SEL[6]
port 616 e
rlabel metal2 -1500 -9760 -1500 -9715 3 ROW_SEL[7]
port 717 e
rlabel metal2 -1500 -11260 -1500 -11215 3 ROW_SEL[8]
port 818 e
rlabel metal2 -1500 -12760 -1500 -12715 3 ROW_SEL[9]
port 919 e
rlabel metal2 -1500 -14260 -1500 -14215 3 ROW_SEL[10]
port 1020 e
rlabel metal2 -1500 -15760 -1500 -15715 3 ROW_SEL[11]
port 1121 e
rlabel metal2 -1500 -17260 -1500 -17215 3 ROW_SEL[12]
port 1222 e
rlabel metal2 -1500 -18760 -1500 -18715 3 ROW_SEL[13]
port 1323 e
rlabel metal2 -1500 -20260 -1500 -20215 3 ROW_SEL[14]
port 1424 e
rlabel metal2 -1500 -21760 -1500 -21715 3 ROW_SEL[15]
port 1525 e
rlabel metal2 -1500 -23260 -1500 -23215 3 ROW_SEL[16]
port 1626 e
rlabel metal2 -1500 -24760 -1500 -24715 3 ROW_SEL[17]
port 1727 e
rlabel metal2 -1500 -26260 -1500 -26215 3 ROW_SEL[18]
port 1828 e
rlabel metal2 -1500 -27760 -1500 -27715 3 ROW_SEL[19]
port 1929 e
rlabel metal2 -1500 -29260 -1500 -29215 3 ROW_SEL[20]
port 2030 e
rlabel metal2 -1500 -30760 -1500 -30715 3 ROW_SEL[21]
port 2131 e
rlabel metal2 -1500 -32260 -1500 -32215 3 ROW_SEL[22]
port 2232 e
rlabel metal2 -1500 -33760 -1500 -33715 3 ROW_SEL[23]
port 2333 e
rlabel metal2 -1500 -35260 -1500 -35215 3 ROW_SEL[24]
port 2434 e
rlabel metal2 -1500 -36760 -1500 -36715 3 ROW_SEL[25]
port 2535 e
rlabel metal2 -1500 -38260 -1500 -38215 3 ROW_SEL[26]
port 2636 e
rlabel metal2 -1500 -39760 -1500 -39715 3 ROW_SEL[27]
port 2737 e
rlabel metal2 -1500 -41260 -1500 -41215 3 ROW_SEL[28]
port 2838 e
rlabel metal2 -1500 -42760 -1500 -42715 3 ROW_SEL[29]
port 2939 e
rlabel metal2 -1500 -44260 -1500 -44215 3 ROW_SEL[30]
port 3040 e
rlabel metal2 -1500 -45760 -1500 -45715 3 ROW_SEL[31]
port 3141 e
rlabel metal2 -1500 -47260 -1500 -47215 3 ROW_SEL[32]
port 3242 e
rlabel metal2 -1500 -48760 -1500 -48715 3 ROW_SEL[33]
port 3343 e
rlabel metal2 -1500 -50260 -1500 -50215 3 ROW_SEL[34]
port 3444 e
rlabel metal2 -1500 -51760 -1500 -51715 3 ROW_SEL[35]
port 3545 e
rlabel metal2 -1500 -53260 -1500 -53215 3 ROW_SEL[36]
port 3646 e
rlabel metal2 -1500 -54760 -1500 -54715 3 ROW_SEL[37]
port 3747 e
rlabel metal2 -1500 -56260 -1500 -56215 3 ROW_SEL[38]
port 3848 e
rlabel metal2 -1500 -57760 -1500 -57715 3 ROW_SEL[39]
port 3949 e
rlabel metal2 -1500 -59260 -1500 -59215 3 ROW_SEL[40]
port 4050 e
rlabel metal2 -1500 -60760 -1500 -60715 3 ROW_SEL[41]
port 4151 e
rlabel metal2 -1500 -62260 -1500 -62215 3 ROW_SEL[42]
port 4252 e
rlabel metal2 -1500 -63760 -1500 -63715 3 ROW_SEL[43]
port 4353 e
rlabel metal2 -1500 -65260 -1500 -65215 3 ROW_SEL[44]
port 4454 e
rlabel metal2 -1500 -66760 -1500 -66715 3 ROW_SEL[45]
port 4555 e
rlabel metal2 -1500 -68260 -1500 -68215 3 ROW_SEL[46]
port 4656 e
rlabel metal2 -1500 -69760 -1500 -69715 3 ROW_SEL[47]
port 4757 e
rlabel metal2 -1500 -71260 -1500 -71215 3 ROW_SEL[48]
port 4858 e
rlabel metal2 -1500 -72760 -1500 -72715 3 ROW_SEL[49]
port 4959 e
rlabel metal2 -1500 -74260 -1500 -74215 3 ROW_SEL[50]
port 5060 e
rlabel metal2 -1500 -75760 -1500 -75715 3 ROW_SEL[51]
port 5161 e
rlabel metal2 -1500 -77260 -1500 -77215 3 ROW_SEL[52]
port 5262 e
rlabel metal2 -1500 -78760 -1500 -78715 3 ROW_SEL[53]
port 5363 e
rlabel metal2 -1500 -80260 -1500 -80215 3 ROW_SEL[54]
port 5464 e
rlabel metal2 -1500 -81760 -1500 -81715 3 ROW_SEL[55]
port 5565 e
rlabel metal2 -1500 -83260 -1500 -83215 3 ROW_SEL[56]
port 5666 e
rlabel metal2 -1500 -84760 -1500 -84715 3 ROW_SEL[57]
port 5767 e
rlabel metal2 -1500 -86260 -1500 -86215 3 ROW_SEL[58]
port 5868 e
rlabel metal2 -1500 -87760 -1500 -87715 3 ROW_SEL[59]
port 5969 e
rlabel metal2 -1500 -89260 -1500 -89215 3 ROW_SEL[60]
port 6070 e
rlabel metal2 -1500 -90760 -1500 -90715 3 ROW_SEL[61]
port 6171 e
rlabel metal2 -1500 -92260 -1500 -92215 3 ROW_SEL[62]
port 6272 e
rlabel metal2 -1500 -93760 -1500 -93715 3 ROW_SEL[63]
port 6373 e
rlabel metal2 -1500 -95260 -1500 -95215 3 ROW_SEL[64]
port 6474 e
rlabel metal2 -1500 -96760 -1500 -96715 3 ROW_SEL[65]
port 6575 e
rlabel metal2 -1500 -98260 -1500 -98215 3 ROW_SEL[66]
port 6676 e
rlabel metal2 -1500 -99760 -1500 -99715 3 ROW_SEL[67]
port 6777 e
rlabel metal2 -1500 -101260 -1500 -101215 3 ROW_SEL[68]
port 6878 e
rlabel metal2 -1500 -102760 -1500 -102715 3 ROW_SEL[69]
port 6979 e
rlabel metal2 -1500 -104260 -1500 -104215 3 ROW_SEL[70]
port 7080 e
rlabel metal2 -1500 -105760 -1500 -105715 3 ROW_SEL[71]
port 7181 e
rlabel metal2 -1500 -107260 -1500 -107215 3 ROW_SEL[72]
port 7282 e
rlabel metal2 -1500 -108760 -1500 -108715 3 ROW_SEL[73]
port 7383 e
rlabel metal2 -1500 -110260 -1500 -110215 3 ROW_SEL[74]
port 7484 e
rlabel metal2 -1500 -111760 -1500 -111715 3 ROW_SEL[75]
port 7585 e
rlabel metal2 -1500 -113260 -1500 -113215 3 ROW_SEL[76]
port 7686 e
rlabel metal2 -1500 -114760 -1500 -114715 3 ROW_SEL[77]
port 7787 e
rlabel metal2 -1500 -116260 -1500 -116215 3 ROW_SEL[78]
port 7888 e
rlabel metal2 -1500 -117760 -1500 -117715 3 ROW_SEL[79]
port 7989 e
rlabel metal2 -1500 -119260 -1500 -119215 3 ROW_SEL[80]
port 8090 e
rlabel metal2 -1500 -120760 -1500 -120715 3 ROW_SEL[81]
port 8191 e
rlabel metal2 -1500 -122260 -1500 -122215 3 ROW_SEL[82]
port 8292 e
rlabel metal2 -1500 -123760 -1500 -123715 3 ROW_SEL[83]
port 8393 e
rlabel metal2 -1500 -125260 -1500 -125215 3 ROW_SEL[84]
port 8494 e
rlabel metal2 -1500 -126760 -1500 -126715 3 ROW_SEL[85]
port 8595 e
rlabel metal2 -1500 -128260 -1500 -128215 3 ROW_SEL[86]
port 8696 e
rlabel metal2 -1500 -129760 -1500 -129715 3 ROW_SEL[87]
port 8797 e
rlabel metal2 -1500 -131260 -1500 -131215 3 ROW_SEL[88]
port 8898 e
rlabel metal2 -1500 -132760 -1500 -132715 3 ROW_SEL[89]
port 8999 e
rlabel metal2 -1500 -134260 -1500 -134215 3 ROW_SEL[90]
port 9100 e
rlabel metal2 -1500 -135760 -1500 -135715 3 ROW_SEL[91]
port 9201 e
rlabel metal2 -1500 -137260 -1500 -137215 3 ROW_SEL[92]
port 9302 e
rlabel metal2 -1500 -138760 -1500 -138715 3 ROW_SEL[93]
port 9403 e
rlabel metal2 -1500 -140260 -1500 -140215 3 ROW_SEL[94]
port 9504 e
rlabel metal2 -1500 -141760 -1500 -141715 3 ROW_SEL[95]
port 9605 e
rlabel metal2 -1500 -143260 -1500 -143215 3 ROW_SEL[96]
port 9706 e
rlabel metal2 -1500 -144760 -1500 -144715 3 ROW_SEL[97]
port 9807 e
rlabel metal2 -1500 -146260 -1500 -146215 3 ROW_SEL[98]
port 9908 e
rlabel metal4 110 -149050 220 -149050 1 COL_SEL[0]
port 10010 n
rlabel metal4 -240 -149300 -240 -149300 1 CSA_VREF
port 10011 n
rlabel metal2 -1500 -147760 -1500 -147715 3 ROW_SEL[99]
port 10012 e
rlabel metal4 1610 -149050 1720 -149050 1 COL_SEL[1]
port 10015 n
rlabel metal4 3110 -149050 3220 -149050 1 COL_SEL[2]
port 10018 n
rlabel metal4 4610 -149050 4720 -149050 1 COL_SEL[3]
port 10021 n
rlabel metal4 6110 -149050 6220 -149050 1 COL_SEL[4]
port 10024 n
rlabel metal4 7610 -149050 7720 -149050 1 COL_SEL[5]
port 10027 n
rlabel metal4 9110 -149050 9220 -149050 1 COL_SEL[6]
port 10030 n
rlabel metal4 10610 -149050 10720 -149050 1 COL_SEL[7]
port 10033 n
rlabel metal4 12110 -149050 12220 -149050 1 COL_SEL[8]
port 10036 n
rlabel metal4 13610 -149050 13720 -149050 1 COL_SEL[9]
port 10039 n
rlabel metal4 15110 -149050 15220 -149050 1 COL_SEL[10]
port 10042 n
rlabel metal4 16610 -149050 16720 -149050 1 COL_SEL[11]
port 10045 n
rlabel metal4 18110 -149050 18220 -149050 1 COL_SEL[12]
port 10048 n
rlabel metal4 19610 -149050 19720 -149050 1 COL_SEL[13]
port 10051 n
rlabel metal4 21110 -149050 21220 -149050 1 COL_SEL[14]
port 10054 n
rlabel metal4 22610 -149050 22720 -149050 1 COL_SEL[15]
port 10057 n
rlabel metal4 24110 -149050 24220 -149050 1 COL_SEL[16]
port 10060 n
rlabel metal4 25610 -149050 25720 -149050 1 COL_SEL[17]
port 10063 n
rlabel metal4 27110 -149050 27220 -149050 1 COL_SEL[18]
port 10066 n
rlabel metal4 28610 -149050 28720 -149050 1 COL_SEL[19]
port 10069 n
rlabel metal4 30110 -149050 30220 -149050 1 COL_SEL[20]
port 10072 n
rlabel metal4 31610 -149050 31720 -149050 1 COL_SEL[21]
port 10075 n
rlabel metal4 33110 -149050 33220 -149050 1 COL_SEL[22]
port 10078 n
rlabel metal4 34610 -149050 34720 -149050 1 COL_SEL[23]
port 10081 n
rlabel metal4 36110 -149050 36220 -149050 1 COL_SEL[24]
port 10084 n
rlabel metal4 37610 -149050 37720 -149050 1 COL_SEL[25]
port 10087 n
rlabel metal4 39110 -149050 39220 -149050 1 COL_SEL[26]
port 10090 n
rlabel metal4 40610 -149050 40720 -149050 1 COL_SEL[27]
port 10093 n
rlabel metal4 42110 -149050 42220 -149050 1 COL_SEL[28]
port 10096 n
rlabel metal4 43610 -149050 43720 -149050 1 COL_SEL[29]
port 10099 n
rlabel metal4 45110 -149050 45220 -149050 1 COL_SEL[30]
port 10102 n
rlabel metal4 46610 -149050 46720 -149050 1 COL_SEL[31]
port 10105 n
rlabel metal4 48110 -149050 48220 -149050 1 COL_SEL[32]
port 10108 n
rlabel metal4 49610 -149050 49720 -149050 1 COL_SEL[33]
port 10111 n
rlabel metal4 51110 -149050 51220 -149050 1 COL_SEL[34]
port 10114 n
rlabel metal4 52610 -149050 52720 -149050 1 COL_SEL[35]
port 10117 n
rlabel metal4 54110 -149050 54220 -149050 1 COL_SEL[36]
port 10120 n
rlabel metal4 55610 -149050 55720 -149050 1 COL_SEL[37]
port 10123 n
rlabel metal4 57110 -149050 57220 -149050 1 COL_SEL[38]
port 10126 n
rlabel metal4 58610 -149050 58720 -149050 1 COL_SEL[39]
port 10129 n
rlabel metal4 60110 -149050 60220 -149050 1 COL_SEL[40]
port 10132 n
rlabel metal4 61610 -149050 61720 -149050 1 COL_SEL[41]
port 10135 n
rlabel metal4 63110 -149050 63220 -149050 1 COL_SEL[42]
port 10138 n
rlabel metal4 64610 -149050 64720 -149050 1 COL_SEL[43]
port 10141 n
rlabel metal4 66110 -149050 66220 -149050 1 COL_SEL[44]
port 10144 n
rlabel metal4 67610 -149050 67720 -149050 1 COL_SEL[45]
port 10147 n
rlabel metal4 69110 -149050 69220 -149050 1 COL_SEL[46]
port 10150 n
rlabel metal4 70610 -149050 70720 -149050 1 COL_SEL[47]
port 10153 n
rlabel metal4 72110 -149050 72220 -149050 1 COL_SEL[48]
port 10156 n
rlabel metal4 73610 -149050 73720 -149050 1 COL_SEL[49]
port 10159 n
rlabel metal4 75110 -149050 75220 -149050 1 COL_SEL[50]
port 10162 n
rlabel metal4 76610 -149050 76720 -149050 1 COL_SEL[51]
port 10165 n
rlabel metal4 78110 -149050 78220 -149050 1 COL_SEL[52]
port 10168 n
rlabel metal4 79610 -149050 79720 -149050 1 COL_SEL[53]
port 10171 n
rlabel metal4 81110 -149050 81220 -149050 1 COL_SEL[54]
port 10174 n
rlabel metal4 82610 -149050 82720 -149050 1 COL_SEL[55]
port 10177 n
rlabel metal4 84110 -149050 84220 -149050 1 COL_SEL[56]
port 10180 n
rlabel metal4 85610 -149050 85720 -149050 1 COL_SEL[57]
port 10183 n
rlabel metal4 87110 -149050 87220 -149050 1 COL_SEL[58]
port 10186 n
rlabel metal4 88610 -149050 88720 -149050 1 COL_SEL[59]
port 10189 n
rlabel metal4 90110 -149050 90220 -149050 1 COL_SEL[60]
port 10192 n
rlabel metal4 91610 -149050 91720 -149050 1 COL_SEL[61]
port 10195 n
rlabel metal4 93110 -149050 93220 -149050 1 COL_SEL[62]
port 10198 n
rlabel metal4 94610 -149050 94720 -149050 1 COL_SEL[63]
port 10201 n
rlabel metal4 96110 -149050 96220 -149050 1 COL_SEL[64]
port 10204 n
rlabel metal4 97610 -149050 97720 -149050 1 COL_SEL[65]
port 10207 n
rlabel metal4 99110 -149050 99220 -149050 1 COL_SEL[66]
port 10210 n
rlabel metal4 100610 -149050 100720 -149050 1 COL_SEL[67]
port 10213 n
rlabel metal4 102110 -149050 102220 -149050 1 COL_SEL[68]
port 10216 n
rlabel metal4 103610 -149050 103720 -149050 1 COL_SEL[69]
port 10219 n
rlabel metal4 105110 -149050 105220 -149050 1 COL_SEL[70]
port 10222 n
rlabel metal4 106610 -149050 106720 -149050 1 COL_SEL[71]
port 10225 n
rlabel metal4 108110 -149050 108220 -149050 1 COL_SEL[72]
port 10228 n
rlabel metal4 109610 -149050 109720 -149050 1 COL_SEL[73]
port 10231 n
rlabel metal4 111110 -149050 111220 -149050 1 COL_SEL[74]
port 10234 n
rlabel metal4 112610 -149050 112720 -149050 1 COL_SEL[75]
port 10237 n
rlabel metal4 114110 -149050 114220 -149050 1 COL_SEL[76]
port 10240 n
rlabel metal4 115610 -149050 115720 -149050 1 COL_SEL[77]
port 10243 n
rlabel metal4 117110 -149050 117220 -149050 1 COL_SEL[78]
port 10246 n
rlabel metal4 118610 -149050 118720 -149050 1 COL_SEL[79]
port 10249 n
rlabel metal4 120110 -149050 120220 -149050 1 COL_SEL[80]
port 10252 n
rlabel metal4 121610 -149050 121720 -149050 1 COL_SEL[81]
port 10255 n
rlabel metal4 123110 -149050 123220 -149050 1 COL_SEL[82]
port 10258 n
rlabel metal4 124610 -149050 124720 -149050 1 COL_SEL[83]
port 10261 n
rlabel metal4 126110 -149050 126220 -149050 1 COL_SEL[84]
port 10264 n
rlabel metal4 127610 -149050 127720 -149050 1 COL_SEL[85]
port 10267 n
rlabel metal4 129110 -149050 129220 -149050 1 COL_SEL[86]
port 10270 n
rlabel metal4 130610 -149050 130720 -149050 1 COL_SEL[87]
port 10273 n
rlabel metal4 132110 -149050 132220 -149050 1 COL_SEL[88]
port 10276 n
rlabel metal4 133610 -149050 133720 -149050 1 COL_SEL[89]
port 10279 n
rlabel metal4 135110 -149050 135220 -149050 1 COL_SEL[90]
port 10282 n
rlabel metal4 136610 -149050 136720 -149050 1 COL_SEL[91]
port 10285 n
rlabel metal4 138110 -149050 138220 -149050 1 COL_SEL[92]
port 10288 n
rlabel metal4 139610 -149050 139720 -149050 1 COL_SEL[93]
port 10291 n
rlabel metal4 141110 -149050 141220 -149050 1 COL_SEL[94]
port 10294 n
rlabel metal4 142610 -149050 142720 -149050 1 COL_SEL[95]
port 10297 n
rlabel metal4 144110 -149050 144220 -149050 1 COL_SEL[96]
port 10300 n
rlabel metal4 145610 -149050 145720 -149050 1 COL_SEL[97]
port 10303 n
rlabel metal4 147110 -149050 147220 -149050 1 COL_SEL[98]
port 10306 n
rlabel metal2 149970 -149050 149970 -149050 1 ARRAY_OUT
port 10309 n
rlabel metal4 148610 -149050 148720 -149050 1 COL_SEL[99]
port 10310 n
rlabel metal3 -573 2441 -573 2441 1 SF_IB
port 10311 n
<< end >>
